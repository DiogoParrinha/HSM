-- Version: v11.7 SP1 11.7.1.14

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_controller is

    port( sha256_controller_0_read_addr_0 : out   std_logic_vector(3 downto 0);
          sha256_controller_0_bytes_o     : out   std_logic_vector(1 to 1);
          state_out_net_0                 : out   std_logic_vector(0 to 0);
          state_4                         : out   std_logic;
          state_3                         : out   std_logic;
          state_1                         : out   std_logic;
          ce_i_i_2                        : out   std_logic;
          ce_i_i_2_i_0                    : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK    : in    std_logic;
          sha256_system_sb_0_GPIO_9_M2F   : in    std_logic;
          sha256_controller_0_end_o       : out   std_logic;
          last_block_0                    : out   std_logic;
          N_88_i_0                        : out   std_logic;
          N_28                            : out   std_logic;
          SHA256_Module_0_di_req_o        : in    std_logic;
          N_89                            : out   std_logic;
          SHA256_Module_0_do_valid_o      : in    std_logic;
          last_block                      : in    std_logic;
          prev_sig                        : in    std_logic;
          first_block                     : in    std_logic;
          SHA256_Module_0_data_out_ready  : in    std_logic;
          prev_sig_0                      : in    std_logic;
          N_87_i_0                        : out   std_logic
        );

end sha256_controller;

architecture DEF_ARCH of sha256_controller is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal un2_rst_n_i, \un2_rst_n\, \blocks_counter[0]_net_1\, 
        \blocks_counter_s[0]\, \ce_i_i_2\, 
        \sha256_controller_0_read_addr_0[0]\, VCC_net_1, 
        un5_rst_n_i, N_139_i_0, GND_net_1, 
        \sha256_controller_0_read_addr_0[1]\, \counter_4[1]\, 
        \sha256_controller_0_read_addr_0[2]\, \counter_4[2]\, 
        \sha256_controller_0_read_addr_0[3]\, N_11_i_0, 
        \state_ns[0]\, \state_4\, N_71_i_0, \state_3\, N_73_i_0, 
        \state[2]_net_1\, \state_ns_i_i[3]_net_1\, \state_1\, 
        \state_ns[4]\, \state[0]_net_1\, \state_ns[5]\, 
        \un1_state_1_0_a2_0_a2\, end_o_1_sqmuxa_i_0, \extra_add\, 
        \un1_extra_add_1_sqmuxa_0_0\, start_o_1_sqmuxa_i_0, 
        \blocks_counter[1]_net_1\, \blocks_counter_s[1]\, 
        \blocks_counter[2]_net_1\, \blocks_counter_s[2]\, 
        \blocks_counter[3]_net_1\, \blocks_counter_s[3]\, 
        \blocks_counter[4]_net_1\, \blocks_counter_s[4]\, 
        \blocks_counter[5]_net_1\, \blocks_counter_s[5]\, 
        \blocks_counter[6]_net_1\, \blocks_counter_s[6]\, 
        \blocks_counter[7]_net_1\, \blocks_counter_s[7]\, 
        \blocks_counter[8]_net_1\, \blocks_counter_s[8]\, 
        \blocks_counter[9]_net_1\, \blocks_counter_s[9]\, 
        \blocks_counter[10]_net_1\, \blocks_counter_s[10]\, 
        \blocks_counter[11]_net_1\, \blocks_counter_s[11]\, 
        \blocks_counter[12]_net_1\, \blocks_counter_s[12]\, 
        \blocks_counter[13]_net_1\, \blocks_counter_s[13]\, 
        \blocks_counter[14]_net_1\, \blocks_counter_s[14]\, 
        \blocks_counter[15]_net_1\, \blocks_counter_s[15]\, 
        \blocks_counter[16]_net_1\, \blocks_counter_s[16]\, 
        \blocks_counter[17]_net_1\, \blocks_counter_s[17]\, 
        \blocks_counter[18]_net_1\, \blocks_counter_s[18]\, 
        \blocks_counter[19]_net_1\, \blocks_counter_s[19]\, 
        \blocks_counter[20]_net_1\, \blocks_counter_s[20]\, 
        \blocks_counter[21]_net_1\, \blocks_counter_s[21]\, 
        \blocks_counter[22]_net_1\, \blocks_counter_s[22]\, 
        \blocks_counter[23]_net_1\, \blocks_counter_s[23]\, 
        \blocks_counter[24]_net_1\, \blocks_counter_s[24]\, 
        \blocks_counter[25]_net_1\, \blocks_counter_s[25]\, 
        \blocks_counter[26]_net_1\, \blocks_counter_s[26]\, 
        \blocks_counter[27]_net_1\, \blocks_counter_s[27]\, 
        \blocks_counter[28]_net_1\, \blocks_counter_s[28]\, 
        \blocks_counter[29]_net_1\, \blocks_counter_s[29]\, 
        \blocks_counter[30]_net_1\, \blocks_counter_s[30]\, 
        \blocks_counter[31]_net_1\, \blocks_counter_s[31]_net_1\, 
        blocks_counter_s_991_FCO, \blocks_counter_cry[1]_net_1\, 
        \blocks_counter_cry[2]_net_1\, 
        \blocks_counter_cry[3]_net_1\, 
        \blocks_counter_cry[4]_net_1\, 
        \blocks_counter_cry[5]_net_1\, 
        \blocks_counter_cry[6]_net_1\, 
        \blocks_counter_cry[7]_net_1\, 
        \blocks_counter_cry[8]_net_1\, 
        \blocks_counter_cry[9]_net_1\, 
        \blocks_counter_cry[10]_net_1\, 
        \blocks_counter_cry[11]_net_1\, 
        \blocks_counter_cry[12]_net_1\, 
        \blocks_counter_cry[13]_net_1\, 
        \blocks_counter_cry[14]_net_1\, 
        \blocks_counter_cry[15]_net_1\, 
        \blocks_counter_cry[16]_net_1\, 
        \blocks_counter_cry[17]_net_1\, 
        \blocks_counter_cry[18]_net_1\, 
        \blocks_counter_cry[19]_net_1\, 
        \blocks_counter_cry[20]_net_1\, 
        \blocks_counter_cry[21]_net_1\, 
        \blocks_counter_cry[22]_net_1\, 
        \blocks_counter_cry[23]_net_1\, 
        \blocks_counter_cry[24]_net_1\, 
        \blocks_counter_cry[25]_net_1\, 
        \blocks_counter_cry[26]_net_1\, 
        \blocks_counter_cry[27]_net_1\, 
        \blocks_counter_cry[28]_net_1\, 
        \blocks_counter_cry[29]_net_1\, 
        \blocks_counter_cry[30]_net_1\, N_141, N_182, N_30, 
        \N_28\, start_o2_23, start_o2_22, start_o2_21, 
        start_o2_20, start_o2_19, start_o2_18, start_o2_17, 
        start_o2_16, \un1_extra_add_1_sqmuxa_0_0_a2_2\, N_29, 
        N_179, start_o2_29, start_o2_28 : std_logic;

begin 

    sha256_controller_0_read_addr_0(3) <= 
        \sha256_controller_0_read_addr_0[3]\;
    sha256_controller_0_read_addr_0(2) <= 
        \sha256_controller_0_read_addr_0[2]\;
    sha256_controller_0_read_addr_0(1) <= 
        \sha256_controller_0_read_addr_0[1]\;
    sha256_controller_0_read_addr_0(0) <= 
        \sha256_controller_0_read_addr_0[0]\;
    state_4 <= \state_4\;
    state_3 <= \state_3\;
    state_1 <= \state_1\;
    ce_i_i_2 <= \ce_i_i_2\;
    N_28 <= \N_28\;

    \op_eq.start_o2_19\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[15]_net_1\, B => 
        \blocks_counter[14]_net_1\, C => 
        \blocks_counter[13]_net_1\, D => 
        \blocks_counter[12]_net_1\, Y => start_o2_19);
    
    \blocks_counter_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[2]_net_1\, S => \blocks_counter_s[3]\, 
        Y => OPEN, FCO => \blocks_counter_cry[3]_net_1\);
    
    \blocks_counter_cry[26]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[26]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[25]_net_1\, S => 
        \blocks_counter_s[26]\, Y => OPEN, FCO => 
        \blocks_counter_cry[26]_net_1\);
    
    \blocks_counter[31]\ : SLE
      port map(D => \blocks_counter_s[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[31]_net_1\);
    
    \blocks_counter_s[31]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[31]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[30]_net_1\, S => 
        \blocks_counter_s[31]_net_1\, Y => OPEN, FCO => OPEN);
    
    \blocks_counter_cry[22]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[22]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[21]_net_1\, S => 
        \blocks_counter_s[22]\, Y => OPEN, FCO => 
        \blocks_counter_cry[22]_net_1\);
    
    \blocks_counter_cry[25]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[25]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[24]_net_1\, S => 
        \blocks_counter_s[25]\, Y => OPEN, FCO => 
        \blocks_counter_cry[25]_net_1\);
    
    un1_state_1_0_a2_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \state[2]_net_1\, B => \state[0]_net_1\, Y
         => \un1_state_1_0_a2_0_a2\);
    
    \op_eq.start_o2_22\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[27]_net_1\, B => 
        \blocks_counter[26]_net_1\, C => 
        \blocks_counter[25]_net_1\, D => 
        \blocks_counter[24]_net_1\, Y => start_o2_22);
    
    \blocks_counter_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        blocks_counter_s_991_FCO, S => \blocks_counter_s[1]\, Y
         => OPEN, FCO => \blocks_counter_cry[1]_net_1\);
    
    \blocks_counter_cry[16]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[16]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[15]_net_1\, S => 
        \blocks_counter_s[16]\, Y => OPEN, FCO => 
        \blocks_counter_cry[16]_net_1\);
    
    \state_RNO[3]\ : CFG4
      generic map(INIT => x"AA20")

      port map(A => SHA256_Module_0_di_req_o, B => N_182, C => 
        \state_3\, D => \state[2]_net_1\, Y => N_73_i_0);
    
    \counter[2]\ : SLE
      port map(D => \counter_4[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        un5_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \sha256_controller_0_read_addr_0[2]\);
    
    \counter_4_0_o2[1]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \sha256_controller_0_read_addr_0[2]\, B => 
        \sha256_controller_0_read_addr_0[3]\, Y => N_141);
    
    \blocks_counter_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[11]_net_1\, S => 
        \blocks_counter_s[12]\, Y => OPEN, FCO => 
        \blocks_counter_cry[12]_net_1\);
    
    \blocks_counter[20]\ : SLE
      port map(D => \blocks_counter_s[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[20]_net_1\);
    
    \blocks_counter[13]\ : SLE
      port map(D => \blocks_counter_s[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[13]_net_1\);
    
    \state[5]\ : SLE
      port map(D => \state_ns[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_0_GPIO_9_M2F, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ce_i_i_2\);
    
    \blocks_counter_cry[15]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[14]_net_1\, S => 
        \blocks_counter_s[15]\, Y => OPEN, FCO => 
        \blocks_counter_cry[15]_net_1\);
    
    \blocks_counter[26]\ : SLE
      port map(D => \blocks_counter_s[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[26]_net_1\);
    
    \blocks_counter[15]\ : SLE
      port map(D => \blocks_counter_s[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[15]_net_1\);
    
    \state_out_a3_0_a2[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \un1_state_1_0_a2_0_a2\, B => \state_4\, Y
         => state_out_net_0(0));
    
    \blocks_counter[30]\ : SLE
      port map(D => \blocks_counter_s[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[30]_net_1\);
    
    \state[4]\ : SLE
      port map(D => N_71_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => sha256_system_sb_0_GPIO_9_M2F, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \state_4\);
    
    \blocks_counter[0]\ : SLE
      port map(D => \blocks_counter_s[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[0]_net_1\);
    
    \blocks_counter_cry[23]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[23]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[22]_net_1\, S => 
        \blocks_counter_s[23]\, Y => OPEN, FCO => 
        \blocks_counter_cry[23]_net_1\);
    
    \counter_RNO[0]\ : CFG4
      generic map(INIT => x"33C4")

      port map(A => \sha256_controller_0_read_addr_0[1]\, B => 
        \sha256_controller_0_read_addr_0[0]\, C => N_141, D => 
        N_29, Y => N_139_i_0);
    
    \state_ns_i_i[3]\ : CFG4
      generic map(INIT => x"FF0E")

      port map(A => \state[2]_net_1\, B => \state_3\, C => 
        SHA256_Module_0_di_req_o, D => \state_4\, Y => 
        \state_ns_i_i[3]_net_1\);
    
    \state[2]\ : SLE
      port map(D => \state_ns_i_i[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_0_GPIO_9_M2F, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[2]_net_1\);
    
    \counter_4_0_o2_0[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \N_28\, B => \extra_add\, Y => N_29);
    
    \op_eq.start_o2_29\ : CFG4
      generic map(INIT => x"8000")

      port map(A => start_o2_23, B => start_o2_22, C => 
        start_o2_21, D => start_o2_20, Y => start_o2_29);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    un1_extra_add_1_sqmuxa_0_0 : CFG4
      generic map(INIT => x"10FF")

      port map(A => \sha256_controller_0_read_addr_0[3]\, B => 
        \sha256_controller_0_read_addr_0[1]\, C => 
        \un1_extra_add_1_sqmuxa_0_0_a2_2\, D => \state[2]_net_1\, 
        Y => \un1_extra_add_1_sqmuxa_0_0\);
    
    \state_RNI2S0E[5]\ : CFG1
      generic map(INIT => "01")

      port map(A => \ce_i_i_2\, Y => ce_i_i_2_i_0);
    
    \blocks_counter[11]\ : SLE
      port map(D => \blocks_counter_s[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[11]_net_1\);
    
    \op_eq.start_o2_18\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[11]_net_1\, B => 
        \blocks_counter[10]_net_1\, C => 
        \blocks_counter[9]_net_1\, D => \blocks_counter[8]_net_1\, 
        Y => start_o2_18);
    
    \state[3]\ : SLE
      port map(D => N_73_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => sha256_system_sb_0_GPIO_9_M2F, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \state_3\);
    
    \blocks_counter_cry[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[12]_net_1\, S => 
        \blocks_counter_s[13]\, Y => OPEN, FCO => 
        \blocks_counter_cry[13]_net_1\);
    
    \counter_4_0_o2[2]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \sha256_controller_0_read_addr_0[0]\, B => 
        \sha256_controller_0_read_addr_0[1]\, Y => N_30);
    
    \blocks_counter_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[1]_net_1\, S => \blocks_counter_s[2]\, 
        Y => OPEN, FCO => \blocks_counter_cry[2]_net_1\);
    
    \blocks_counter_cry[27]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[27]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[26]_net_1\, S => 
        \blocks_counter_s[27]\, Y => OPEN, FCO => 
        \blocks_counter_cry[27]_net_1\);
    
    \op_eq.start_o2_23\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[31]_net_1\, B => 
        \blocks_counter[30]_net_1\, C => 
        \blocks_counter[29]_net_1\, D => 
        \blocks_counter[28]_net_1\, Y => start_o2_23);
    
    \blocks_counter[24]\ : SLE
      port map(D => \blocks_counter_s[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[24]_net_1\);
    
    \blocks_counter_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[5]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[4]_net_1\, S => \blocks_counter_s[5]\, 
        Y => OPEN, FCO => \blocks_counter_cry[5]_net_1\);
    
    \blocks_counter_cry[28]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[28]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[27]_net_1\, S => 
        \blocks_counter_s[28]\, Y => OPEN, FCO => 
        \blocks_counter_cry[28]_net_1\);
    
    \blocks_counter[22]\ : SLE
      port map(D => \blocks_counter_s[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[22]_net_1\);
    
    \op_eq.start_o2_20\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[19]_net_1\, B => 
        \blocks_counter[18]_net_1\, C => 
        \blocks_counter[17]_net_1\, D => 
        \blocks_counter[16]_net_1\, Y => start_o2_20);
    
    \blocks_counter_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[8]_net_1\, S => \blocks_counter_s[9]\, 
        Y => OPEN, FCO => \blocks_counter_cry[9]_net_1\);
    
    un2_rst_n_RNIE1K2 : CLKINT
      port map(A => \un2_rst_n\, Y => un2_rst_n_i);
    
    \blocks_counter_cry[17]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[17]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[16]_net_1\, S => 
        \blocks_counter_s[17]\, Y => OPEN, FCO => 
        \blocks_counter_cry[17]_net_1\);
    
    \blocks_counter[5]\ : SLE
      port map(D => \blocks_counter_s[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[5]_net_1\);
    
    \blocks_counter[10]\ : SLE
      port map(D => \blocks_counter_s[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[10]_net_1\);
    
    \blocks_counter[16]\ : SLE
      port map(D => \blocks_counter_s[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[16]_net_1\);
    
    \counter_4_0[1]\ : CFG4
      generic map(INIT => x"66A2")

      port map(A => \sha256_controller_0_read_addr_0[1]\, B => 
        \sha256_controller_0_read_addr_0[0]\, C => N_141, D => 
        N_29, Y => \counter_4[1]\);
    
    sel_di_i_a3_0_a2 : CFG3
      generic map(INIT => x"01")

      port map(A => \state_1\, B => \state_4\, C => \state_3\, Y
         => N_89);
    
    \blocks_counter_cry[18]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[18]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[17]_net_1\, S => 
        \blocks_counter_s[18]\, Y => OPEN, FCO => 
        \blocks_counter_cry[18]_net_1\);
    
    \state_ns_a3_0_a2[4]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SHA256_Module_0_di_req_o, B => N_182, C => 
        \state_3\, Y => \state_ns[4]\);
    
    \op_eq.start_o2_28\ : CFG4
      generic map(INIT => x"8000")

      port map(A => start_o2_19, B => start_o2_18, C => 
        start_o2_17, D => start_o2_16, Y => start_o2_28);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \blocks_counter[1]\ : SLE
      port map(D => \blocks_counter_s[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[1]_net_1\);
    
    \blocks_counter[8]\ : SLE
      port map(D => \blocks_counter_s[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[8]_net_1\);
    
    \state[0]\ : SLE
      port map(D => \state_ns[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_0_GPIO_9_M2F, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[0]_net_1\);
    
    \blocks_counter[2]\ : SLE
      port map(D => \blocks_counter_s[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[2]_net_1\);
    
    end_o_1_sqmuxa_i : CFG2
      generic map(INIT => x"B")

      port map(A => last_block, B => \state_1\, Y => 
        end_o_1_sqmuxa_i_0);
    
    \blocks_counter[27]\ : SLE
      port map(D => \blocks_counter_s[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[27]_net_1\);
    
    \blocks_counter[3]\ : SLE
      port map(D => \blocks_counter_s[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[3]_net_1\);
    
    start_o : SLE
      port map(D => \state_4\, CLK => start_o_1_sqmuxa_i_0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        last_block_0);
    
    un1_extra_add_1_sqmuxa_0_0_a2_2 : CFG3
      generic map(INIT => x"02")

      port map(A => SHA256_Module_0_di_req_o, B => 
        \sha256_controller_0_read_addr_0[2]\, C => 
        \sha256_controller_0_read_addr_0[0]\, Y => 
        \un1_extra_add_1_sqmuxa_0_0_a2_2\);
    
    \counter_RNO[3]\ : CFG4
      generic map(INIT => x"A6A2")

      port map(A => \sha256_controller_0_read_addr_0[3]\, B => 
        \sha256_controller_0_read_addr_0[2]\, C => N_30, D => 
        N_29, Y => N_11_i_0);
    
    \state_RNIQ72A1[0]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \state[0]_net_1\, B => \state[2]_net_1\, C
         => \state_1\, Y => N_88_i_0);
    
    blocks_counter_s_991 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => blocks_counter_s_991_FCO);
    
    \blocks_counter_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[7]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[6]_net_1\, S => \blocks_counter_s[7]\, 
        Y => OPEN, FCO => \blocks_counter_cry[7]_net_1\);
    
    \blocks_counter_cry[30]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[30]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[29]_net_1\, S => 
        \blocks_counter_s[30]\, Y => OPEN, FCO => 
        \blocks_counter_cry[30]_net_1\);
    
    \blocks_counter[14]\ : SLE
      port map(D => \blocks_counter_s[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[14]_net_1\);
    
    \counter[1]\ : SLE
      port map(D => \counter_4[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        un5_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \sha256_controller_0_read_addr_0[1]\);
    
    \blocks_counter[12]\ : SLE
      port map(D => \blocks_counter_s[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[12]_net_1\);
    
    \counter[3]\ : SLE
      port map(D => N_11_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => un5_rst_n_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sha256_controller_0_read_addr_0[3]\);
    
    \blocks_counter_cry[21]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[21]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[20]_net_1\, S => 
        \blocks_counter_s[21]\, Y => OPEN, FCO => 
        \blocks_counter_cry[21]_net_1\);
    
    \op_eq.start_o2_16\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[3]_net_1\, B => 
        \blocks_counter[2]_net_1\, C => \blocks_counter[1]_net_1\, 
        D => \blocks_counter[0]_net_1\, Y => start_o2_16);
    
    \counter_4_i_a2_0[3]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \sha256_controller_0_read_addr_0[0]\, B => 
        N_141, C => \sha256_controller_0_read_addr_0[1]\, Y => 
        N_182);
    
    \state_RNO[4]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \ce_i_i_2\, B => 
        SHA256_Module_0_data_out_ready, C => prev_sig_0, Y => 
        N_71_i_0);
    
    \blocks_counter_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \blocks_counter[0]_net_1\, Y => 
        \blocks_counter_s[0]\);
    
    \blocks_counter_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[4]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[3]_net_1\, S => \blocks_counter_s[4]\, 
        Y => OPEN, FCO => \blocks_counter_cry[4]_net_1\);
    
    \blocks_counter_cry[29]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[29]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[28]_net_1\, S => 
        \blocks_counter_s[29]\, Y => OPEN, FCO => 
        \blocks_counter_cry[29]_net_1\);
    
    \blocks_counter[28]\ : SLE
      port map(D => \blocks_counter_s[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[28]_net_1\);
    
    \state_ns_0_a2[0]\ : CFG3
      generic map(INIT => x"C8")

      port map(A => SHA256_Module_0_di_req_o, B => 
        \state[0]_net_1\, C => SHA256_Module_0_do_valid_o, Y => 
        N_179);
    
    extra_add : SLE
      port map(D => \state[2]_net_1\, CLK => 
        \un1_extra_add_1_sqmuxa_0_0\, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => VCC_net_1, Q => \extra_add\);
    
    \blocks_counter_cry[20]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[20]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[19]_net_1\, S => 
        \blocks_counter_s[20]\, Y => OPEN, FCO => 
        \blocks_counter_cry[20]_net_1\);
    
    \blocks_counter[29]\ : SLE
      port map(D => \blocks_counter_s[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[29]_net_1\);
    
    \state[1]\ : SLE
      port map(D => \state_ns[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_0_GPIO_9_M2F, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state_1\);
    
    \blocks_counter_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[6]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[5]_net_1\, S => \blocks_counter_s[6]\, 
        Y => OPEN, FCO => \blocks_counter_cry[6]_net_1\);
    
    \blocks_counter[6]\ : SLE
      port map(D => \blocks_counter_s[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[6]_net_1\);
    
    \op_eq.start_o2_17\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[7]_net_1\, B => 
        \blocks_counter[6]_net_1\, C => \blocks_counter[5]_net_1\, 
        D => \blocks_counter[4]_net_1\, Y => start_o2_17);
    
    \blocks_counter_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[10]_net_1\, S => 
        \blocks_counter_s[11]\, Y => OPEN, FCO => 
        \blocks_counter_cry[11]_net_1\);
    
    \blocks_counter_cry[19]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[19]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[18]_net_1\, S => 
        \blocks_counter_s[19]\, Y => OPEN, FCO => 
        \blocks_counter_cry[19]_net_1\);
    
    \blocks_counter[17]\ : SLE
      port map(D => \blocks_counter_s[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[17]_net_1\);
    
    \blocks_counter_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[9]_net_1\, S => 
        \blocks_counter_s[10]\, Y => OPEN, FCO => 
        \blocks_counter_cry[10]_net_1\);
    
    start_o_1_sqmuxa_i : CFG3
      generic map(INIT => x"D5")

      port map(A => \state_4\, B => start_o2_29, C => start_o2_28, 
        Y => start_o_1_sqmuxa_i_0);
    
    \blocks_counter_cry[24]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[24]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[23]_net_1\, S => 
        \blocks_counter_s[24]\, Y => OPEN, FCO => 
        \blocks_counter_cry[24]_net_1\);
    
    \state_RNIUH1S[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \state_1\, B => \state_3\, Y => \N_28\);
    
    \blocks_counter[7]\ : SLE
      port map(D => \blocks_counter_s[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[7]_net_1\);
    
    un5_rst_n : CFG2
      generic map(INIT => x"4")

      port map(A => \ce_i_i_2\, B => 
        sha256_system_sb_0_GPIO_9_M2F, Y => un5_rst_n_i);
    
    \state_ns_0[5]\ : CFG4
      generic map(INIT => x"AAAE")

      port map(A => \state_1\, B => \state[0]_net_1\, C => 
        SHA256_Module_0_di_req_o, D => SHA256_Module_0_do_valid_o, 
        Y => \state_ns[5]\);
    
    \blocks_counter_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[7]_net_1\, S => \blocks_counter_s[8]\, 
        Y => OPEN, FCO => \blocks_counter_cry[8]_net_1\);
    
    \blocks_counter_cry[14]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[13]_net_1\, S => 
        \blocks_counter_s[14]\, Y => OPEN, FCO => 
        \blocks_counter_cry[14]_net_1\);
    
    \blocks_counter[23]\ : SLE
      port map(D => \blocks_counter_s[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[23]_net_1\);
    
    \op_eq.start_o2_21\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[23]_net_1\, B => 
        \blocks_counter[22]_net_1\, C => 
        \blocks_counter[21]_net_1\, D => 
        \blocks_counter[20]_net_1\, Y => start_o2_21);
    
    \blocks_counter[25]\ : SLE
      port map(D => \blocks_counter_s[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[25]_net_1\);
    
    \counter_4_0[2]\ : CFG4
      generic map(INIT => x"C3C4")

      port map(A => \sha256_controller_0_read_addr_0[3]\, B => 
        \sha256_controller_0_read_addr_0[2]\, C => N_30, D => 
        N_29, Y => \counter_4[2]\);
    
    \state_RNIUB2A1[0]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \state[0]_net_1\, B => \state_3\, C => 
        \state_4\, Y => N_87_i_0);
    
    end_o : SLE
      port map(D => \state_1\, CLK => end_o_1_sqmuxa_i_0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        sha256_controller_0_end_o);
    
    \blocks_counter[4]\ : SLE
      port map(D => \blocks_counter_s[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[4]_net_1\);
    
    \blocks_counter[18]\ : SLE
      port map(D => \blocks_counter_s[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[18]_net_1\);
    
    un2_rst_n : CFG3
      generic map(INIT => x"8A")

      port map(A => sha256_system_sb_0_GPIO_9_M2F, B => prev_sig, 
        C => first_block, Y => \un2_rst_n\);
    
    \blocks_counter[19]\ : SLE
      port map(D => \blocks_counter_s[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[19]_net_1\);
    
    \bytes_o[0]\ : SLE
      port map(D => GND_net_1, CLK => \un1_state_1_0_a2_0_a2\, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        sha256_controller_0_bytes_o(1));
    
    \counter[0]\ : SLE
      port map(D => N_139_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        un5_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \sha256_controller_0_read_addr_0[0]\);
    
    \blocks_counter[9]\ : SLE
      port map(D => \blocks_counter_s[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[9]_net_1\);
    
    \blocks_counter[21]\ : SLE
      port map(D => \blocks_counter_s[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \state_4\, ALn => 
        un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[21]_net_1\);
    
    \state_ns_0[0]\ : CFG4
      generic map(INIT => x"FDCC")

      port map(A => SHA256_Module_0_data_out_ready, B => N_179, C
         => prev_sig_0, D => \ce_i_i_2\, Y => \state_ns[0]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_control is

    port( hash_control_st_reg_i           : out   std_logic_vector(6 to 6);
          msg_bitlen                      : out   std_logic_vector(63 downto 3);
          Kt_addr                         : out   std_logic_vector(5 downto 0);
          st_cnt_reg                      : out   std_logic_vector(6 to 6);
          Kt_addr_fast                    : out   std_logic_vector(5 downto 0);
          sha256_controller_0_bytes_o     : in    std_logic_vector(1 to 1);
          hash_control_st_reg_ns_i_0_a2_0 : out   std_logic_vector(4 to 4);
          hash_control_st_reg_ns_i_0_a2_2 : in    std_logic_vector(4 to 4);
          hash_control_st_reg_2           : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK    : in    std_logic;
          one_insert                      : out   std_logic;
          sha_last_blk_reg                : out   std_logic;
          SHA256_Module_0_di_req_o        : out   std_logic;
          SHA256_Module_0_do_valid_o      : out   std_logic;
          Kt_addr_2_rep1                  : out   std_logic;
          Kt_addr_2_rep2                  : out   std_logic;
          Kt_addr_1_rep1                  : out   std_logic;
          Kt_addr_1_rep2                  : out   std_logic;
          Kt_addr_3_rep1                  : out   std_logic;
          Kt_addr_3_rep2                  : out   std_logic;
          Kt_addr_5_rep1                  : out   std_logic;
          Kt_addr_0_rep1                  : out   std_logic;
          Kt_addr_0_rep2                  : out   std_logic;
          Kt_addr_4_rep1                  : out   std_logic;
          Kt_addr_4_rep2                  : out   std_logic;
          sha256_controller_0_end_o       : in    std_logic;
          last_block_0                    : in    std_logic;
          N_168_i_0                       : out   std_logic;
          ce_i_i_2                        : in    std_logic;
          pad_one_reg_0_0_a2_0            : out   std_logic;
          sha_last_blk_next_0_o2_0        : out   std_logic;
          oregs_ce_i_a2_0_a2              : out   std_logic;
          N_102                           : out   std_logic;
          N_28                            : in    std_logic;
          N_387                           : out   std_logic;
          N_388                           : in    std_logic;
          W_m4_e_2                        : in    std_logic;
          N_105                           : in    std_logic;
          N_111                           : out   std_logic;
          core_ce_o_iv_i_0                : out   std_logic;
          N_244_i_0                       : out   std_logic;
          SHA256_Module_0_error_o         : out   std_logic;
          ld_i_i_3                        : out   std_logic
        );

end sha256_control;

architecture DEF_ARCH of sha256_control is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \padding_reg\, VCC_net_1, \padding_reg_0_0\, 
        GND_net_1, \hash_control_st_reg_i[6]_net_1\, \one_insert\, 
        \pad_one_reg_0_0\, \msg_bitlen[3]\, 
        un1_msg_bit_cnt_reg_cry_0_Y, \msg_bitlen[4]\, 
        un1_msg_bit_cnt_reg_cry_1_S, \msg_bitlen[5]\, 
        un1_msg_bit_cnt_reg_cry_2_S, \msg_bitlen[6]\, 
        un1_msg_bit_cnt_reg_cry_3_S, \msg_bitlen[7]\, 
        un1_msg_bit_cnt_reg_cry_4_S, \msg_bitlen[8]\, 
        un1_msg_bit_cnt_reg_cry_5_S, \msg_bitlen[9]\, 
        un1_msg_bit_cnt_reg_cry_6_S, \msg_bitlen[10]\, 
        un1_msg_bit_cnt_reg_cry_7_S, \msg_bitlen[11]\, 
        un1_msg_bit_cnt_reg_cry_8_S, \msg_bitlen[12]\, 
        un1_msg_bit_cnt_reg_cry_9_S, \msg_bitlen[13]\, 
        un1_msg_bit_cnt_reg_cry_10_S, \msg_bitlen[14]\, 
        un1_msg_bit_cnt_reg_cry_11_S, \msg_bitlen[15]\, 
        un1_msg_bit_cnt_reg_cry_12_S, \msg_bitlen[16]\, 
        un1_msg_bit_cnt_reg_cry_13_S, \msg_bitlen[17]\, 
        un1_msg_bit_cnt_reg_cry_14_S, \msg_bitlen[18]\, 
        un1_msg_bit_cnt_reg_cry_15_S, \msg_bitlen[19]\, 
        un1_msg_bit_cnt_reg_cry_16_S, \msg_bitlen[20]\, 
        un1_msg_bit_cnt_reg_cry_17_S, \msg_bitlen[21]\, 
        un1_msg_bit_cnt_reg_cry_18_S, \msg_bitlen[22]\, 
        un1_msg_bit_cnt_reg_cry_19_S, \msg_bitlen[23]\, 
        un1_msg_bit_cnt_reg_cry_20_S, \msg_bitlen[24]\, 
        un1_msg_bit_cnt_reg_cry_21_S, \msg_bitlen[25]\, 
        un1_msg_bit_cnt_reg_cry_22_S, \msg_bitlen[26]\, 
        un1_msg_bit_cnt_reg_cry_23_S, \msg_bitlen[27]\, 
        un1_msg_bit_cnt_reg_cry_24_S, \msg_bitlen[28]\, 
        un1_msg_bit_cnt_reg_cry_25_S, \msg_bitlen[29]\, 
        un1_msg_bit_cnt_reg_cry_26_S, \msg_bitlen[30]\, 
        un1_msg_bit_cnt_reg_cry_27_S, \msg_bitlen[31]\, 
        un1_msg_bit_cnt_reg_cry_28_S, \msg_bitlen[32]\, 
        un1_msg_bit_cnt_reg_cry_29_S, \msg_bitlen[33]\, 
        un1_msg_bit_cnt_reg_cry_30_S, \msg_bitlen[34]\, 
        un1_msg_bit_cnt_reg_cry_31_S, \msg_bitlen[35]\, 
        un1_msg_bit_cnt_reg_cry_32_S, \msg_bitlen[36]\, 
        un1_msg_bit_cnt_reg_cry_33_S, \msg_bitlen[37]\, 
        un1_msg_bit_cnt_reg_cry_34_S, \msg_bitlen[38]\, 
        un1_msg_bit_cnt_reg_cry_35_S, \msg_bitlen[39]\, 
        un1_msg_bit_cnt_reg_cry_36_S, \msg_bitlen[40]\, 
        un1_msg_bit_cnt_reg_cry_37_S, \msg_bitlen[41]\, 
        un1_msg_bit_cnt_reg_cry_38_S, \msg_bitlen[42]\, 
        un1_msg_bit_cnt_reg_cry_39_S, \msg_bitlen[43]\, 
        un1_msg_bit_cnt_reg_cry_40_S, \msg_bitlen[44]\, 
        un1_msg_bit_cnt_reg_cry_41_S, \msg_bitlen[45]\, 
        un1_msg_bit_cnt_reg_cry_42_S, \msg_bitlen[46]\, 
        un1_msg_bit_cnt_reg_cry_43_S, \msg_bitlen[47]\, 
        un1_msg_bit_cnt_reg_cry_44_S, \msg_bitlen[48]\, 
        un1_msg_bit_cnt_reg_cry_45_S, \msg_bitlen[49]\, 
        un1_msg_bit_cnt_reg_cry_46_S, \msg_bitlen[50]\, 
        un1_msg_bit_cnt_reg_cry_47_S, \msg_bitlen[51]\, 
        un1_msg_bit_cnt_reg_cry_48_S, \msg_bitlen[52]\, 
        un1_msg_bit_cnt_reg_cry_49_S, \msg_bitlen[53]\, 
        un1_msg_bit_cnt_reg_cry_50_S, \msg_bitlen[54]\, 
        un1_msg_bit_cnt_reg_cry_51_S, \msg_bitlen[55]\, 
        un1_msg_bit_cnt_reg_cry_52_S, \msg_bitlen[56]\, 
        un1_msg_bit_cnt_reg_cry_53_S, \msg_bitlen[57]\, 
        un1_msg_bit_cnt_reg_cry_54_S, \msg_bitlen[58]\, 
        un1_msg_bit_cnt_reg_cry_55_S, \msg_bitlen[59]\, 
        un1_msg_bit_cnt_reg_cry_56_S, \msg_bitlen[60]\, 
        un1_msg_bit_cnt_reg_cry_57_S, \msg_bitlen[61]\, 
        un1_msg_bit_cnt_reg_cry_58_S, \msg_bitlen[62]\, 
        un1_msg_bit_cnt_reg_cry_59_S, \msg_bitlen[63]\, 
        un1_msg_bit_cnt_reg_s_60_S, 
        \hash_control_st_reg_nsss_i_0[0]\, sha_last_blk_reg_net_1, 
        \sha_last_blk_reg_RNO\, \sha_last_blk_regce\, 
        \Kt_addr[0]\, \st_cnt_reg_s[0]\, st_cnt_rege, 
        \Kt_addr[1]\, \st_cnt_reg_s[1]\, \Kt_addr[2]\, 
        \st_cnt_reg_s[2]\, \Kt_addr[3]\, \st_cnt_reg_s[3]\, 
        \Kt_addr[4]\, \st_cnt_reg_s[4]\, \Kt_addr[5]\, 
        \st_cnt_reg_s[5]\, \st_cnt_reg[6]_net_1\, 
        \st_cnt_reg_s[6]_net_1\, \SHA256_Module_0_di_req_o\, 
        hash_control_st_reg_4, \hash_control_st_reg[0]_net_1\, 
        hash_control_st_reg_3, \SHA256_Module_0_do_valid_o\, 
        hash_control_st_reg_2_0, \hash_control_st_reg_2\, 
        hash_control_st_reg_1, \hash_control_st_reg[3]_net_1\, 
        hash_control_st_reg_0, \hash_control_st_reg[4]_net_1\, 
        hash_control_st_reg, \Kt_addr_fast[2]\, \Kt_addr_fast[1]\, 
        \Kt_addr_fast[3]\, \Kt_addr_0_rep2\, st_cnt_reg_cry_cy, 
        st_cnt_clr, \st_cnt_reg_cry[0]_net_1\, 
        \st_cnt_reg_cry[1]_net_1\, \st_cnt_reg_cry[2]_net_1\, 
        \st_cnt_reg_cry[3]_net_1\, \st_cnt_reg_cry[4]_net_1\, 
        \st_cnt_reg_cry[5]_net_1\, \un1_msg_bit_cnt_reg_cry_0\, 
        N_229, \un1_msg_bit_cnt_reg_cry_1\, 
        \un1_msg_bit_cnt_reg_cry_2\, \un1_msg_bit_cnt_reg_cry_3\, 
        \un1_msg_bit_cnt_reg_cry_4\, \un1_msg_bit_cnt_reg_cry_5\, 
        \un1_msg_bit_cnt_reg_cry_6\, \un1_msg_bit_cnt_reg_cry_7\, 
        \un1_msg_bit_cnt_reg_cry_8\, \un1_msg_bit_cnt_reg_cry_9\, 
        \un1_msg_bit_cnt_reg_cry_10\, 
        \un1_msg_bit_cnt_reg_cry_11\, 
        \un1_msg_bit_cnt_reg_cry_12\, 
        \un1_msg_bit_cnt_reg_cry_13\, 
        \un1_msg_bit_cnt_reg_cry_14\, 
        \un1_msg_bit_cnt_reg_cry_15\, 
        \un1_msg_bit_cnt_reg_cry_16\, 
        \un1_msg_bit_cnt_reg_cry_17\, 
        \un1_msg_bit_cnt_reg_cry_18\, 
        \un1_msg_bit_cnt_reg_cry_19\, 
        \un1_msg_bit_cnt_reg_cry_20\, 
        \un1_msg_bit_cnt_reg_cry_21\, 
        \un1_msg_bit_cnt_reg_cry_22\, 
        \un1_msg_bit_cnt_reg_cry_23\, 
        \un1_msg_bit_cnt_reg_cry_24\, 
        \un1_msg_bit_cnt_reg_cry_25\, 
        \un1_msg_bit_cnt_reg_cry_26\, 
        \un1_msg_bit_cnt_reg_cry_27\, 
        \un1_msg_bit_cnt_reg_cry_28\, 
        \un1_msg_bit_cnt_reg_cry_29\, 
        \un1_msg_bit_cnt_reg_cry_30\, 
        \un1_msg_bit_cnt_reg_cry_31\, 
        \un1_msg_bit_cnt_reg_cry_32\, 
        \un1_msg_bit_cnt_reg_cry_33\, 
        \un1_msg_bit_cnt_reg_cry_34\, 
        \un1_msg_bit_cnt_reg_cry_35\, 
        \un1_msg_bit_cnt_reg_cry_36\, 
        \un1_msg_bit_cnt_reg_cry_37\, 
        \un1_msg_bit_cnt_reg_cry_38\, 
        \un1_msg_bit_cnt_reg_cry_39\, 
        \un1_msg_bit_cnt_reg_cry_40\, 
        \un1_msg_bit_cnt_reg_cry_41\, 
        \un1_msg_bit_cnt_reg_cry_42\, 
        \un1_msg_bit_cnt_reg_cry_43\, 
        \un1_msg_bit_cnt_reg_cry_44\, 
        \un1_msg_bit_cnt_reg_cry_45\, 
        \un1_msg_bit_cnt_reg_cry_46\, 
        \un1_msg_bit_cnt_reg_cry_47\, 
        \un1_msg_bit_cnt_reg_cry_48\, 
        \un1_msg_bit_cnt_reg_cry_49\, 
        \un1_msg_bit_cnt_reg_cry_50\, 
        \un1_msg_bit_cnt_reg_cry_51\, 
        \un1_msg_bit_cnt_reg_cry_52\, 
        \un1_msg_bit_cnt_reg_cry_53\, 
        \un1_msg_bit_cnt_reg_cry_54\, 
        \un1_msg_bit_cnt_reg_cry_55\, 
        \un1_msg_bit_cnt_reg_cry_56\, 
        \un1_msg_bit_cnt_reg_cry_57\, 
        \un1_msg_bit_cnt_reg_cry_58\, 
        \un1_msg_bit_cnt_reg_cry_59\, N_389, N_228, 
        \hash_control_st_reg_r_1[4]_net_1\, 
        \hash_control_st_reg_ns_0_0_a4_1_2[2]_net_1\, N_373, 
        N_104, N_115, \sha_last_blk_next_0_a4_1\, 
        \pad_one_reg_0_0_o2_0\, \sha_last_blk_next_0_o2_0\, 
        oregs_ce_i_a2_0_a2_net_1, N_119, N_233, N_149, N_398, 
        \hash_control_st_reg_ns_i_0_a4_1_1[4]_net_1\, 
        \hash_control_st_reg_ns_0_0_a4_0_0[6]_net_1\, \N_102\, 
        N_399, N_363, N_402, N_217, N_391, \N_387\, 
        \hash_control_st_reg_ns_i_0_0[4]_net_1\, 
        \pad_one_reg_0_0_a4_1_1\, N_368, N_340, N_357, N_338, 
        N_341, N_375, \hash_control_st_reg_ns_i_0_0[1]_net_1\, 
        N_367, N_355, \N_111\, N_118, 
        \hash_control_st_reg_ns_i_0_1[1]_net_1\, N_358
         : std_logic;

begin 

    hash_control_st_reg_i(6) <= \hash_control_st_reg_i[6]_net_1\;
    msg_bitlen(63) <= \msg_bitlen[63]\;
    msg_bitlen(62) <= \msg_bitlen[62]\;
    msg_bitlen(61) <= \msg_bitlen[61]\;
    msg_bitlen(60) <= \msg_bitlen[60]\;
    msg_bitlen(59) <= \msg_bitlen[59]\;
    msg_bitlen(58) <= \msg_bitlen[58]\;
    msg_bitlen(57) <= \msg_bitlen[57]\;
    msg_bitlen(56) <= \msg_bitlen[56]\;
    msg_bitlen(55) <= \msg_bitlen[55]\;
    msg_bitlen(54) <= \msg_bitlen[54]\;
    msg_bitlen(53) <= \msg_bitlen[53]\;
    msg_bitlen(52) <= \msg_bitlen[52]\;
    msg_bitlen(51) <= \msg_bitlen[51]\;
    msg_bitlen(50) <= \msg_bitlen[50]\;
    msg_bitlen(49) <= \msg_bitlen[49]\;
    msg_bitlen(48) <= \msg_bitlen[48]\;
    msg_bitlen(47) <= \msg_bitlen[47]\;
    msg_bitlen(46) <= \msg_bitlen[46]\;
    msg_bitlen(45) <= \msg_bitlen[45]\;
    msg_bitlen(44) <= \msg_bitlen[44]\;
    msg_bitlen(43) <= \msg_bitlen[43]\;
    msg_bitlen(42) <= \msg_bitlen[42]\;
    msg_bitlen(41) <= \msg_bitlen[41]\;
    msg_bitlen(40) <= \msg_bitlen[40]\;
    msg_bitlen(39) <= \msg_bitlen[39]\;
    msg_bitlen(38) <= \msg_bitlen[38]\;
    msg_bitlen(37) <= \msg_bitlen[37]\;
    msg_bitlen(36) <= \msg_bitlen[36]\;
    msg_bitlen(35) <= \msg_bitlen[35]\;
    msg_bitlen(34) <= \msg_bitlen[34]\;
    msg_bitlen(33) <= \msg_bitlen[33]\;
    msg_bitlen(32) <= \msg_bitlen[32]\;
    msg_bitlen(31) <= \msg_bitlen[31]\;
    msg_bitlen(30) <= \msg_bitlen[30]\;
    msg_bitlen(29) <= \msg_bitlen[29]\;
    msg_bitlen(28) <= \msg_bitlen[28]\;
    msg_bitlen(27) <= \msg_bitlen[27]\;
    msg_bitlen(26) <= \msg_bitlen[26]\;
    msg_bitlen(25) <= \msg_bitlen[25]\;
    msg_bitlen(24) <= \msg_bitlen[24]\;
    msg_bitlen(23) <= \msg_bitlen[23]\;
    msg_bitlen(22) <= \msg_bitlen[22]\;
    msg_bitlen(21) <= \msg_bitlen[21]\;
    msg_bitlen(20) <= \msg_bitlen[20]\;
    msg_bitlen(19) <= \msg_bitlen[19]\;
    msg_bitlen(18) <= \msg_bitlen[18]\;
    msg_bitlen(17) <= \msg_bitlen[17]\;
    msg_bitlen(16) <= \msg_bitlen[16]\;
    msg_bitlen(15) <= \msg_bitlen[15]\;
    msg_bitlen(14) <= \msg_bitlen[14]\;
    msg_bitlen(13) <= \msg_bitlen[13]\;
    msg_bitlen(12) <= \msg_bitlen[12]\;
    msg_bitlen(11) <= \msg_bitlen[11]\;
    msg_bitlen(10) <= \msg_bitlen[10]\;
    msg_bitlen(9) <= \msg_bitlen[9]\;
    msg_bitlen(8) <= \msg_bitlen[8]\;
    msg_bitlen(7) <= \msg_bitlen[7]\;
    msg_bitlen(6) <= \msg_bitlen[6]\;
    msg_bitlen(5) <= \msg_bitlen[5]\;
    msg_bitlen(4) <= \msg_bitlen[4]\;
    msg_bitlen(3) <= \msg_bitlen[3]\;
    Kt_addr(5) <= \Kt_addr[5]\;
    Kt_addr(4) <= \Kt_addr[4]\;
    Kt_addr(3) <= \Kt_addr[3]\;
    Kt_addr(2) <= \Kt_addr[2]\;
    Kt_addr(1) <= \Kt_addr[1]\;
    Kt_addr(0) <= \Kt_addr[0]\;
    st_cnt_reg(6) <= \st_cnt_reg[6]_net_1\;
    Kt_addr_fast(3) <= \Kt_addr_fast[3]\;
    Kt_addr_fast(2) <= \Kt_addr_fast[2]\;
    Kt_addr_fast(1) <= \Kt_addr_fast[1]\;
    hash_control_st_reg_2 <= \hash_control_st_reg_2\;
    one_insert <= \one_insert\;
    sha_last_blk_reg <= sha_last_blk_reg_net_1;
    SHA256_Module_0_di_req_o <= \SHA256_Module_0_di_req_o\;
    SHA256_Module_0_do_valid_o <= \SHA256_Module_0_do_valid_o\;
    Kt_addr_0_rep2 <= \Kt_addr_0_rep2\;
    sha_last_blk_next_0_o2_0 <= \sha_last_blk_next_0_o2_0\;
    oregs_ce_i_a2_0_a2 <= oregs_ce_i_a2_0_a2_net_1;
    N_102 <= \N_102\;
    N_387 <= \N_387\;
    N_111 <= \N_111\;

    pad_one_reg_0_0_a4_1_1 : CFG3
      generic map(INIT => x"80")

      port map(A => \hash_control_st_reg_i[6]_net_1\, B => N_399, 
        C => N_388, Y => \pad_one_reg_0_0_a4_1_1\);
    
    \msg_bit_cnt_reg[42]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_39_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[42]\);
    
    \hash_control_st_reg_r[3]\ : CFG4
      generic map(INIT => x"4454")

      port map(A => last_block_0, B => N_363, C => N_389, D => 
        N_228, Y => hash_control_st_reg_0);
    
    un1_msg_bit_cnt_reg_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[17]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_13\, S => 
        un1_msg_bit_cnt_reg_cry_14_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_14\);
    
    un1_msg_bit_cnt_reg_cry_18 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[21]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_17\, S => 
        un1_msg_bit_cnt_reg_cry_18_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_18\);
    
    un1_msg_bit_cnt_reg_cry_16 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[19]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_15\, S => 
        un1_msg_bit_cnt_reg_cry_16_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_16\);
    
    un1_msg_bit_cnt_reg_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[14]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_10\, S => 
        un1_msg_bit_cnt_reg_cry_11_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_11\);
    
    \msg_bit_cnt_reg[35]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_32_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[35]\);
    
    \hash_control_st_reg_ns_i_0_o2[4]\ : CFG4
      generic map(INIT => x"C0AA")

      port map(A => N_399, B => 
        hash_control_st_reg_ns_i_0_a2_2(4), C => \Kt_addr[3]\, D
         => \Kt_addr[0]\, Y => N_118);
    
    sha_last_blk_regce : CFG4
      generic map(INIT => x"0BBB")

      port map(A => N_338, B => \N_111\, C => ce_i_i_2, D => 
        \hash_control_st_reg_i[6]_net_1\, Y => 
        \sha_last_blk_regce\);
    
    un1_msg_bit_cnt_reg_cry_20 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[23]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_19\, S => 
        un1_msg_bit_cnt_reg_cry_20_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_20\);
    
    \msg_bit_cnt_reg[63]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_s_60_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[63]\);
    
    \pad_one_reg_0_0_a2_0\ : CFG3
      generic map(INIT => x"70")

      port map(A => sha256_controller_0_bytes_o(1), B => 
        sha256_controller_0_end_o, C => 
        \SHA256_Module_0_di_req_o\, Y => \N_387\);
    
    \msg_bit_cnt_reg[48]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_45_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[48]\);
    
    st_cnt_reg_1_rep2 : SLE
      port map(D => \st_cnt_reg_s[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_1_rep2);
    
    \msg_bit_cnt_reg[39]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_36_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[39]\);
    
    sch_ld_o_i_0_0 : CFG4
      generic map(INIT => x"DCCC")

      port map(A => \Kt_addr[0]\, B => 
        \hash_control_st_reg[4]_net_1\, C => N_399, D => N_402, Y
         => ld_i_i_3);
    
    st_cnt_reg_0_rep2 : SLE
      port map(D => \st_cnt_reg_s[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \Kt_addr_0_rep2\);
    
    \hash_control_st_reg_ns_i_0_0[1]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => ce_i_i_2, B => \SHA256_Module_0_di_req_o\, C
         => \hash_control_st_reg_i[6]_net_1\, D => N_217, Y => 
        \hash_control_st_reg_ns_i_0_0[1]_net_1\);
    
    un1_msg_bit_cnt_reg_cry_49 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[52]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_48\, S => 
        un1_msg_bit_cnt_reg_cry_49_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_49\);
    
    \st_cnt_reg_cry_cy[0]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => st_cnt_clr, C => GND_net_1, D
         => GND_net_1, FCI => VCC_net_1, S => OPEN, Y => OPEN, 
        FCO => st_cnt_reg_cry_cy);
    
    un1_msg_bit_cnt_reg_cry_57 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[60]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_56\, S => 
        un1_msg_bit_cnt_reg_cry_57_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_57\);
    
    un1_msg_bit_cnt_reg_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_3\, S => 
        un1_msg_bit_cnt_reg_cry_4_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_4\);
    
    st_cnt_reg_4_rep1 : SLE
      port map(D => \st_cnt_reg_s[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_4_rep1);
    
    \msg_bit_cnt_reg[34]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_31_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[34]\);
    
    \hash_control_st_reg_ns_0_0_a4_0_0[6]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \SHA256_Module_0_do_valid_o\, B => 
        \SHA256_Module_0_di_req_o\, C => N_398, Y => 
        \hash_control_st_reg_ns_0_0_a4_0_0[6]_net_1\);
    
    pad_one_reg_0_0_a2 : CFG4
      generic map(INIT => x"0004")

      port map(A => \Kt_addr[1]\, B => \Kt_addr[4]\, C => 
        \Kt_addr[3]\, D => \Kt_addr[2]\, Y => N_399);
    
    \msg_bit_cnt_reg[4]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_1_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[4]\);
    
    sha_last_blk_next_0_a4_1 : CFG2
      generic map(INIT => x"2")

      port map(A => \Kt_addr[0]\, B => \Kt_addr[4]\, Y => 
        \sha_last_blk_next_0_a4_1\);
    
    \hash_control_st_reg_ns_0_0_a4_0[2]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => N_402, B => N_118, C => ce_i_i_2, D => N_28, 
        Y => N_373);
    
    \hash_control_st_reg[0]\ : SLE
      port map(D => hash_control_st_reg_3, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \hash_control_st_reg[0]_net_1\);
    
    \st_cnt_reg_fast[4]\ : SLE
      port map(D => \st_cnt_reg_s[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_fast(4));
    
    un1_msg_bit_cnt_reg_cry_45 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[48]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_44\, S => 
        un1_msg_bit_cnt_reg_cry_45_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_45\);
    
    sch_ld_o_i_0_0_a2_0 : CFG3
      generic map(INIT => x"02")

      port map(A => \hash_control_st_reg_2\, B => \Kt_addr[5]\, C
         => \st_cnt_reg[6]_net_1\, Y => N_402);
    
    \hash_control_st_reg_r_1[4]\ : CFG4
      generic map(INIT => x"3331")

      port map(A => \hash_control_st_reg_ns_0_0_a4_1_2[2]_net_1\, 
        B => N_373, C => N_104, D => N_115, Y => 
        \hash_control_st_reg_r_1[4]_net_1\);
    
    \msg_bit_cnt_reg[23]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_20_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[23]\);
    
    un1_msg_bit_cnt_reg_cry_23 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[26]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_22\, S => 
        un1_msg_bit_cnt_reg_cry_23_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_23\);
    
    \state_counter_proc.un15_ce_i_i_0_a2_RNIKNCQ\ : CFG2
      generic map(INIT => x"7")

      port map(A => N_115, B => N_398, Y => N_244_i_0);
    
    \msg_bit_cnt_reg[10]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_7_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[10]\);
    
    \hash_control_st_reg[3]\ : SLE
      port map(D => hash_control_st_reg_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \hash_control_st_reg[3]_net_1\);
    
    \hash_control_st_reg_nsss_i[0]\ : CFG3
      generic map(INIT => x"51")

      port map(A => last_block_0, B => ce_i_i_2, C => 
        \hash_control_st_reg_i[6]_net_1\, Y => 
        \hash_control_st_reg_nsss_i_0[0]\);
    
    \st_cnt_reg[2]\ : SLE
      port map(D => \st_cnt_reg_s[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \Kt_addr[2]\);
    
    st_cnt_reg_2_rep2 : SLE
      port map(D => \st_cnt_reg_s[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_2_rep2);
    
    un1_msg_bit_cnt_reg_cry_44 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[47]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_43\, S => 
        un1_msg_bit_cnt_reg_cry_44_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_44\);
    
    un1_msg_bit_cnt_reg_cry_48 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[51]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_47\, S => 
        un1_msg_bit_cnt_reg_cry_48_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_48\);
    
    un1_msg_bit_cnt_reg_cry_46 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[49]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_45\, S => 
        un1_msg_bit_cnt_reg_cry_46_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_46\);
    
    un1_msg_bit_cnt_reg_cry_37 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[40]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_36\, S => 
        un1_msg_bit_cnt_reg_cry_37_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_37\);
    
    un1_msg_bit_cnt_reg_cry_41 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[44]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_40\, S => 
        un1_msg_bit_cnt_reg_cry_41_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_41\);
    
    \msg_bit_cnt_reg[11]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_8_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[11]\);
    
    un1_msg_bit_cnt_reg_s_60 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[63]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_59\, S => 
        un1_msg_bit_cnt_reg_s_60_S, Y => OPEN, FCO => OPEN);
    
    \msg_bit_cnt_reg[40]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_37_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[40]\);
    
    \st_cnt_reg_fast[0]\ : SLE
      port map(D => \st_cnt_reg_s[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_fast(0));
    
    \msg_bit_cnt_reg[52]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_49_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[52]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un1_msg_bit_cnt_reg_cry_29 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[32]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_28\, S => 
        un1_msg_bit_cnt_reg_cry_29_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_29\);
    
    \st_cnt_reg_cry[4]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[4]\, 
        D => GND_net_1, FCI => \st_cnt_reg_cry[3]_net_1\, S => 
        \st_cnt_reg_s[4]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[4]_net_1\);
    
    un1_msg_bit_cnt_reg_cry_2 : ARI1
      generic map(INIT => x"5EA15")

      port map(A => \msg_bitlen[5]\, B => N_229, C => 
        sha256_controller_0_bytes_o(1), D => 
        sha256_controller_0_end_o, FCI => 
        \un1_msg_bit_cnt_reg_cry_1\, S => 
        un1_msg_bit_cnt_reg_cry_2_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_2\);
    
    \hash_control_st_reg_ns_i_0_a2_0[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \Kt_addr_fast[1]\, B => \Kt_addr_fast[2]\, Y
         => hash_control_st_reg_ns_i_0_a2_0(4));
    
    \msg_bit_cnt_reg[41]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_38_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[41]\);
    
    \msg_bit_cnt_reg[58]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_55_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[58]\);
    
    \st_cnt_reg[3]\ : SLE
      port map(D => \st_cnt_reg_s[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \Kt_addr[3]\);
    
    \st_cnt_reg_fast[3]\ : SLE
      port map(D => \st_cnt_reg_s[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \Kt_addr_fast[3]\);
    
    \msg_bit_cnt_reg[27]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_24_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[27]\);
    
    un1_msg_bit_cnt_reg_cry_25 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[28]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_24\, S => 
        un1_msg_bit_cnt_reg_cry_25_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_25\);
    
    \msg_bit_cnt_reg[26]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_23_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[26]\);
    
    \msg_bit_cnt_reg[3]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_0_Y, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[3]\);
    
    st_cnt_clr_0_a2_0_a4 : CFG3
      generic map(INIT => x"10")

      port map(A => \SHA256_Module_0_do_valid_o\, B => 
        \SHA256_Module_0_di_req_o\, C => N_398, Y => st_cnt_clr);
    
    \hash_control_st_reg_ns_0_0_a4_1_2[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => sha256_controller_0_bytes_o(1), B => 
        sha256_controller_0_end_o, C => \Kt_addr[5]\, D => N_149, 
        Y => \hash_control_st_reg_ns_0_0_a4_1_2[2]_net_1\);
    
    un1_msg_bit_cnt_reg_cry_24 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[27]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_23\, S => 
        un1_msg_bit_cnt_reg_cry_24_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_24\);
    
    un1_msg_bit_cnt_reg_cry_28 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[31]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_27\, S => 
        un1_msg_bit_cnt_reg_cry_28_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_28\);
    
    un1_msg_bit_cnt_reg_cry_26 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[29]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_25\, S => 
        un1_msg_bit_cnt_reg_cry_26_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_26\);
    
    \state_counter_proc.un15_ce_i_i_0_o2\ : CFG2
      generic map(INIT => x"7")

      port map(A => N_28, B => \SHA256_Module_0_di_req_o\, Y => 
        N_115);
    
    un1_msg_bit_cnt_reg_cry_21 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[24]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_20\, S => 
        un1_msg_bit_cnt_reg_cry_21_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_21\);
    
    \msg_bit_cnt_reg[6]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_3_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[6]\);
    
    un1_msg_bit_cnt_reg_cry_17 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[20]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_16\, S => 
        un1_msg_bit_cnt_reg_cry_17_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_17\);
    
    \st_cnt_reg_s[6]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => 
        \st_cnt_reg[6]_net_1\, D => GND_net_1, FCI => 
        \st_cnt_reg_cry[5]_net_1\, S => \st_cnt_reg_s[6]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    un1_msg_bit_cnt_reg_cry_52 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[55]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_51\, S => 
        un1_msg_bit_cnt_reg_cry_52_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_52\);
    
    \hash_control_st_reg_ns_i_0_o2_1[4]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \SHA256_Module_0_di_req_o\, B => 
        sha256_controller_0_end_o, Y => N_233);
    
    \msg_bit_cnt_reg[32]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_29_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[32]\);
    
    \msg_bit_cnt_reg[25]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_22_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[25]\);
    
    \hash_control_st_reg_ns_i_0_o2_1[1]\ : CFG2
      generic map(INIT => x"B")

      port map(A => sha_last_blk_reg_net_1, B => 
        \hash_control_st_reg[3]_net_1\, Y => N_119);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    st_cnt_reg_3_rep2 : SLE
      port map(D => \st_cnt_reg_s[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_3_rep2);
    
    sha_last_blk_next_0_o2_0_1 : CFG2
      generic map(INIT => x"E")

      port map(A => \Kt_addr_0_rep2\, B => \one_insert\, Y => 
        \sha_last_blk_next_0_o2_0\);
    
    un1_msg_bit_cnt_reg_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_5\, S => 
        un1_msg_bit_cnt_reg_cry_6_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_6\);
    
    un1_msg_bit_cnt_reg_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_7\, S => 
        un1_msg_bit_cnt_reg_cry_8_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_8\);
    
    \st_cnt_reg_fast[1]\ : SLE
      port map(D => \st_cnt_reg_s[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \Kt_addr_fast[1]\);
    
    \msg_bit_cnt_reg[50]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_47_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[50]\);
    
    \msg_bit_cnt_reg[29]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_26_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[29]\);
    
    \st_cnt_reg_cry[2]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[2]\, 
        D => GND_net_1, FCI => \st_cnt_reg_cry[1]_net_1\, S => 
        \st_cnt_reg_s[2]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[2]_net_1\);
    
    \st_cnt_reg[5]\ : SLE
      port map(D => \st_cnt_reg_s[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \Kt_addr[5]\);
    
    \msg_bit_cnt_reg[38]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_35_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[38]\);
    
    \hash_control_st_reg_ns_i_0_a4_1[4]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \hash_control_st_reg_ns_i_0_a4_1_1[4]_net_1\, 
        B => ce_i_i_2, C => N_118, D => N_28, Y => N_358);
    
    \hash_control_st_reg_ns_0_0_a2[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_28, B => \hash_control_st_reg[4]_net_1\, Y
         => N_389);
    
    \msg_bit_cnt_reg[13]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_10_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[13]\);
    
    \st_cnt_reg[6]\ : SLE
      port map(D => \st_cnt_reg_s[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \st_cnt_reg[6]_net_1\);
    
    \hash_control_st_reg_ns_i_0_a4_1_1[4]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \hash_control_st_reg[3]_net_1\, B => 
        \Kt_addr[5]\, C => \st_cnt_reg[6]_net_1\, Y => 
        \hash_control_st_reg_ns_i_0_a4_1_1[4]_net_1\);
    
    \msg_bit_cnt_reg[51]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_48_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[51]\);
    
    \msg_bit_cnt_reg[24]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_21_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[24]\);
    
    pad_one_reg_0_0 : CFG4
      generic map(INIT => x"FEEE")

      port map(A => N_367, B => N_368, C => N_402, D => 
        \pad_one_reg_0_0_a4_1_1\, Y => \pad_one_reg_0_0\);
    
    \hash_control_st_reg[4]\ : SLE
      port map(D => hash_control_st_reg, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \hash_control_st_reg[4]_net_1\);
    
    \hash_control_st_reg_ns_0_0_o2_0[2]\ : CFG4
      generic map(INIT => x"F7FF")

      port map(A => \Kt_addr_fast[2]\, B => \Kt_addr_fast[1]\, C
         => \st_cnt_reg[6]_net_1\, D => \Kt_addr_fast[3]\, Y => 
        \N_102\);
    
    un1_msg_bit_cnt_reg_cry_32 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[35]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_31\, S => 
        un1_msg_bit_cnt_reg_cry_32_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_32\);
    
    \hash_control_st_reg_ns_i_0_o2[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_119, B => \padding_reg\, Y => N_217);
    
    \hash_control_st_reg_ns_i_0_0[4]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => \hash_control_st_reg_2\, B => ce_i_i_2, C => 
        N_28, D => N_233, Y => 
        \hash_control_st_reg_ns_i_0_0[4]_net_1\);
    
    \st_cnt_reg_cry[0]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[0]\, 
        D => GND_net_1, FCI => st_cnt_reg_cry_cy, S => 
        \st_cnt_reg_s[0]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[0]_net_1\);
    
    \msg_bit_cnt_reg[43]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_40_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[43]\);
    
    \hash_control_st_reg[2]\ : SLE
      port map(D => hash_control_st_reg_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \hash_control_st_reg_2\);
    
    \hash_control_st_reg_ns_i_0_1[1]\ : CFG4
      generic map(INIT => x"FF20")

      port map(A => sha256_controller_0_end_o, B => ce_i_i_2, C
         => N_391, D => \hash_control_st_reg_ns_i_0_0[1]_net_1\, 
        Y => \hash_control_st_reg_ns_i_0_1[1]_net_1\);
    
    un1_msg_bit_cnt_reg_cry_47 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[50]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_46\, S => 
        un1_msg_bit_cnt_reg_cry_47_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_47\);
    
    un1_msg_bit_cnt_reg_cry_0 : ARI1
      generic map(INIT => x"5BF40")

      port map(A => \msg_bitlen[3]\, B => N_229, C => 
        sha256_controller_0_bytes_o(1), D => 
        sha256_controller_0_end_o, FCI => GND_net_1, S => OPEN, Y
         => un1_msg_bit_cnt_reg_cry_0_Y, FCO => 
        \un1_msg_bit_cnt_reg_cry_0\);
    
    \st_cnt_reg[1]\ : SLE
      port map(D => \st_cnt_reg_s[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \Kt_addr[1]\);
    
    sha_last_blk_reg_RNO : CFG2
      generic map(INIT => x"B")

      port map(A => \sha_last_blk_regce\, B => 
        \hash_control_st_reg_i[6]_net_1\, Y => 
        \sha_last_blk_reg_RNO\);
    
    un1_msg_bit_cnt_reg_cry_50 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[53]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_49\, S => 
        un1_msg_bit_cnt_reg_cry_50_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_50\);
    
    \hash_control_st_reg_ns_0_0_o2[2]\ : CFG4
      generic map(INIT => x"FFF7")

      port map(A => \Kt_addr[4]\, B => \Kt_addr[5]\, C => N_149, 
        D => \N_102\, Y => N_228);
    
    pad_one_reg : SLE
      port map(D => \pad_one_reg_0_0\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => VCC_net_1, LAT
         => GND_net_1, Q => \one_insert\);
    
    \hash_control_st_reg_ns_0_0_a4[6]\ : CFG4
      generic map(INIT => x"44C4")

      port map(A => \SHA256_Module_0_di_req_o\, B => N_391, C => 
        sha256_controller_0_bytes_o(1), D => 
        sha256_controller_0_end_o, Y => N_341);
    
    \hash_control_st_reg_ns_0_0_a4_0[5]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => ce_i_i_2, B => N_28, C => 
        \hash_control_st_reg[3]_net_1\, D => 
        sha_last_blk_reg_net_1, Y => N_340);
    
    \msg_bit_cnt_reg[17]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_14_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[17]\);
    
    \msg_bit_cnt_reg[16]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_13_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[16]\);
    
    un1_msg_bit_cnt_reg_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_8\, S => 
        un1_msg_bit_cnt_reg_cry_9_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_9\);
    
    \msg_bit_cnt_reg[30]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_27_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[30]\);
    
    sha_last_blk_next_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => N_105, B => \sha_last_blk_next_0_o2_0\, Y => 
        \N_111\);
    
    st_cnt_reg_4_rep2 : SLE
      port map(D => \st_cnt_reg_s[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_4_rep2);
    
    oregs_ce_i_a2_0_a2_i : CFG2
      generic map(INIT => x"D")

      port map(A => \hash_control_st_reg_i[6]_net_1\, B => 
        \hash_control_st_reg[3]_net_1\, Y => N_168_i_0);
    
    \hash_control_st_reg[1]\ : SLE
      port map(D => hash_control_st_reg_2_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_Module_0_do_valid_o\);
    
    \hash_control_st_reg_r[0]\ : CFG4
      generic map(INIT => x"3230")

      port map(A => \hash_control_st_reg_ns_0_0_a4_0_0[6]_net_1\, 
        B => last_block_0, C => N_341, D => 
        oregs_ce_i_a2_0_a2_net_1, Y => hash_control_st_reg_3);
    
    \msg_bit_cnt_reg[31]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_28_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[31]\);
    
    \hash_control_st_reg_RNI42JO1[0]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => \SHA256_Module_0_do_valid_o\, B => 
        \hash_control_st_reg[0]_net_1\, C => N_28, D => 
        \SHA256_Module_0_di_req_o\, Y => core_ce_o_iv_i_0);
    
    \un1_ce_i_i_o4[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_115, B => ce_i_i_2, Y => N_229);
    
    st_cnt_reg_1_rep1 : SLE
      port map(D => \st_cnt_reg_s[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_1_rep1);
    
    \msg_bit_cnt_reg[47]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_44_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[47]\);
    
    \st_cnt_reg[4]\ : SLE
      port map(D => \st_cnt_reg_s[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \Kt_addr[4]\);
    
    \sha_last_blk_reg\ : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => 
        \sha_last_blk_reg_RNO\, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => \hash_control_st_reg_i[6]_net_1\, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        sha_last_blk_reg_net_1);
    
    pad_one_reg_0_0_o2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => ce_i_i_2, B => \hash_control_st_reg[4]_net_1\, 
        Y => \pad_one_reg_0_0_o2_0\);
    
    \st_cnt_reg_cry[1]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[1]\, 
        D => GND_net_1, FCI => \st_cnt_reg_cry[0]_net_1\, S => 
        \st_cnt_reg_s[1]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[1]_net_1\);
    
    un1_msg_bit_cnt_reg_cry_30 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[33]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_29\, S => 
        un1_msg_bit_cnt_reg_cry_30_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_30\);
    
    \msg_bit_cnt_reg[46]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_43_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[46]\);
    
    st_cnt_reg_0_rep1 : SLE
      port map(D => \st_cnt_reg_s[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_0_rep1);
    
    \msg_bit_cnt_reg[62]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_59_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[62]\);
    
    un1_msg_bit_cnt_reg_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[15]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_11\, S => 
        un1_msg_bit_cnt_reg_cry_12_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_12\);
    
    \hash_control_st_reg_ns_i_0_o2_0[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \N_102\, B => \Kt_addr[4]\, Y => N_104);
    
    un1_msg_bit_cnt_reg_cry_53 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[56]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_52\, S => 
        un1_msg_bit_cnt_reg_cry_53_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_53\);
    
    padding_reg : SLE
      port map(D => \padding_reg_0_0\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \padding_reg\);
    
    sha_last_blk_next_0_a4 : CFG4
      generic map(INIT => x"4000")

      port map(A => \Kt_addr[1]\, B => \Kt_addr[3]\, C => 
        W_m4_e_2, D => \sha_last_blk_next_0_a4_1\, Y => N_338);
    
    un1_msg_bit_cnt_reg_cry_27 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[30]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_26\, S => 
        un1_msg_bit_cnt_reg_cry_27_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_27\);
    
    \msg_bit_cnt_reg[15]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_12_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[15]\);
    
    \hash_control_st_reg_ns_i_0_a4_2[1]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \Kt_addr[5]\, B => N_149, C => N_104, D => 
        N_391, Y => N_355);
    
    \st_cnt_reg_cry[3]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[3]\, 
        D => GND_net_1, FCI => \st_cnt_reg_cry[2]_net_1\, S => 
        \st_cnt_reg_s[3]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[3]_net_1\);
    
    \msg_bit_cnt_reg[53]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_50_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[53]\);
    
    \msg_bit_cnt_reg[19]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_16_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[19]\);
    
    \hash_control_st_reg_r[1]\ : CFG4
      generic map(INIT => x"5504")

      port map(A => last_block_0, B => 
        \SHA256_Module_0_do_valid_o\, C => N_28, D => N_340, Y
         => hash_control_st_reg_2_0);
    
    \st_cnt_reg_fast[2]\ : SLE
      port map(D => \st_cnt_reg_s[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \Kt_addr_fast[2]\);
    
    un1_msg_bit_cnt_reg_cry_59 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[62]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_58\, S => 
        un1_msg_bit_cnt_reg_cry_59_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_59\);
    
    \msg_bit_cnt_reg[45]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_42_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[45]\);
    
    \msg_bit_cnt_reg[22]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_19_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[22]\);
    
    \hash_control_st_reg_r[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => N_357, B => last_block_0, C => N_358, D => 
        \hash_control_st_reg_ns_i_0_0[4]_net_1\, Y => 
        hash_control_st_reg_1);
    
    st_cnt_reg_2_rep1 : SLE
      port map(D => \st_cnt_reg_s[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_2_rep1);
    
    un1_msg_bit_cnt_reg_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_4\, S => 
        un1_msg_bit_cnt_reg_cry_5_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_5\);
    
    un1_msg_bit_cnt_reg_cry_33 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[36]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_32\, S => 
        un1_msg_bit_cnt_reg_cry_33_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_33\);
    
    \msg_bit_cnt_reg[14]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_11_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[14]\);
    
    \state_counter_proc.un15_ce_i_i_0_a2\ : CFG2
      generic map(INIT => x"1")

      port map(A => \hash_control_st_reg_2\, B => 
        \hash_control_st_reg[4]_net_1\, Y => N_398);
    
    \msg_bit_cnt_reg[49]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_46_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[49]\);
    
    \hash_control_st_reg_i[6]\ : SLE
      port map(D => \hash_control_st_reg_nsss_i_0[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \hash_control_st_reg_i[6]_net_1\);
    
    \st_cnt_reg_cry[5]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[5]\, 
        D => GND_net_1, FCI => \st_cnt_reg_cry[4]_net_1\, S => 
        \st_cnt_reg_s[5]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[5]_net_1\);
    
    \oregs_ce_i_a2_0_a2\ : CFG2
      generic map(INIT => x"2")

      port map(A => \hash_control_st_reg_i[6]_net_1\, B => 
        \hash_control_st_reg[3]_net_1\, Y => 
        oregs_ce_i_a2_0_a2_net_1);
    
    un1_msg_bit_cnt_reg_cry_55 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[58]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_54\, S => 
        un1_msg_bit_cnt_reg_cry_55_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_55\);
    
    \msg_bit_cnt_reg[28]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_25_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[28]\);
    
    un1_msg_bit_cnt_reg_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_6\, S => 
        un1_msg_bit_cnt_reg_cry_7_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_7\);
    
    \state_counter_proc.un15_ce_i_i_0_a2_RNIM61C1\ : CFG4
      generic map(INIT => x"FF15")

      port map(A => ce_i_i_2, B => N_398, C => N_115, D => 
        st_cnt_clr, Y => st_cnt_rege);
    
    un1_msg_bit_cnt_reg_cry_42 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[45]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_41\, S => 
        un1_msg_bit_cnt_reg_cry_42_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_42\);
    
    \msg_bit_cnt_reg[44]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_41_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[44]\);
    
    \hash_control_st_reg_r[5]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => last_block_0, B => N_341, C => N_355, D => 
        \hash_control_st_reg_ns_i_0_1[1]_net_1\, Y => 
        hash_control_st_reg_4);
    
    \hash_control_st_reg_ns_0_0_a2[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \hash_control_st_reg_i[6]_net_1\, B => N_28, 
        Y => N_391);
    
    un1_msg_bit_cnt_reg_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[13]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_9\, S => 
        un1_msg_bit_cnt_reg_cry_10_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_10\);
    
    \hash_control_st_reg_ns_0_0_a4[3]\ : CFG3
      generic map(INIT => x"20")

      port map(A => ce_i_i_2, B => N_28, C => 
        \hash_control_st_reg[3]_net_1\, Y => N_363);
    
    st_cnt_reg_5_rep1 : SLE
      port map(D => \st_cnt_reg_s[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_5_rep1);
    
    un1_msg_bit_cnt_reg_cry_54 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[57]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_53\, S => 
        un1_msg_bit_cnt_reg_cry_54_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_54\);
    
    \msg_bit_cnt_reg[57]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_54_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[57]\);
    
    un1_msg_bit_cnt_reg_cry_58 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[61]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_57\, S => 
        un1_msg_bit_cnt_reg_cry_58_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_58\);
    
    un1_msg_bit_cnt_reg_cry_56 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[59]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_55\, S => 
        un1_msg_bit_cnt_reg_cry_56_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_56\);
    
    un1_msg_bit_cnt_reg_cry_39 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[42]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_38\, S => 
        un1_msg_bit_cnt_reg_cry_39_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_39\);
    
    un1_msg_bit_cnt_reg_cry_51 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[54]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_50\, S => 
        un1_msg_bit_cnt_reg_cry_51_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_51\);
    
    \msg_bit_cnt_reg[60]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_57_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[60]\);
    
    un1_msg_bit_cnt_reg_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_2\, S => 
        un1_msg_bit_cnt_reg_cry_3_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_3\);
    
    \msg_bit_cnt_reg[56]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_53_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[56]\);
    
    \msg_bit_cnt_reg[5]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_2_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[5]\);
    
    \msg_bit_cnt_reg[33]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_30_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[33]\);
    
    \msg_bit_cnt_reg[61]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_58_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[61]\);
    
    un1_msg_bit_cnt_reg_cry_35 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[38]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_34\, S => 
        un1_msg_bit_cnt_reg_cry_35_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_35\);
    
    pad_one_reg_0_0_a4_0 : CFG4
      generic map(INIT => x"0800")

      port map(A => \hash_control_st_reg_i[6]_net_1\, B => N_115, 
        C => \hash_control_st_reg_2\, D => \one_insert\, Y => 
        N_368);
    
    \hash_control_st_reg[5]\ : SLE
      port map(D => hash_control_st_reg_4, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_Module_0_di_req_o\);
    
    \msg_bit_cnt_reg[8]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_5_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[8]\);
    
    \st_cnt_reg[0]\ : SLE
      port map(D => \st_cnt_reg_s[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \Kt_addr[0]\);
    
    un1_msg_bit_cnt_reg_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[16]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_12\, S => 
        un1_msg_bit_cnt_reg_cry_13_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_13\);
    
    un1_msg_bit_cnt_reg_cry_34 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[37]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_33\, S => 
        un1_msg_bit_cnt_reg_cry_34_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_34\);
    
    un1_msg_bit_cnt_reg_cry_38 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[41]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_37\, S => 
        un1_msg_bit_cnt_reg_cry_38_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_38\);
    
    un1_msg_bit_cnt_reg_cry_36 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[39]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_35\, S => 
        un1_msg_bit_cnt_reg_cry_36_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_36\);
    
    un1_msg_bit_cnt_reg_cry_31 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[34]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_30\, S => 
        un1_msg_bit_cnt_reg_cry_31_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_31\);
    
    padding_reg_0_0 : CFG4
      generic map(INIT => x"AEFF")

      port map(A => \padding_reg\, B => \hash_control_st_reg_2\, 
        C => ce_i_i_2, D => \hash_control_st_reg_i[6]_net_1\, Y
         => \padding_reg_0_0\);
    
    \msg_bit_cnt_reg[20]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_17_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[20]\);
    
    \msg_bit_cnt_reg[55]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_52_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[55]\);
    
    un1_msg_bit_cnt_reg_cry_22 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[25]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_21\, S => 
        un1_msg_bit_cnt_reg_cry_22_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_22\);
    
    
        \core_error_combi_proc.core_error_combi_proc.un9_core_error_0_a4\ : 
        CFG3
      generic map(INIT => x"10")

      port map(A => sha256_controller_0_end_o, B => N_115, C => 
        sha256_controller_0_bytes_o(1), Y => N_375);
    
    \msg_bit_cnt_reg[7]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_4_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[7]\);
    
    un1_msg_bit_cnt_reg_cry_40 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[43]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_39\, S => 
        un1_msg_bit_cnt_reg_cry_40_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_40\);
    
    st_cnt_reg_3_rep1 : SLE
      port map(D => \st_cnt_reg_s[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_3_rep1);
    
    \msg_bit_cnt_reg[59]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_56_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[59]\);
    
    \msg_bit_cnt_reg[21]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_18_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[21]\);
    
    \msg_bit_cnt_reg[9]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_6_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[9]\);
    
    \hash_control_st_reg_ns_i_0_o2_2[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \Kt_addr[0]\, B => ce_i_i_2, Y => N_149);
    
    \msg_bit_cnt_reg[37]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_34_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[37]\);
    
    un1_msg_bit_cnt_reg_cry_19 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[22]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_18\, S => 
        un1_msg_bit_cnt_reg_cry_19_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_19\);
    
    \msg_bit_cnt_reg[54]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_51_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[54]\);
    
    \msg_bit_cnt_reg[36]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_33_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[36]\);
    
    un1_msg_bit_cnt_reg_cry_1 : ARI1
      generic map(INIT => x"5BF40")

      port map(A => \msg_bitlen[4]\, B => N_229, C => 
        sha256_controller_0_bytes_o(1), D => 
        sha256_controller_0_end_o, FCI => 
        \un1_msg_bit_cnt_reg_cry_0\, S => 
        un1_msg_bit_cnt_reg_cry_1_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_1\);
    
    pad_one_reg_0_0_a4 : CFG4
      generic map(INIT => x"C800")

      port map(A => \pad_one_reg_0_0_o2_0\, B => \one_insert\, C
         => \N_387\, D => \hash_control_st_reg_i[6]_net_1\, Y => 
        N_367);
    
    \msg_bit_cnt_reg[12]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_9_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[12]\);
    
    \hash_control_st_reg_ns_i_0_a4_0[4]\ : CFG4
      generic map(INIT => x"0023")

      port map(A => N_119, B => N_28, C => \padding_reg\, D => 
        \hash_control_st_reg_2\, Y => N_357);
    
    \st_cnt_reg_fast[5]\ : SLE
      port map(D => \st_cnt_reg_s[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => st_cnt_rege, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => Kt_addr_fast(5));
    
    un1_msg_bit_cnt_reg_cry_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[18]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_14\, S => 
        un1_msg_bit_cnt_reg_cry_15_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_15\);
    
    \hash_control_st_reg_r[4]\ : CFG4
      generic map(INIT => x"4055")

      port map(A => last_block_0, B => N_389, C => N_228, D => 
        \hash_control_st_reg_r_1[4]_net_1\, Y => 
        hash_control_st_reg);
    
    un1_msg_bit_cnt_reg_cry_43 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[46]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_42\, S => 
        un1_msg_bit_cnt_reg_cry_43_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_43\);
    
    \msg_bit_cnt_reg[18]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_15_S, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[18]\);
    
    pad_one_reg_0_0_a2_0_0 : CFG2
      generic map(INIT => x"1")

      port map(A => \Kt_addr_fast[1]\, B => \Kt_addr_fast[2]\, Y
         => pad_one_reg_0_0_a2_0);
    
    
        \core_error_combi_proc.core_error_combi_proc.un9_core_error_0\ : 
        CFG4
      generic map(INIT => x"FCFE")

      port map(A => N_391, B => N_375, C => 
        \hash_control_st_reg[0]_net_1\, D => 
        \SHA256_Module_0_di_req_o\, Y => SHA256_Module_0_error_o);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_hash_core is

    port( R1_data                      : out   std_logic_vector(31 downto 0);
          R2_data                      : out   std_logic_vector(31 downto 0);
          R3_data                      : out   std_logic_vector(31 downto 0);
          R5_data                      : out   std_logic_vector(31 downto 0);
          R6_data                      : out   std_logic_vector(31 downto 0);
          R7_data                      : out   std_logic_vector(31 downto 0);
          R0_data                      : out   std_logic_vector(31 downto 0);
          R4_data                      : out   std_logic_vector(31 downto 0);
          N4_data                      : in    std_logic_vector(31 downto 1);
          N0_data                      : in    std_logic_vector(31 downto 1);
          W_out_i_0                    : in    std_logic_vector(0 to 0);
          Kt_addr                      : in    std_logic_vector(5 to 5);
          N3_data                      : in    std_logic_vector(31 downto 1);
          N2_data                      : in    std_logic_vector(31 downto 1);
          N1_data                      : in    std_logic_vector(31 downto 1);
          N7_data                      : in    std_logic_vector(31 downto 1);
          N6_data                      : in    std_logic_vector(31 downto 1);
          N5_data                      : in    std_logic_vector(31 downto 1);
          Wt_data                      : in    std_logic_vector(31 downto 0);
          Kt_data_15                   : in    std_logic;
          Kt_data_24                   : in    std_logic;
          Kt_data_0                    : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK : in    std_logic;
          core_ce_o_iv_i_0             : in    std_logic;
          oregs_ce_i_a2_0_a2           : in    std_logic;
          next_reg_H4_cry_0_0_Y        : in    std_logic;
          next_reg_H0_cry_0_0_Y        : in    std_logic;
          next_r0_0_cry_0_Y            : in    std_logic;
          ld_i_i_3                     : in    std_logic;
          N_98                         : in    std_logic;
          m10_bm                       : in    std_logic;
          m20_1                        : in    std_logic;
          m10_am                       : in    std_logic;
          m34                          : in    std_logic;
          m49_am                       : in    std_logic;
          m49_bm                       : in    std_logic;
          Kt_addr_5_rep1               : in    std_logic;
          m62_am                       : in    std_logic;
          m62_bm                       : in    std_logic;
          m67_ns                       : in    std_logic;
          m73                          : in    std_logic;
          m78                          : in    std_logic;
          m83_ns                       : in    std_logic;
          m95_1_0                      : in    std_logic;
          m95_1_1                      : in    std_logic;
          m104_am                      : in    std_logic;
          m104_bm                      : in    std_logic;
          m110_ns                      : in    std_logic;
          m114                         : in    std_logic;
          m119_ns                      : in    std_logic;
          m124                         : in    std_logic;
          m137_am                      : in    std_logic;
          m137_bm                      : in    std_logic;
          m141                         : in    std_logic;
          m144_ns                      : in    std_logic;
          m157                         : in    std_logic;
          m168_1_0                     : in    std_logic;
          m168_1_1                     : in    std_logic;
          m172_ns                      : in    std_logic;
          m177                         : in    std_logic;
          m197_1_0                     : in    std_logic;
          m197_1_1                     : in    std_logic;
          m207_1_0                     : in    std_logic;
          m207_1_1                     : in    std_logic;
          m215_am                      : in    std_logic;
          m215_bm                      : in    std_logic;
          m219                         : in    std_logic;
          m222_ns                      : in    std_logic;
          m226_ns                      : in    std_logic;
          m230                         : in    std_logic;
          m235_ns                      : in    std_logic;
          m239                         : in    std_logic;
          m250_am                      : in    std_logic;
          m250_bm                      : in    std_logic;
          m254                         : in    std_logic;
          m258_ns                      : in    std_logic;
          m273                         : in    std_logic;
          m276_ns                      : in    std_logic;
          m281_ns                      : in    std_logic;
          m285                         : in    std_logic;
          m289                         : in    std_logic;
          m292_ns                      : in    std_logic;
          m296                         : in    std_logic;
          m300_ns                      : in    std_logic;
          m304                         : in    std_logic;
          i3_mux_1                     : in    std_logic;
          m325                         : in    std_logic;
          m316                         : in    std_logic;
          next_reg_H3_cry_0_0_Y        : in    std_logic;
          next_reg_H2_cry_0_0_Y        : in    std_logic;
          next_reg_H1_cry_0_0_Y        : in    std_logic;
          next_reg_H7_cry_0_0_Y        : in    std_logic;
          next_reg_H6_cry_0_0_Y        : in    std_logic;
          next_reg_H5_cry_0_0_Y        : in    std_logic
        );

end sha256_hash_core;

architecture DEF_ARCH of sha256_hash_core is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \R1_data[31]\, VCC_net_1, \next_reg_b[31]_net_1\, 
        GND_net_1, \R1_data[16]\, \next_reg_b[16]_net_1\, 
        \R1_data[17]\, \next_reg_b[17]_net_1\, \R1_data[18]\, 
        \next_reg_b[18]_net_1\, \R1_data[19]\, 
        \next_reg_b[19]_net_1\, \R1_data[20]\, 
        \next_reg_b[20]_net_1\, \R1_data[21]\, 
        \next_reg_b[21]_net_1\, \R1_data[22]\, 
        \next_reg_b[22]_net_1\, \R1_data[23]\, 
        \next_reg_b[23]_net_1\, \R1_data[24]\, 
        \next_reg_b[24]_net_1\, \R1_data[25]\, 
        \next_reg_b[25]_net_1\, \R1_data[26]\, 
        \next_reg_b[26]_net_1\, \R1_data[27]\, 
        \next_reg_b[27]_net_1\, \R1_data[28]\, 
        \next_reg_b[28]_net_1\, \R1_data[29]\, 
        \next_reg_b[29]_net_1\, \R1_data[30]\, 
        \next_reg_b[30]_net_1\, \R1_data[1]\, 
        \next_reg_b[1]_net_1\, \R1_data[2]\, 
        \next_reg_b[2]_net_1\, \R1_data[3]\, 
        \next_reg_b[3]_net_1\, \R1_data[4]\, 
        \next_reg_b[4]_net_1\, \R1_data[5]\, 
        \next_reg_b[5]_net_1\, \R1_data[6]\, 
        \next_reg_b[6]_net_1\, \R1_data[7]\, 
        \next_reg_b[7]_net_1\, \R1_data[8]\, 
        \next_reg_b[8]_net_1\, \R1_data[9]\, 
        \next_reg_b[9]_net_1\, \R1_data[10]\, 
        \next_reg_b[10]_net_1\, \R1_data[11]\, 
        \next_reg_b[11]_net_1\, \R1_data[12]\, 
        \next_reg_b[12]_net_1\, \R1_data[13]\, 
        \next_reg_b[13]_net_1\, \R1_data[14]\, 
        \next_reg_b[14]_net_1\, \R1_data[15]\, 
        \next_reg_b[15]_net_1\, \R2_data[18]\, 
        \next_reg_c[18]_net_1\, \R2_data[19]\, 
        \next_reg_c[19]_net_1\, \R2_data[20]\, 
        \next_reg_c[20]_net_1\, \R2_data[21]\, 
        \next_reg_c[21]_net_1\, \R2_data[22]\, 
        \next_reg_c[22]_net_1\, \R2_data[23]\, 
        \next_reg_c[23]_net_1\, \R2_data[24]\, 
        \next_reg_c[24]_net_1\, \R2_data[25]\, 
        \next_reg_c[25]_net_1\, \R2_data[26]\, 
        \next_reg_c[26]_net_1\, \R2_data[27]\, 
        \next_reg_c[27]_net_1\, \R2_data[28]\, 
        \next_reg_c[28]_net_1\, \R2_data[29]\, 
        \next_reg_c[29]_net_1\, \R2_data[30]\, 
        \next_reg_c[30]_net_1\, \R2_data[31]\, 
        \next_reg_c[31]_net_1\, \R1_data[0]\, 
        \next_reg_b[0]_net_1\, \R2_data[3]\, 
        \next_reg_c[3]_net_1\, \R2_data[4]\, 
        \next_reg_c[4]_net_1\, \R2_data[5]\, 
        \next_reg_c[5]_net_1\, \R2_data[6]\, 
        \next_reg_c[6]_net_1\, \R2_data[7]\, 
        \next_reg_c[7]_net_1\, \R2_data[8]\, 
        \next_reg_c[8]_net_1\, \R2_data[9]\, 
        \next_reg_c[9]_net_1\, \R2_data[10]\, 
        \next_reg_c[10]_net_1\, \R2_data[11]\, 
        \next_reg_c[11]_net_1\, \R2_data[12]\, 
        \next_reg_c[12]_net_1\, \R2_data[13]\, 
        \next_reg_c[13]_net_1\, \R2_data[14]\, 
        \next_reg_c[14]_net_1\, \R2_data[15]\, 
        \next_reg_c[15]_net_1\, \R2_data[16]\, 
        \next_reg_c[16]_net_1\, \R2_data[17]\, 
        \next_reg_c[17]_net_1\, \R3_data[20]\, 
        \next_reg_d[20]_net_1\, \R3_data[21]\, 
        \next_reg_d[21]_net_1\, \R3_data[22]\, 
        \next_reg_d[22]_net_1\, \R3_data[23]\, 
        \next_reg_d[23]_net_1\, \R3_data[24]\, 
        \next_reg_d[24]_net_1\, \R3_data[25]\, 
        \next_reg_d[25]_net_1\, \R3_data[26]\, 
        \next_reg_d[26]_net_1\, \R3_data[27]\, 
        \next_reg_d[27]_net_1\, \R3_data[28]\, 
        \next_reg_d[28]_net_1\, \R3_data[29]\, 
        \next_reg_d[29]_net_1\, \R3_data[30]\, 
        \next_reg_d[30]_net_1\, \R3_data[31]\, 
        \next_reg_d[31]_net_1\, \R2_data[0]\, 
        \next_reg_c[0]_net_1\, \R2_data[1]\, 
        \next_reg_c[1]_net_1\, \R2_data[2]\, 
        \next_reg_c[2]_net_1\, \R3_data[5]\, 
        \next_reg_d[5]_net_1\, \R3_data[6]\, 
        \next_reg_d[6]_net_1\, \R3_data[7]\, 
        \next_reg_d[7]_net_1\, \R3_data[8]\, 
        \next_reg_d[8]_net_1\, \R3_data[9]\, 
        \next_reg_d[9]_net_1\, \R3_data[10]\, 
        \next_reg_d[10]_net_1\, \R3_data[11]\, 
        \next_reg_d[11]_net_1\, \R3_data[12]\, 
        \next_reg_d[12]_net_1\, \R3_data[13]\, 
        \next_reg_d[13]_net_1\, \R3_data[14]\, 
        \next_reg_d[14]_net_1\, \R3_data[15]\, 
        \next_reg_d[15]_net_1\, \R3_data[16]\, 
        \next_reg_d[16]_net_1\, \R3_data[17]\, 
        \next_reg_d[17]_net_1\, \R3_data[18]\, 
        \next_reg_d[18]_net_1\, \R3_data[19]\, 
        \next_reg_d[19]_net_1\, \R5_data[22]\, 
        \next_reg_f[22]_net_1\, \R5_data[23]\, 
        \next_reg_f[23]_net_1\, \R5_data[24]\, 
        \next_reg_f[24]_net_1\, \R5_data[25]\, 
        \next_reg_f[25]_net_1\, \R5_data[26]\, 
        \next_reg_f[26]_net_1\, \R5_data[27]\, 
        \next_reg_f[27]_net_1\, \R5_data[28]\, 
        \next_reg_f[28]_net_1\, \R5_data[29]\, 
        \next_reg_f[29]_net_1\, \R5_data[30]\, 
        \next_reg_f[30]_net_1\, \R5_data[31]\, 
        \next_reg_f[31]_net_1\, \R3_data[0]\, 
        \next_reg_d[0]_net_1\, \R3_data[1]\, 
        \next_reg_d[1]_net_1\, \R3_data[2]\, 
        \next_reg_d[2]_net_1\, \R3_data[3]\, 
        \next_reg_d[3]_net_1\, \R3_data[4]\, 
        \next_reg_d[4]_net_1\, \R5_data[7]\, 
        \next_reg_f[7]_net_1\, \R5_data[8]\, 
        \next_reg_f[8]_net_1\, \R5_data[9]\, 
        \next_reg_f[9]_net_1\, \R5_data[10]\, 
        \next_reg_f[10]_net_1\, \R5_data[11]\, 
        \next_reg_f[11]_net_1\, \R5_data[12]\, 
        \next_reg_f[12]_net_1\, \R5_data[13]\, 
        \next_reg_f[13]_net_1\, \R5_data[14]\, 
        \next_reg_f[14]_net_1\, \R5_data[15]\, 
        \next_reg_f[15]_net_1\, \R5_data[16]\, 
        \next_reg_f[16]_net_1\, \R5_data[17]\, 
        \next_reg_f[17]_net_1\, \R5_data[18]\, 
        \next_reg_f[18]_net_1\, \R5_data[19]\, 
        \next_reg_f[19]_net_1\, \R5_data[20]\, 
        \next_reg_f[20]_net_1\, \R5_data[21]\, 
        \next_reg_f[21]_net_1\, \R6_data[24]\, 
        \next_reg_g[24]_net_1\, \R6_data[25]\, 
        \next_reg_g[25]_net_1\, \R6_data[26]\, 
        \next_reg_g[26]_net_1\, \R6_data[27]\, 
        \next_reg_g[27]_net_1\, \R6_data[28]\, 
        \next_reg_g[28]_net_1\, \R6_data[29]\, 
        \next_reg_g[29]_net_1\, \R6_data[30]\, 
        \next_reg_g[30]_net_1\, \R6_data[31]\, 
        \next_reg_g[31]_net_1\, \R5_data[0]\, 
        \next_reg_f[0]_net_1\, \R5_data[1]\, 
        \next_reg_f[1]_net_1\, \R5_data[2]\, 
        \next_reg_f[2]_net_1\, \R5_data[3]\, 
        \next_reg_f[3]_net_1\, \R5_data[4]\, 
        \next_reg_f[4]_net_1\, \R5_data[5]\, 
        \next_reg_f[5]_net_1\, \R5_data[6]\, 
        \next_reg_f[6]_net_1\, \R6_data[9]\, 
        \next_reg_g[9]_net_1\, \R6_data[10]\, 
        \next_reg_g[10]_net_1\, \R6_data[11]\, 
        \next_reg_g[11]_net_1\, \R6_data[12]\, 
        \next_reg_g[12]_net_1\, \R6_data[13]\, 
        \next_reg_g[13]_net_1\, \R6_data[14]\, 
        \next_reg_g[14]_net_1\, \R6_data[15]\, 
        \next_reg_g[15]_net_1\, \R6_data[16]\, 
        \next_reg_g[16]_net_1\, \R6_data[17]\, 
        \next_reg_g[17]_net_1\, \R6_data[18]\, 
        \next_reg_g[18]_net_1\, \R6_data[19]\, 
        \next_reg_g[19]_net_1\, \R6_data[20]\, 
        \next_reg_g[20]_net_1\, \R6_data[21]\, 
        \next_reg_g[21]_net_1\, \R6_data[22]\, 
        \next_reg_g[22]_net_1\, \R6_data[23]\, 
        \next_reg_g[23]_net_1\, \R7_data[26]\, 
        \next_reg_h[26]_net_1\, \R7_data[27]\, 
        \next_reg_h[27]_net_1\, \R7_data[28]\, 
        \next_reg_h[28]_net_1\, \R7_data[29]\, 
        \next_reg_h[29]_net_1\, \R7_data[30]\, 
        \next_reg_h[30]_net_1\, \R7_data[31]\, 
        \next_reg_h[31]_net_1\, \R6_data[0]\, 
        \next_reg_g[0]_net_1\, \R6_data[1]\, 
        \next_reg_g[1]_net_1\, \R6_data[2]\, 
        \next_reg_g[2]_net_1\, \R6_data[3]\, 
        \next_reg_g[3]_net_1\, \R6_data[4]\, 
        \next_reg_g[4]_net_1\, \R6_data[5]\, 
        \next_reg_g[5]_net_1\, \R6_data[6]\, 
        \next_reg_g[6]_net_1\, \R6_data[7]\, 
        \next_reg_g[7]_net_1\, \R6_data[8]\, 
        \next_reg_g[8]_net_1\, \R7_data[11]\, 
        \next_reg_h[11]_net_1\, \R7_data[12]\, 
        \next_reg_h[12]_net_1\, \R7_data[13]\, 
        \next_reg_h[13]_net_1\, \R7_data[14]\, 
        \next_reg_h[14]_net_1\, \R7_data[15]\, 
        \next_reg_h[15]_net_1\, \R7_data[16]\, 
        \next_reg_h[16]_net_1\, \R7_data[17]\, 
        \next_reg_h[17]_net_1\, \R7_data[18]\, 
        \next_reg_h[18]_net_1\, \R7_data[19]\, 
        \next_reg_h[19]_net_1\, \R7_data[20]\, 
        \next_reg_h[20]_net_1\, \R7_data[21]\, 
        \next_reg_h[21]_net_1\, \R7_data[22]\, 
        \next_reg_h[22]_net_1\, \R7_data[23]\, 
        \next_reg_h[23]_net_1\, \R7_data[24]\, 
        \next_reg_h[24]_net_1\, \R7_data[25]\, 
        \next_reg_h[25]_net_1\, \R0_data[28]\, \next_reg_a[28]\, 
        \R0_data[29]\, \next_reg_a[29]\, \R0_data[30]\, 
        \next_reg_a[30]\, \R0_data[31]\, \next_reg_a[31]\, 
        \R7_data[0]\, \next_reg_h[0]_net_1\, \R7_data[1]\, 
        \next_reg_h[1]_net_1\, \R7_data[2]\, 
        \next_reg_h[2]_net_1\, \R7_data[3]\, 
        \next_reg_h[3]_net_1\, \R7_data[4]\, 
        \next_reg_h[4]_net_1\, \R7_data[5]\, 
        \next_reg_h[5]_net_1\, \R7_data[6]\, 
        \next_reg_h[6]_net_1\, \R7_data[7]\, 
        \next_reg_h[7]_net_1\, \R7_data[8]\, 
        \next_reg_h[8]_net_1\, \R7_data[9]\, 
        \next_reg_h[9]_net_1\, \R7_data[10]\, 
        \next_reg_h[10]_net_1\, \R0_data[13]\, \next_reg_a[13]\, 
        \R0_data[14]\, \next_reg_a[14]\, \R0_data[15]\, 
        \next_reg_a[15]\, \R0_data[16]\, \next_reg_a[16]\, 
        \R0_data[17]\, \next_reg_a[17]\, \R0_data[18]\, 
        \next_reg_a[18]\, \R0_data[19]\, \next_reg_a[19]\, 
        \R0_data[20]\, \next_reg_a[20]\, \R0_data[21]\, 
        \next_reg_a[21]\, \R0_data[22]\, \next_reg_a[22]\, 
        \R0_data[23]\, \next_reg_a[23]\, \R0_data[24]\, 
        \next_reg_a[24]\, \R0_data[25]\, \next_reg_a[25]\, 
        \R0_data[26]\, \next_reg_a[26]\, \R0_data[27]\, 
        \next_reg_a[27]\, \R4_data[30]\, \next_reg_e[30]\, 
        \R4_data[31]\, \next_reg_e[31]\, \R0_data[0]\, 
        next_reg_a_cry_0_0_Y, \R0_data[1]\, \next_reg_a[1]\, 
        \R0_data[2]\, \next_reg_a[2]\, \R0_data[3]\, 
        \next_reg_a[3]\, \R0_data[4]\, \next_reg_a[4]\, 
        \R0_data[5]\, \next_reg_a[5]\, \R0_data[6]\, 
        \next_reg_a[6]\, \R0_data[7]\, \next_reg_a[7]\, 
        \R0_data[8]\, \next_reg_a[8]\, \R0_data[9]\, 
        \next_reg_a[9]\, \R0_data[10]\, \next_reg_a[10]\, 
        \R0_data[11]\, \next_reg_a[11]\, \R0_data[12]\, 
        \next_reg_a[12]\, \R4_data[15]\, \next_reg_e[15]\, 
        \R4_data[16]\, \next_reg_e[16]\, \R4_data[17]\, 
        \next_reg_e[17]\, \R4_data[18]\, \next_reg_e[18]\, 
        \R4_data[19]\, \next_reg_e[19]\, \R4_data[20]\, 
        \next_reg_e[20]\, \R4_data[21]\, \next_reg_e[21]\, 
        \R4_data[22]\, \next_reg_e[22]\, \R4_data[23]\, 
        \next_reg_e[23]\, \R4_data[24]\, \next_reg_e[24]\, 
        \R4_data[25]\, \next_reg_e[25]\, \R4_data[26]\, 
        \next_reg_e[26]\, \R4_data[27]\, \next_reg_e[27]\, 
        \R4_data[28]\, \next_reg_e[28]\, \R4_data[29]\, 
        \next_reg_e[29]\, \R4_data[0]\, next_reg_e_cry_0_0_Y, 
        \R4_data[1]\, \next_reg_e[1]\, \R4_data[2]\, 
        \next_reg_e[2]\, \R4_data[3]\, \next_reg_e[3]\, 
        \R4_data[4]\, \next_reg_e[4]\, \R4_data[5]\, 
        \next_reg_e[5]\, \R4_data[6]\, \next_reg_e[6]\, 
        \R4_data[7]\, \next_reg_e[7]\, \R4_data[8]\, 
        \next_reg_e[8]\, \R4_data[9]\, \next_reg_e[9]\, 
        \R4_data[10]\, \next_reg_e[10]\, \R4_data[11]\, 
        \next_reg_e[11]\, \R4_data[12]\, \next_reg_e[12]\, 
        \R4_data[13]\, \next_reg_e[13]\, \R4_data[14]\, 
        \next_reg_e[14]\, next_reg_e_cry_0, sum3_cry_0_Y, 
        next_reg_e_cry_1, \sum3[1]\, next_reg_e_cry_2, \sum3[2]\, 
        next_reg_e_cry_3, \sum3[3]\, next_reg_e_cry_4, \sum3[4]\, 
        next_reg_e_cry_5, \sum3[5]\, next_reg_e_cry_6, \sum3[6]\, 
        next_reg_e_cry_7, \sum3[7]\, next_reg_e_cry_8, \sum3[8]\, 
        next_reg_e_cry_9, \sum3[9]\, next_reg_e_cry_10, 
        \sum3[10]\, next_reg_e_cry_11, \sum3[11]\, 
        next_reg_e_cry_12, \sum3[12]\, next_reg_e_cry_13, 
        \sum3[13]\, next_reg_e_cry_14, \sum3[14]\, 
        next_reg_e_cry_15, \sum3[15]\, next_reg_e_cry_16, 
        \sum3[16]\, next_reg_e_cry_17, \sum3[17]\, 
        next_reg_e_cry_18, \sum3[18]\, next_reg_e_cry_19, 
        \sum3[19]\, next_reg_e_cry_20, \sum3[20]\, 
        next_reg_e_cry_21, \sum3[21]\, next_reg_e_cry_22, 
        \sum3[22]\, next_reg_e_cry_23, \sum3[23]\, 
        next_reg_e_cry_24, \sum3[24]\, next_reg_e_cry_25, 
        \sum3[25]\, next_reg_e_cry_26, \sum3[26]\, 
        next_reg_e_cry_27, \sum3[27]\, next_reg_e_cry_28, 
        \sum3[28]\, next_reg_e_cry_29, \sum3[29]\, \sum3[31]\, 
        next_reg_e_cry_30, \sum3[30]\, next_reg_a_cry_0, 
        sum0_4_cry_0_Y_0, next_reg_a_cry_1, \sum0_4[1]\, 
        next_reg_a_cry_2, \sum0_4[2]\, next_reg_a_cry_3, 
        \sum0_4[3]\, next_reg_a_cry_4, \sum0_4[4]\, 
        next_reg_a_cry_5, \sum0_4[5]\, next_reg_a_cry_6, 
        \sum0_4[6]\, next_reg_a_cry_7, \sum0_4[7]\, 
        next_reg_a_cry_8, \sum0_4[8]\, next_reg_a_cry_9, 
        \sum0_4[9]\, next_reg_a_cry_10, \sum0_4[10]\, 
        next_reg_a_cry_11, \sum0_4[11]\, next_reg_a_cry_12, 
        \sum0_4[12]\, next_reg_a_cry_13, \sum0_4[13]\, 
        next_reg_a_cry_14, \sum0_4[14]\, next_reg_a_cry_15, 
        \sum0_4[15]\, next_reg_a_cry_16, \sum0_4[16]\, 
        next_reg_a_cry_17, \sum0_4[17]\, next_reg_a_cry_18, 
        \sum0_4[18]\, next_reg_a_cry_19, \sum0_4[19]\, 
        next_reg_a_cry_20, \sum0_4[20]\, next_reg_a_cry_21, 
        \sum0_4[21]\, next_reg_a_cry_22, \sum0_4[22]\, 
        next_reg_a_cry_23, \sum0_4[23]\, next_reg_a_cry_24, 
        \sum0_4[24]\, next_reg_a_cry_25, \sum0_4[25]\, 
        next_reg_a_cry_26, \sum0_4[26]\, next_reg_a_cry_27, 
        \sum0_4[27]\, next_reg_a_cry_28, \sum0_4[28]\, 
        next_reg_a_cry_29, \sum0_4[29]\, \sum0_4[31]\, 
        next_reg_a_cry_30, \sum0_4[30]\, \sum0_4_cry_0\, sum0_4_0, 
        \sum0_4[0]\, \sum0_4_cry_1\, \SIG0_0[1]\, \sum0_4_axb_1\, 
        \sum0_4_cry_2\, \SIG0_0[2]\, \sum0_4_axb_2\, 
        \sum0_4_cry_3\, \SIG0_0[3]\, \sum0_4_axb_3\, 
        \sum0_4_cry_4\, \SIG0_0[4]\, \sum0_4_axb_4\, 
        \sum0_4_cry_5\, \SIG0_0[5]\, \sum0_4_axb_5\, 
        \sum0_4_cry_6\, \SIG0_0[6]\, \sum0_4_axb_6\, 
        \sum0_4_cry_7\, \SIG0_0[7]\, \sum0_4_axb_7\, 
        \sum0_4_cry_8\, \SIG0_0[8]\, \sum0_4_axb_8\, 
        \sum0_4_cry_9\, \SIG0_0[9]\, \sum0_4_axb_9\, 
        \sum0_4_cry_10\, \SIG0_0[10]\, \sum0_4_axb_10\, 
        \sum0_4_cry_11\, \SIG0_0[11]\, \sum0_4_axb_11\, 
        \sum0_4_cry_12\, \SIG0_0[12]\, \sum0_4_axb_12\, 
        \sum0_4_cry_13\, \SIG0_0[13]\, \sum0_4_axb_13\, 
        \sum0_4_cry_14\, \SIG0_0[14]\, \sum0_4_axb_14\, 
        \sum0_4_cry_15\, \SIG0_0[15]\, \sum0_4_axb_15\, 
        \sum0_4_cry_16\, \SIG0_0[16]\, \sum0_4_axb_16\, 
        \sum0_4_cry_17\, \SIG0_0[17]\, \sum0_4_axb_17\, 
        \sum0_4_cry_18\, \SIG0_0[18]\, \sum0_4_axb_18\, 
        \sum0_4_cry_19\, \SIG0_0[19]\, \sum0_4_axb_19\, 
        \sum0_4_cry_20\, \SIG0_0[20]\, \sum0_4_axb_20\, 
        \sum0_4_cry_21\, \SIG0_0[21]\, \sum0_4_axb_21\, 
        \sum0_4_cry_22\, \SIG0_0[22]\, \sum0_4_axb_22\, 
        \sum0_4_cry_23\, \SIG0_0[23]\, \sum0_4_axb_23\, 
        \sum0_4_cry_24\, \SIG0_0[24]\, \sum0_4_axb_24\, 
        \sum0_4_cry_25\, \SIG0_0[25]\, \sum0_4_axb_25\, 
        \sum0_4_cry_26\, \SIG0_0[26]\, \sum0_4_axb_26\, 
        \sum0_4_cry_27\, \SIG0_0[27]\, \sum0_4_axb_27\, 
        \sum0_4_cry_28\, \SIG0_0[28]\, \sum0_4_axb_28\, 
        \sum0_4_cry_29\, \SIG0_0[29]\, \sum0_4_axb_29\, 
        \Maj[31]_net_1\, \sum0_4_cry_30\, \SIG0_0[30]\, 
        \sum0_4_axb_30\, \sum3_6_0_cry_0\, sum3_6_0_cry_0_Y, 
        \sum3_6_0_cry_1\, \sum3_6_0[1]\, \sum3_6_0_cry_2\, 
        \sum3_6_0[2]\, \sum3_6_0_cry_3\, \sum3_6_0[3]\, 
        \sum3_6_0_cry_4\, \sum3_6_0[4]\, \sum3_6_0_cry_5\, 
        \sum3_6_0[5]\, \sum3_6_0_cry_6\, \sum3_6_0[6]\, 
        \sum3_6_0_cry_7\, \sum3_6_0[7]\, \sum3_6_0_cry_8\, 
        \sum3_6_0[8]\, \sum3_6_0_cry_9\, \sum3_6_0[9]\, 
        \sum3_6_0_cry_10\, \sum3_6_0[10]\, \sum3_6_0_cry_11\, 
        \sum3_6_0[11]\, \sum3_6_0_cry_12\, \sum3_6_0[12]\, 
        \sum3_6_0_cry_13\, \sum3_6_0[13]\, \sum3_6_0_cry_14\, 
        \sum3_6_0[14]\, \sum3_6_0_cry_15\, \sum3_6_0[15]\, 
        \sum3_6_0_cry_16\, \sum3_6_0[16]\, \sum3_6_0_cry_17\, 
        \sum3_6_0[17]\, \sum3_6_0_cry_18\, \sum3_6_0[18]\, 
        \sum3_6_0_cry_19\, \sum3_6_0[19]\, \sum3_6_0_cry_20\, 
        \sum3_6_0[20]\, \sum3_6_0_cry_21\, \sum3_6_0[21]\, 
        \sum3_6_0_cry_22\, \sum3_6_0[22]\, \sum3_6_0_cry_23\, 
        \sum3_6_0[23]\, \sum3_6_0_cry_24\, \sum3_6_0[24]\, 
        \sum3_6_0_cry_25\, \sum3_6_0[25]\, \sum3_6_0_cry_26\, 
        \sum3_6_0[26]\, \sum3_6_0_cry_27\, \sum3_6_0[27]\, 
        \sum3_6_0_cry_28\, \sum3_6_0[28]\, \sum3_6_0_cry_29\, 
        \sum3_6_0[29]\, \sum3_6_0[31]\, \sum3_6_0_cry_30\, 
        \sum3_6_0[30]\, \sum3_cry_0\, \Wt_data_0[0]\, \sum3[0]\, 
        \sum3_cry_1\, \sum3_4[1]\, \sum3_cry_2\, \sum3_4[2]\, 
        \sum3_cry_3\, \sum3_4[3]\, \sum3_cry_4\, \sum3_4[4]\, 
        \sum3_cry_5\, \sum3_4[5]\, \sum3_cry_6\, \sum3_4[6]\, 
        \sum3_cry_7\, \sum3_4[7]\, \sum3_cry_8\, \sum3_4[8]\, 
        \sum3_cry_9\, \sum3_4[9]\, \sum3_cry_10\, \sum3_4[10]\, 
        \sum3_cry_11\, \sum3_4[11]\, \sum3_cry_12\, \sum3_4[12]\, 
        \sum3_cry_13\, \sum3_4[13]\, \sum3_cry_14\, \sum3_4[14]\, 
        \sum3_cry_15\, \sum3_4[15]\, \sum3_cry_16\, \sum3_4[16]\, 
        \sum3_cry_17\, \sum3_4[17]\, \sum3_cry_18\, \sum3_4[18]\, 
        \sum3_cry_19\, \sum3_4[19]\, \sum3_cry_20\, \sum3_4[20]\, 
        \sum3_cry_21\, \sum3_4[21]\, \sum3_cry_22\, \sum3_4[22]\, 
        \sum3_cry_23\, \sum3_4[23]\, \sum3_cry_24\, \sum3_4[24]\, 
        \sum3_cry_25\, \sum3_4[25]\, \sum3_cry_26\, \sum3_4[26]\, 
        \sum3_cry_27\, \sum3_4[27]\, \sum3_cry_28\, \sum3_4[28]\, 
        \sum3_cry_29\, \sum3_4[29]\, \sum3_4[31]\, \sum3_cry_30\, 
        \sum3_4[30]\, \sum3_4_cry_0\, sum3_4_cry_0_Y, 
        \Kt_data_0[0]\, \sum3_4[0]\, \sum3_4_cry_1\, \sum3_6[1]\, 
        \sum3_4_cry_2\, \sum3_6[2]\, \sum3_4_cry_3\, \sum3_6[3]\, 
        \sum3_4_cry_4\, \sum3_6[4]\, \sum3_4_cry_5\, \sum3_6[5]\, 
        \sum3_4_cry_6\, \sum3_6[6]\, \sum3_4_cry_7\, \sum3_6[7]\, 
        \sum3_4_cry_8\, \sum3_6[8]\, \sum3_4_cry_9\, \sum3_6[9]\, 
        \sum3_4_cry_10\, \sum3_6[10]\, \sum3_4_cry_11\, 
        \sum3_6[11]\, \sum3_4_cry_12\, \sum3_6[12]\, 
        \sum3_4_cry_13\, \sum3_6[13]\, \sum3_4_cry_14\, 
        \sum3_6[14]\, \sum3_4_cry_15\, \sum3_6[15]\, 
        \sum3_4_cry_16\, \sum3_6[16]\, \sum3_4_cry_17\, 
        \sum3_6[17]\, \sum3_4_cry_18\, \sum3_6[18]\, 
        \sum3_4_cry_19\, \sum3_6[19]\, \sum3_4_cry_20\, 
        \sum3_6[20]\, \sum3_4_cry_21\, \sum3_6[21]\, 
        \sum3_4_cry_22\, \sum3_6[22]\, \sum3_4_cry_23\, 
        \sum3_6[23]\, \sum3_4_cry_24\, \sum3_6[24]\, 
        \sum3_4_cry_25\, \sum3_6[25]\, \sum3_4_cry_26\, 
        \sum3_6[26]\, \sum3_4_cry_27\, \sum3_6[27]\, 
        \sum3_4_cry_28\, \sum3_6[28]\, \sum3_4_cry_29\, 
        \sum3_6[29]\, \sum3_6[31]\, \sum3_4_cry_30\, \sum3_6[30]\, 
        \sum3_6_cry_0\, sum3_6_cry_0_Y, sum3_6_0, \sum3_6[0]\, 
        \sum3_6_cry_1\, \sum3_6_cry_2\, \sum3_6_cry_3\, 
        \sum3_6_cry_4\, \sum3_6_cry_5\, \sum3_6_cry_6\, 
        \sum3_6_cry_7\, \sum3_6_cry_8\, \sum3_6_cry_9\, 
        \sum3_6_cry_10\, \sum3_6_cry_11\, \sum3_6_cry_12\, 
        \sum3_6_cry_13\, \sum3_6_cry_14\, \sum3_6_cry_15\, 
        \sum3_6_cry_16\, \sum3_6_cry_17\, \sum3_6_cry_18\, 
        \sum3_6_cry_19\, \sum3_6_cry_20\, \sum3_6_cry_21\, 
        \sum3_6_cry_22\, \sum3_6_cry_23\, \sum3_6_cry_24\, 
        \sum3_6_cry_25\, \sum3_6_cry_26\, \sum3_6_cry_27\, 
        \sum3_6_cry_28\, \sum3_6_cry_29\, \sum3_6_cry_30\, 
        \SIG0[15]_net_1\, \SIG0[14]_net_1\, \SIG0[12]_net_1\, 
        \SIG0[2]_net_1\, \SIG0[30]_net_1\, \SIG0[25]_net_1\, 
        \SIG0[23]_net_1\, \SIG0[19]_net_1\, \SIG0[16]_net_1\, 
        \SIG0[18]_net_1\, \SIG0[27]_net_1\, \SIG0[28]_net_1\, 
        \SIG0[29]_net_1\, \SIG0[4]_net_1\, \SIG0[6]_net_1\, 
        \SIG0[7]_net_1\, \SIG0[17]_net_1\, \SIG0[20]_net_1\, 
        \SIG0[26]_net_1\, \SIG0[5]_net_1\, \SIG0[8]_net_1\, 
        \SIG0[21]_net_1\, \SIG0[9]_net_1\, \SIG0[10]_net_1\, 
        \SIG0[11]_net_1\, sum0_4, \SIG0[22]_net_1\, 
        \SIG0[24]_net_1\, \SIG0[1]_net_1\, \SIG0[3]_net_1\, 
        \SIG0[13]_net_1\ : std_logic;

begin 

    R1_data(31) <= \R1_data[31]\;
    R1_data(30) <= \R1_data[30]\;
    R1_data(29) <= \R1_data[29]\;
    R1_data(28) <= \R1_data[28]\;
    R1_data(27) <= \R1_data[27]\;
    R1_data(26) <= \R1_data[26]\;
    R1_data(25) <= \R1_data[25]\;
    R1_data(24) <= \R1_data[24]\;
    R1_data(23) <= \R1_data[23]\;
    R1_data(22) <= \R1_data[22]\;
    R1_data(21) <= \R1_data[21]\;
    R1_data(20) <= \R1_data[20]\;
    R1_data(19) <= \R1_data[19]\;
    R1_data(18) <= \R1_data[18]\;
    R1_data(17) <= \R1_data[17]\;
    R1_data(16) <= \R1_data[16]\;
    R1_data(15) <= \R1_data[15]\;
    R1_data(14) <= \R1_data[14]\;
    R1_data(13) <= \R1_data[13]\;
    R1_data(12) <= \R1_data[12]\;
    R1_data(11) <= \R1_data[11]\;
    R1_data(10) <= \R1_data[10]\;
    R1_data(9) <= \R1_data[9]\;
    R1_data(8) <= \R1_data[8]\;
    R1_data(7) <= \R1_data[7]\;
    R1_data(6) <= \R1_data[6]\;
    R1_data(5) <= \R1_data[5]\;
    R1_data(4) <= \R1_data[4]\;
    R1_data(3) <= \R1_data[3]\;
    R1_data(2) <= \R1_data[2]\;
    R1_data(1) <= \R1_data[1]\;
    R1_data(0) <= \R1_data[0]\;
    R2_data(31) <= \R2_data[31]\;
    R2_data(30) <= \R2_data[30]\;
    R2_data(29) <= \R2_data[29]\;
    R2_data(28) <= \R2_data[28]\;
    R2_data(27) <= \R2_data[27]\;
    R2_data(26) <= \R2_data[26]\;
    R2_data(25) <= \R2_data[25]\;
    R2_data(24) <= \R2_data[24]\;
    R2_data(23) <= \R2_data[23]\;
    R2_data(22) <= \R2_data[22]\;
    R2_data(21) <= \R2_data[21]\;
    R2_data(20) <= \R2_data[20]\;
    R2_data(19) <= \R2_data[19]\;
    R2_data(18) <= \R2_data[18]\;
    R2_data(17) <= \R2_data[17]\;
    R2_data(16) <= \R2_data[16]\;
    R2_data(15) <= \R2_data[15]\;
    R2_data(14) <= \R2_data[14]\;
    R2_data(13) <= \R2_data[13]\;
    R2_data(12) <= \R2_data[12]\;
    R2_data(11) <= \R2_data[11]\;
    R2_data(10) <= \R2_data[10]\;
    R2_data(9) <= \R2_data[9]\;
    R2_data(8) <= \R2_data[8]\;
    R2_data(7) <= \R2_data[7]\;
    R2_data(6) <= \R2_data[6]\;
    R2_data(5) <= \R2_data[5]\;
    R2_data(4) <= \R2_data[4]\;
    R2_data(3) <= \R2_data[3]\;
    R2_data(2) <= \R2_data[2]\;
    R2_data(1) <= \R2_data[1]\;
    R2_data(0) <= \R2_data[0]\;
    R3_data(31) <= \R3_data[31]\;
    R3_data(30) <= \R3_data[30]\;
    R3_data(29) <= \R3_data[29]\;
    R3_data(28) <= \R3_data[28]\;
    R3_data(27) <= \R3_data[27]\;
    R3_data(26) <= \R3_data[26]\;
    R3_data(25) <= \R3_data[25]\;
    R3_data(24) <= \R3_data[24]\;
    R3_data(23) <= \R3_data[23]\;
    R3_data(22) <= \R3_data[22]\;
    R3_data(21) <= \R3_data[21]\;
    R3_data(20) <= \R3_data[20]\;
    R3_data(19) <= \R3_data[19]\;
    R3_data(18) <= \R3_data[18]\;
    R3_data(17) <= \R3_data[17]\;
    R3_data(16) <= \R3_data[16]\;
    R3_data(15) <= \R3_data[15]\;
    R3_data(14) <= \R3_data[14]\;
    R3_data(13) <= \R3_data[13]\;
    R3_data(12) <= \R3_data[12]\;
    R3_data(11) <= \R3_data[11]\;
    R3_data(10) <= \R3_data[10]\;
    R3_data(9) <= \R3_data[9]\;
    R3_data(8) <= \R3_data[8]\;
    R3_data(7) <= \R3_data[7]\;
    R3_data(6) <= \R3_data[6]\;
    R3_data(5) <= \R3_data[5]\;
    R3_data(4) <= \R3_data[4]\;
    R3_data(3) <= \R3_data[3]\;
    R3_data(2) <= \R3_data[2]\;
    R3_data(1) <= \R3_data[1]\;
    R3_data(0) <= \R3_data[0]\;
    R5_data(31) <= \R5_data[31]\;
    R5_data(30) <= \R5_data[30]\;
    R5_data(29) <= \R5_data[29]\;
    R5_data(28) <= \R5_data[28]\;
    R5_data(27) <= \R5_data[27]\;
    R5_data(26) <= \R5_data[26]\;
    R5_data(25) <= \R5_data[25]\;
    R5_data(24) <= \R5_data[24]\;
    R5_data(23) <= \R5_data[23]\;
    R5_data(22) <= \R5_data[22]\;
    R5_data(21) <= \R5_data[21]\;
    R5_data(20) <= \R5_data[20]\;
    R5_data(19) <= \R5_data[19]\;
    R5_data(18) <= \R5_data[18]\;
    R5_data(17) <= \R5_data[17]\;
    R5_data(16) <= \R5_data[16]\;
    R5_data(15) <= \R5_data[15]\;
    R5_data(14) <= \R5_data[14]\;
    R5_data(13) <= \R5_data[13]\;
    R5_data(12) <= \R5_data[12]\;
    R5_data(11) <= \R5_data[11]\;
    R5_data(10) <= \R5_data[10]\;
    R5_data(9) <= \R5_data[9]\;
    R5_data(8) <= \R5_data[8]\;
    R5_data(7) <= \R5_data[7]\;
    R5_data(6) <= \R5_data[6]\;
    R5_data(5) <= \R5_data[5]\;
    R5_data(4) <= \R5_data[4]\;
    R5_data(3) <= \R5_data[3]\;
    R5_data(2) <= \R5_data[2]\;
    R5_data(1) <= \R5_data[1]\;
    R5_data(0) <= \R5_data[0]\;
    R6_data(31) <= \R6_data[31]\;
    R6_data(30) <= \R6_data[30]\;
    R6_data(29) <= \R6_data[29]\;
    R6_data(28) <= \R6_data[28]\;
    R6_data(27) <= \R6_data[27]\;
    R6_data(26) <= \R6_data[26]\;
    R6_data(25) <= \R6_data[25]\;
    R6_data(24) <= \R6_data[24]\;
    R6_data(23) <= \R6_data[23]\;
    R6_data(22) <= \R6_data[22]\;
    R6_data(21) <= \R6_data[21]\;
    R6_data(20) <= \R6_data[20]\;
    R6_data(19) <= \R6_data[19]\;
    R6_data(18) <= \R6_data[18]\;
    R6_data(17) <= \R6_data[17]\;
    R6_data(16) <= \R6_data[16]\;
    R6_data(15) <= \R6_data[15]\;
    R6_data(14) <= \R6_data[14]\;
    R6_data(13) <= \R6_data[13]\;
    R6_data(12) <= \R6_data[12]\;
    R6_data(11) <= \R6_data[11]\;
    R6_data(10) <= \R6_data[10]\;
    R6_data(9) <= \R6_data[9]\;
    R6_data(8) <= \R6_data[8]\;
    R6_data(7) <= \R6_data[7]\;
    R6_data(6) <= \R6_data[6]\;
    R6_data(5) <= \R6_data[5]\;
    R6_data(4) <= \R6_data[4]\;
    R6_data(3) <= \R6_data[3]\;
    R6_data(2) <= \R6_data[2]\;
    R6_data(1) <= \R6_data[1]\;
    R6_data(0) <= \R6_data[0]\;
    R7_data(31) <= \R7_data[31]\;
    R7_data(30) <= \R7_data[30]\;
    R7_data(29) <= \R7_data[29]\;
    R7_data(28) <= \R7_data[28]\;
    R7_data(27) <= \R7_data[27]\;
    R7_data(26) <= \R7_data[26]\;
    R7_data(25) <= \R7_data[25]\;
    R7_data(24) <= \R7_data[24]\;
    R7_data(23) <= \R7_data[23]\;
    R7_data(22) <= \R7_data[22]\;
    R7_data(21) <= \R7_data[21]\;
    R7_data(20) <= \R7_data[20]\;
    R7_data(19) <= \R7_data[19]\;
    R7_data(18) <= \R7_data[18]\;
    R7_data(17) <= \R7_data[17]\;
    R7_data(16) <= \R7_data[16]\;
    R7_data(15) <= \R7_data[15]\;
    R7_data(14) <= \R7_data[14]\;
    R7_data(13) <= \R7_data[13]\;
    R7_data(12) <= \R7_data[12]\;
    R7_data(11) <= \R7_data[11]\;
    R7_data(10) <= \R7_data[10]\;
    R7_data(9) <= \R7_data[9]\;
    R7_data(8) <= \R7_data[8]\;
    R7_data(7) <= \R7_data[7]\;
    R7_data(6) <= \R7_data[6]\;
    R7_data(5) <= \R7_data[5]\;
    R7_data(4) <= \R7_data[4]\;
    R7_data(3) <= \R7_data[3]\;
    R7_data(2) <= \R7_data[2]\;
    R7_data(1) <= \R7_data[1]\;
    R7_data(0) <= \R7_data[0]\;
    R0_data(31) <= \R0_data[31]\;
    R0_data(30) <= \R0_data[30]\;
    R0_data(29) <= \R0_data[29]\;
    R0_data(28) <= \R0_data[28]\;
    R0_data(27) <= \R0_data[27]\;
    R0_data(26) <= \R0_data[26]\;
    R0_data(25) <= \R0_data[25]\;
    R0_data(24) <= \R0_data[24]\;
    R0_data(23) <= \R0_data[23]\;
    R0_data(22) <= \R0_data[22]\;
    R0_data(21) <= \R0_data[21]\;
    R0_data(20) <= \R0_data[20]\;
    R0_data(19) <= \R0_data[19]\;
    R0_data(18) <= \R0_data[18]\;
    R0_data(17) <= \R0_data[17]\;
    R0_data(16) <= \R0_data[16]\;
    R0_data(15) <= \R0_data[15]\;
    R0_data(14) <= \R0_data[14]\;
    R0_data(13) <= \R0_data[13]\;
    R0_data(12) <= \R0_data[12]\;
    R0_data(11) <= \R0_data[11]\;
    R0_data(10) <= \R0_data[10]\;
    R0_data(9) <= \R0_data[9]\;
    R0_data(8) <= \R0_data[8]\;
    R0_data(7) <= \R0_data[7]\;
    R0_data(6) <= \R0_data[6]\;
    R0_data(5) <= \R0_data[5]\;
    R0_data(4) <= \R0_data[4]\;
    R0_data(3) <= \R0_data[3]\;
    R0_data(2) <= \R0_data[2]\;
    R0_data(1) <= \R0_data[1]\;
    R0_data(0) <= \R0_data[0]\;
    R4_data(31) <= \R4_data[31]\;
    R4_data(30) <= \R4_data[30]\;
    R4_data(29) <= \R4_data[29]\;
    R4_data(28) <= \R4_data[28]\;
    R4_data(27) <= \R4_data[27]\;
    R4_data(26) <= \R4_data[26]\;
    R4_data(25) <= \R4_data[25]\;
    R4_data(24) <= \R4_data[24]\;
    R4_data(23) <= \R4_data[23]\;
    R4_data(22) <= \R4_data[22]\;
    R4_data(21) <= \R4_data[21]\;
    R4_data(20) <= \R4_data[20]\;
    R4_data(19) <= \R4_data[19]\;
    R4_data(18) <= \R4_data[18]\;
    R4_data(17) <= \R4_data[17]\;
    R4_data(16) <= \R4_data[16]\;
    R4_data(15) <= \R4_data[15]\;
    R4_data(14) <= \R4_data[14]\;
    R4_data(13) <= \R4_data[13]\;
    R4_data(12) <= \R4_data[12]\;
    R4_data(11) <= \R4_data[11]\;
    R4_data(10) <= \R4_data[10]\;
    R4_data(9) <= \R4_data[9]\;
    R4_data(8) <= \R4_data[8]\;
    R4_data(7) <= \R4_data[7]\;
    R4_data(6) <= \R4_data[6]\;
    R4_data(5) <= \R4_data[5]\;
    R4_data(4) <= \R4_data[4]\;
    R4_data(3) <= \R4_data[3]\;
    R4_data(2) <= \R4_data[2]\;
    R4_data(1) <= \R4_data[1]\;
    R4_data(0) <= \R4_data[0]\;

    sum3_6_0_cry_24 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[24]\, B => \R4_data[24]\, C => 
        \R5_data[24]\, D => \R6_data[24]\, FCI => 
        \sum3_6_0_cry_23\, S => \sum3_6_0[24]\, Y => OPEN, FCO
         => \sum3_6_0_cry_24\);
    
    \next_reg_h[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(11), B => \R6_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[11]_net_1\);
    
    sum3_cry_24 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[24]\, B => Wt_data(24), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_23\, S => 
        \sum3[24]\, Y => OPEN, FCO => \sum3_cry_24\);
    
    \reg_f[12]\ : SLE
      port map(D => \next_reg_f[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[12]\);
    
    sum3_cry_30 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[30]\, B => Wt_data(30), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_29\, S => 
        \sum3[30]\, Y => OPEN, FCO => \sum3_cry_30\);
    
    \next_reg_c[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(14), B => \R1_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[14]_net_1\);
    
    \reg_f[11]\ : SLE
      port map(D => \next_reg_f[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[11]\);
    
    sum3_6_0_cry_21 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[21]\, B => \R4_data[21]\, C => 
        \R5_data[21]\, D => \R6_data[21]\, FCI => 
        \sum3_6_0_cry_20\, S => \sum3_6_0[21]\, Y => OPEN, FCO
         => \sum3_6_0_cry_21\);
    
    \reg_h[22]\ : SLE
      port map(D => \next_reg_h[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[22]\);
    
    sum0_4_cry_0 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => sum0_4_0, C => \sum0_4[0]\, D
         => GND_net_1, FCI => GND_net_1, S => OPEN, Y => 
        sum0_4_cry_0_Y_0, FCO => \sum0_4_cry_0\);
    
    \reg_e[14]\ : SLE
      port map(D => \next_reg_e[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[14]\);
    
    \reg_h[21]\ : SLE
      port map(D => \next_reg_h[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[21]\);
    
    sum3_6_cry_11 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[11]\, B => \R4_data[4]\, C => 
        \R4_data[17]\, D => \R4_data[22]\, FCI => \sum3_6_cry_10\, 
        S => \sum3_6[11]\, Y => OPEN, FCO => \sum3_6_cry_11\);
    
    \SIG0[26]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[16]\, C => 
        \R0_data[7]\, Y => \SIG0[26]_net_1\);
    
    \next_reg_f[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(9), B => \R4_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[9]_net_1\);
    
    next_reg_a_cry_23_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[23]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[23]\, D => N0_data(23), FCI => next_reg_a_cry_22, S
         => \next_reg_a[23]\, Y => OPEN, FCO => next_reg_a_cry_23);
    
    \next_reg_g[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[0]\, B => next_reg_H6_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_g[0]_net_1\);
    
    \next_reg_g[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(10), B => \R5_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[10]_net_1\);
    
    \next_reg_b[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(27), B => \R0_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[27]_net_1\);
    
    \next_reg_b[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(25), B => \R0_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[25]_net_1\);
    
    sum3_cry_26 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[26]\, B => Wt_data(26), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_25\, S => 
        \sum3[26]\, Y => OPEN, FCO => \sum3_cry_26\);
    
    \reg_d[17]\ : SLE
      port map(D => \next_reg_d[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[17]\);
    
    sum3_4_cry_5 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[5]\, B => m78, C => m83_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_4\, S => \sum3_4[5]\, Y
         => OPEN, FCO => \sum3_4_cry_5\);
    
    \reg_f[3]\ : SLE
      port map(D => \next_reg_f[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[3]\);
    
    \next_reg_f[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(27), B => \R4_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[27]_net_1\);
    
    sum0_4_cry_20 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[20]\, C => 
        \sum0_4_axb_20\, D => GND_net_1, FCI => \sum0_4_cry_19\, 
        S => \sum0_4[20]\, Y => OPEN, FCO => \sum0_4_cry_20\);
    
    sum3_6_cry_29 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[29]\, B => \R4_data[3]\, C => 
        \R4_data[8]\, D => \R4_data[22]\, FCI => \sum3_6_cry_28\, 
        S => \sum3_6[29]\, Y => OPEN, FCO => \sum3_6_cry_29\);
    
    \reg_g[13]\ : SLE
      port map(D => \next_reg_g[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[13]\);
    
    \next_reg_f[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(25), B => \R4_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[25]_net_1\);
    
    \reg_c[23]\ : SLE
      port map(D => \next_reg_c[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[23]\);
    
    next_reg_e_cry_11_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[11]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(11), D => \R3_data[11]\, FCI => next_reg_e_cry_10, 
        S => \next_reg_e[11]\, Y => OPEN, FCO => 
        next_reg_e_cry_11);
    
    \reg_f[16]\ : SLE
      port map(D => \next_reg_f[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[16]\);
    
    \next_reg_d[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(13), B => \R2_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[13]_net_1\);
    
    \reg_b[29]\ : SLE
      port map(D => \next_reg_b[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[29]\);
    
    \reg_h[26]\ : SLE
      port map(D => \next_reg_h[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[26]\);
    
    sum3_6_cry_26 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[26]\, B => \R4_data[0]\, C => 
        \R4_data[5]\, D => \R4_data[19]\, FCI => \sum3_6_cry_25\, 
        S => \sum3_6[26]\, Y => OPEN, FCO => \sum3_6_cry_26\);
    
    \reg_a[15]\ : SLE
      port map(D => \next_reg_a[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[15]\);
    
    \reg_e[22]\ : SLE
      port map(D => \next_reg_e[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[22]\);
    
    \next_reg_h[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(20), B => \R6_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[20]_net_1\);
    
    \next_reg_g[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(12), B => \R5_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[12]_net_1\);
    
    \reg_e[21]\ : SLE
      port map(D => \next_reg_e[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[21]\);
    
    \next_reg_g[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(21), B => \R5_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[21]_net_1\);
    
    next_reg_a_cry_13_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[13]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[13]\, D => N0_data(13), FCI => next_reg_a_cry_12, S
         => \next_reg_a[13]\, Y => OPEN, FCO => next_reg_a_cry_13);
    
    \reg_d[8]\ : SLE
      port map(D => \next_reg_d[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[8]\);
    
    next_reg_e_cry_18_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[18]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(18), D => \R3_data[18]\, FCI => next_reg_e_cry_17, 
        S => \next_reg_e[18]\, Y => OPEN, FCO => 
        next_reg_e_cry_18);
    
    \next_reg_c[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(8), B => \R1_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[8]_net_1\);
    
    \reg_a[25]\ : SLE
      port map(D => \next_reg_a[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[25]\);
    
    \next_reg_g[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(31), B => \R5_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[31]_net_1\);
    
    \next_reg_c[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[2]\, B => N2_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[2]_net_1\);
    
    sum3_6_0_cry_2 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[2]\, B => \R4_data[2]\, C => 
        \R5_data[2]\, D => \R6_data[2]\, FCI => \sum3_6_0_cry_1\, 
        S => \sum3_6_0[2]\, Y => OPEN, FCO => \sum3_6_0_cry_2\);
    
    \next_reg_b[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(14), B => \R0_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[14]_net_1\);
    
    sum3_6_axb_0 : CFG4
      generic map(INIT => x"6996")

      port map(A => \R4_data[25]\, B => \R4_data[11]\, C => 
        \R4_data[6]\, D => sum3_6_0_cry_0_Y, Y => \sum3_6[0]\);
    
    \next_reg_b[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(7), B => \R0_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[7]_net_1\);
    
    sum0_4_cry_23 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[23]\, C => 
        \sum0_4_axb_23\, D => GND_net_1, FCI => \sum0_4_cry_22\, 
        S => \sum0_4[23]\, Y => OPEN, FCO => \sum0_4_cry_23\);
    
    \reg_f[18]\ : SLE
      port map(D => \next_reg_f[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[18]\);
    
    \reg_b[4]\ : SLE
      port map(D => \next_reg_b[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[4]\);
    
    \next_reg_f[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(31), B => \R4_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[31]_net_1\);
    
    sum0_4_cry_0_1003 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[24]\, B => \R0_data[3]\, C => 
        \R0_data[12]\, Y => \SIG0_0[22]\);
    
    \SIG0[14]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[16]\, C => 
        \R0_data[4]\, Y => \SIG0[14]_net_1\);
    
    \reg_h[28]\ : SLE
      port map(D => \next_reg_h[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[28]\);
    
    \reg_b[7]\ : SLE
      port map(D => \next_reg_b[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[7]\);
    
    sum0_4_cry_17 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[17]\, C => 
        \sum0_4_axb_17\, D => GND_net_1, FCI => \sum0_4_cry_16\, 
        S => \sum0_4[17]\, Y => OPEN, FCO => \sum0_4_cry_17\);
    
    \reg_g[14]\ : SLE
      port map(D => \next_reg_g[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[14]\);
    
    sum0_4_cry_0_1020 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[18]\, C => 
        \R0_data[7]\, Y => \SIG0_0[5]\);
    
    \reg_c[24]\ : SLE
      port map(D => \next_reg_c[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[24]\);
    
    \next_reg_b[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(9), B => \R0_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[9]_net_1\);
    
    sum0_4_cry_0_996 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[19]\, C => 
        \R0_data[10]\, Y => \SIG0_0[29]\);
    
    \reg_h[15]\ : SLE
      port map(D => \next_reg_h[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[15]\);
    
    next_reg_e_cry_3_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[3]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(3), D => \R3_data[3]\, FCI => next_reg_e_cry_2, S
         => \next_reg_e[3]\, Y => OPEN, FCO => next_reg_e_cry_3);
    
    sum0_4_cry_0_1010 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[17]\, C => 
        \R0_data[5]\, Y => \SIG0_0[15]\);
    
    \next_reg_h[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(22), B => \R6_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[22]_net_1\);
    
    sum0_4_cry_28 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[28]\, C => 
        \sum0_4_axb_28\, D => GND_net_1, FCI => \sum0_4_cry_27\, 
        S => \sum0_4[28]\, Y => OPEN, FCO => \sum0_4_cry_28\);
    
    \reg_f[23]\ : SLE
      port map(D => \next_reg_f[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[23]\);
    
    \reg_e[26]\ : SLE
      port map(D => \next_reg_e[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[26]\);
    
    sum3_6_cry_8 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[8]\, B => \R4_data[1]\, C => 
        \R4_data[14]\, D => \R4_data[19]\, FCI => \sum3_6_cry_7\, 
        S => \sum3_6[8]\, Y => OPEN, FCO => \sum3_6_cry_8\);
    
    sum0_4_cry_0_1008 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[19]\, C => 
        \R0_data[7]\, Y => \SIG0_0[17]\);
    
    sum3_6_cry_22 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[22]\, B => \R4_data[1]\, C => 
        \R4_data[15]\, D => \R4_data[28]\, FCI => \sum3_6_cry_21\, 
        S => \sum3_6[22]\, Y => OPEN, FCO => \sum3_6_cry_22\);
    
    \reg_e[9]\ : SLE
      port map(D => \next_reg_e[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[9]\);
    
    \reg_g[9]\ : SLE
      port map(D => \next_reg_g[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[9]\);
    
    \reg_d[22]\ : SLE
      port map(D => \next_reg_d[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[22]\);
    
    \next_reg_d[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(7), B => \R2_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[7]_net_1\);
    
    \next_reg_c[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(7), B => \R1_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[7]_net_1\);
    
    \reg_d[21]\ : SLE
      port map(D => \next_reg_d[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[21]\);
    
    sum3_4_cry_11 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[11]\, B => m141, C => m144_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_10\, S => \sum3_4[11]\, Y
         => OPEN, FCO => \sum3_4_cry_11\);
    
    \next_reg_c[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(17), B => \R1_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[17]_net_1\);
    
    \next_reg_h[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(31), B => \R6_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[31]_net_1\);
    
    \next_reg_c[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(15), B => \R1_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[15]_net_1\);
    
    \next_reg_b[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(20), B => \R0_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[20]_net_1\);
    
    \reg_e[19]\ : SLE
      port map(D => \next_reg_e[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[19]\);
    
    sum3_cry_10 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[10]\, B => Wt_data(10), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_9\, S => 
        \sum3[10]\, Y => OPEN, FCO => \sum3_cry_10\);
    
    sum3_cry_2 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[2]\, B => Wt_data(2), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_1\, S => \sum3[2]\, Y
         => OPEN, FCO => \sum3_cry_2\);
    
    \next_reg_d[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(18), B => \R2_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[18]_net_1\);
    
    \reg_e[28]\ : SLE
      port map(D => \next_reg_e[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[28]\);
    
    sum3_cry_27 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[27]\, B => Wt_data(27), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_26\, S => 
        \sum3[27]\, Y => OPEN, FCO => \sum3_cry_27\);
    
    \reg_e[8]\ : SLE
      port map(D => \next_reg_e[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[8]\);
    
    sum0_4_cry_0_1002 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[13]\, C => 
        \R0_data[4]\, Y => \SIG0_0[23]\);
    
    \next_reg_d[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[0]\, B => next_reg_H3_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_d[0]_net_1\);
    
    \next_reg_f[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(20), B => \R4_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[20]_net_1\);
    
    \reg_b[27]\ : SLE
      port map(D => \next_reg_b[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[27]\);
    
    \next_reg_h[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(9), B => \R6_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[9]_net_1\);
    
    \next_reg_b[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[0]\, B => next_reg_H1_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_b[0]_net_1\);
    
    \reg_b[13]\ : SLE
      port map(D => \next_reg_b[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[13]\);
    
    \reg_e[31]\ : SLE
      port map(D => \next_reg_e[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[31]\);
    
    sum3_6_0_cry_30 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[30]\, B => \R4_data[30]\, C => 
        \R5_data[30]\, D => \R6_data[30]\, FCI => 
        \sum3_6_0_cry_29\, S => \sum3_6_0[30]\, Y => OPEN, FCO
         => \sum3_6_0_cry_30\);
    
    sum3_6_0_cry_13 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[13]\, B => \R4_data[13]\, C => 
        \R5_data[13]\, D => \R6_data[13]\, FCI => 
        \sum3_6_0_cry_12\, S => \sum3_6_0[13]\, Y => OPEN, FCO
         => \sum3_6_0_cry_13\);
    
    \reg_f[24]\ : SLE
      port map(D => \next_reg_f[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[24]\);
    
    \next_reg_d[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(29), B => \R2_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[29]_net_1\);
    
    \next_reg_f[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(11), B => \R4_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[11]_net_1\);
    
    \SIG0[15]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[17]\, C => 
        \R0_data[5]\, Y => \SIG0[15]_net_1\);
    
    \reg_a[10]\ : SLE
      port map(D => \next_reg_a[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[10]\);
    
    \next_reg_f[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[6]\, B => N5_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[6]_net_1\);
    
    \reg_d[9]\ : SLE
      port map(D => \next_reg_d[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[9]\);
    
    \reg_d[26]\ : SLE
      port map(D => \next_reg_d[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[26]\);
    
    \reg_a[20]\ : SLE
      port map(D => \next_reg_a[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[20]\);
    
    \next_reg_b[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(22), B => \R0_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[22]_net_1\);
    
    \next_reg_c[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(24), B => \R1_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[24]_net_1\);
    
    sum0_4_cry_0_1021 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[17]\, C => 
        \R0_data[6]\, Y => \SIG0_0[4]\);
    
    \reg_f[1]\ : SLE
      port map(D => \next_reg_f[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[1]\);
    
    sum0_4_cry_0_1011 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[16]\, C => 
        \R0_data[4]\, Y => \SIG0_0[14]\);
    
    sum3_6_0_cry_25 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[25]\, B => \R4_data[25]\, C => 
        \R5_data[25]\, D => \R6_data[25]\, FCI => 
        \sum3_6_0_cry_24\, S => \sum3_6_0[25]\, Y => OPEN, FCO
         => \sum3_6_0_cry_25\);
    
    sum3_4_cry_4 : ARI1
      generic map(INIT => x"5C53A")

      port map(A => \sum3_6[4]\, B => m67_ns, C => m73, D => 
        Kt_addr(5), FCI => \sum3_4_cry_3\, S => \sum3_4[4]\, Y
         => OPEN, FCO => \sum3_4_cry_4\);
    
    \next_reg_f[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(22), B => \R4_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[22]_net_1\);
    
    sum0_4_axb_28 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[28]\, B => \R1_data[28]\, C => 
        \R0_data[28]\, D => \SIG0[28]_net_1\, Y => 
        \sum0_4_axb_28\);
    
    sum0_4_cry_14 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[14]\, C => 
        \sum0_4_axb_14\, D => GND_net_1, FCI => \sum0_4_cry_13\, 
        S => \sum0_4[14]\, Y => OPEN, FCO => \sum0_4_cry_14\);
    
    sum3_6_cry_30 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[30]\, B => \R4_data[4]\, C => 
        \R4_data[9]\, D => \R4_data[23]\, FCI => \sum3_6_cry_29\, 
        S => \sum3_6[30]\, Y => OPEN, FCO => \sum3_6_cry_30\);
    
    \next_reg_b[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(17), B => \R0_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[17]_net_1\);
    
    \reg_a[0]\ : SLE
      port map(D => next_reg_a_cry_0_0_Y, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[0]\);
    
    \reg_h[10]\ : SLE
      port map(D => \next_reg_h[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[10]\);
    
    \reg_b[14]\ : SLE
      port map(D => \next_reg_b[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[14]\);
    
    \next_reg_b[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(15), B => \R0_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[15]_net_1\);
    
    sum3_6_cry_10 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[10]\, B => \R4_data[3]\, C => 
        \R4_data[16]\, D => \R4_data[21]\, FCI => \sum3_6_cry_9\, 
        S => \sum3_6[10]\, Y => OPEN, FCO => \sum3_6_cry_10\);
    
    \reg_d[28]\ : SLE
      port map(D => \next_reg_d[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[28]\);
    
    \reg_d[2]\ : SLE
      port map(D => \next_reg_d[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[2]\);
    
    next_reg_e_cry_26_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[26]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(26), D => \R3_data[26]\, FCI => next_reg_e_cry_25, 
        S => \next_reg_e[26]\, Y => OPEN, FCO => 
        next_reg_e_cry_26);
    
    \reg_f[4]\ : SLE
      port map(D => \next_reg_f[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[4]\);
    
    \next_reg_c[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[5]\, B => N2_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[5]_net_1\);
    
    sum3_4_cry_0_993 : CFG4
      generic map(INIT => x"C1CD")

      port map(A => m10_bm, B => m20_1, C => Kt_addr(5), D => 
        m10_am, Y => \Kt_data_0[0]\);
    
    \reg_f[9]\ : SLE
      port map(D => \next_reg_f[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[9]\);
    
    sum3_4_cry_27 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[27]\, B => m289, C => m292_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_26\, S => \sum3_4[27]\, Y
         => OPEN, FCO => \sum3_4_cry_27\);
    
    sum3_6_0_cry_6 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[6]\, B => \R4_data[6]\, C => 
        \R5_data[6]\, D => \R6_data[6]\, FCI => \sum3_6_0_cry_5\, 
        S => \sum3_6_0[6]\, Y => OPEN, FCO => \sum3_6_0_cry_6\);
    
    \reg_g[19]\ : SLE
      port map(D => \next_reg_g[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[19]\);
    
    \next_reg_d[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(16), B => \R2_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[16]_net_1\);
    
    \next_reg_c[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[4]\, B => N2_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[4]_net_1\);
    
    \reg_c[29]\ : SLE
      port map(D => \next_reg_c[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[29]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \next_reg_g[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(8), B => \R5_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[8]_net_1\);
    
    sum0_4_cry_29 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[29]\, C => 
        \sum0_4_axb_29\, D => GND_net_1, FCI => \sum0_4_cry_28\, 
        S => \sum0_4[29]\, Y => OPEN, FCO => \sum0_4_cry_29\);
    
    \next_reg_g[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(11), B => \R5_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[11]_net_1\);
    
    \reg_e[17]\ : SLE
      port map(D => \next_reg_e[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[17]\);
    
    \reg_g[1]\ : SLE
      port map(D => \next_reg_g[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[1]\);
    
    \next_reg_b[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[3]\, B => N1_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[3]_net_1\);
    
    sum3_cry_0_994 : CFG4
      generic map(INIT => x"A3A0")

      port map(A => next_r0_0_cry_0_Y, B => W_out_i_0(0), C => 
        ld_i_i_3, D => N_98, Y => \Wt_data_0[0]\);
    
    sum3_cry_19 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[19]\, B => Wt_data(19), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_18\, S => 
        \sum3[19]\, Y => OPEN, FCO => \sum3_cry_19\);
    
    sum0_4_cry_26 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[26]\, C => 
        \sum0_4_axb_26\, D => GND_net_1, FCI => \sum0_4_cry_25\, 
        S => \sum0_4[26]\, Y => OPEN, FCO => \sum0_4_cry_26\);
    
    \next_reg_c[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(10), B => \R1_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[10]_net_1\);
    
    sum3_cry_18 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[18]\, B => Wt_data(18), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_17\, S => 
        \sum3[18]\, Y => OPEN, FCO => \sum3_cry_18\);
    
    \reg_a[31]\ : SLE
      port map(D => \next_reg_a[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[31]\);
    
    \next_reg_h[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(13), B => \R6_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[13]_net_1\);
    
    sum3_6_cry_13 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[13]\, B => \R4_data[6]\, C => 
        \R4_data[19]\, D => \R4_data[24]\, FCI => \sum3_6_cry_12\, 
        S => \sum3_6[13]\, Y => OPEN, FCO => \sum3_6_cry_13\);
    
    sum0_4_cry_0_1004 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[11]\, C => 
        \R0_data[2]\, Y => \SIG0_0[21]\);
    
    sum0_4_axb_6 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[6]\, B => \R1_data[6]\, C => 
        \R0_data[6]\, D => \SIG0[6]_net_1\, Y => \sum0_4_axb_6\);
    
    \reg_g[25]\ : SLE
      port map(D => \next_reg_g[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[25]\);
    
    \next_reg_h[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(21), B => \R6_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[21]_net_1\);
    
    sum3_6_cry_18 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[18]\, B => \R4_data[11]\, C => 
        \R4_data[24]\, D => \R4_data[29]\, FCI => \sum3_6_cry_17\, 
        S => \sum3_6[18]\, Y => OPEN, FCO => \sum3_6_cry_18\);
    
    \reg_h[0]\ : SLE
      port map(D => \next_reg_h[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[0]\);
    
    sum3_4_cry_6 : ARI1
      generic map(INIT => x"53AC5")

      port map(A => \sum3_6[6]\, B => m95_1_0, C => m95_1_1, D
         => Kt_addr_5_rep1, FCI => \sum3_4_cry_5\, S => 
        \sum3_4[6]\, Y => OPEN, FCO => \sum3_4_cry_6\);
    
    \reg_c[31]\ : SLE
      port map(D => \next_reg_c[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[31]\);
    
    \next_reg_c[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(12), B => \R1_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[12]_net_1\);
    
    \reg_f[29]\ : SLE
      port map(D => \next_reg_f[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[29]\);
    
    next_reg_e_cry_21_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[21]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(21), D => \R3_data[21]\, FCI => next_reg_e_cry_20, 
        S => \next_reg_e[21]\, Y => OPEN, FCO => 
        next_reg_e_cry_21);
    
    sum3_6_cry_4 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[4]\, B => \R4_data[10]\, C => 
        \R4_data[15]\, D => \R4_data[29]\, FCI => \sum3_6_cry_3\, 
        S => \sum3_6[4]\, Y => OPEN, FCO => \sum3_6_cry_4\);
    
    sum0_4_cry_22 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[22]\, C => 
        \sum0_4_axb_22\, D => GND_net_1, FCI => \sum0_4_cry_21\, 
        S => \sum0_4[22]\, Y => OPEN, FCO => \sum0_4_cry_22\);
    
    \next_reg_c[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(27), B => \R1_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[27]_net_1\);
    
    sum3_cry_7 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[7]\, B => Wt_data(7), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_6\, S => \sum3[7]\, Y
         => OPEN, FCO => \sum3_cry_7\);
    
    \reg_g[6]\ : SLE
      port map(D => \next_reg_g[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[6]\);
    
    \next_reg_c[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(25), B => \R1_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[25]_net_1\);
    
    next_reg_e_cry_28_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[28]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(28), D => \R3_data[28]\, FCI => next_reg_e_cry_27, 
        S => \next_reg_e[28]\, Y => OPEN, FCO => 
        next_reg_e_cry_28);
    
    \next_reg_g[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(23), B => \R5_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[23]_net_1\);
    
    \next_reg_b[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(10), B => \R0_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[10]_net_1\);
    
    \SIG0[12]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[14]\, C => 
        \R0_data[2]\, Y => \SIG0[12]_net_1\);
    
    \reg_g[17]\ : SLE
      port map(D => \next_reg_g[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[17]\);
    
    \reg_c[27]\ : SLE
      port map(D => \next_reg_c[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[27]\);
    
    sum3_4_cry_24 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_6[24]\, B => Kt_data_24, C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_4_cry_23\, S => \sum3_4[24]\, 
        Y => OPEN, FCO => \sum3_4_cry_24\);
    
    \reg_d[0]\ : SLE
      port map(D => \next_reg_d[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[0]\);
    
    sum3_4_cry_10 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[10]\, B => m137_am, C => m137_bm, D
         => Kt_addr_5_rep1, FCI => \sum3_4_cry_9\, S => 
        \sum3_4[10]\, Y => OPEN, FCO => \sum3_4_cry_10\);
    
    \next_reg_d[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[2]\, B => N3_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[2]_net_1\);
    
    \reg_a[13]\ : SLE
      port map(D => \next_reg_a[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[13]\);
    
    sum0_4_cry_0_1009 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[18]\, C => 
        \R0_data[6]\, Y => \SIG0_0[16]\);
    
    \reg_h[4]\ : SLE
      port map(D => \next_reg_h[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[4]\);
    
    \reg_b[19]\ : SLE
      port map(D => \next_reg_b[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[19]\);
    
    \next_reg_h[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[6]\, B => N7_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[6]_net_1\);
    
    \next_reg_h[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(18), B => \R6_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[18]_net_1\);
    
    \reg_a[23]\ : SLE
      port map(D => \next_reg_a[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[23]\);
    
    sum3_cry_15 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[15]\, B => Wt_data(15), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_14\, S => 
        \sum3[15]\, Y => OPEN, FCO => \sum3_cry_15\);
    
    \next_reg_b[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(21), B => \R0_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[21]_net_1\);
    
    sum3_6_0_cry_28 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[28]\, B => \R4_data[28]\, C => 
        \R5_data[28]\, D => \R6_data[28]\, FCI => 
        \sum3_6_0_cry_27\, S => \sum3_6_0[28]\, Y => OPEN, FCO
         => \sum3_6_0_cry_28\);
    
    \reg_b[5]\ : SLE
      port map(D => \next_reg_b[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[5]\);
    
    \reg_b[3]\ : SLE
      port map(D => \next_reg_b[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[3]\);
    
    next_reg_a_cry_26_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[26]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[26]\, D => N0_data(26), FCI => next_reg_a_cry_25, S
         => \next_reg_a[26]\, Y => OPEN, FCO => next_reg_a_cry_26);
    
    sum3_6_cry_5 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[5]\, B => \R4_data[11]\, C => 
        \R4_data[16]\, D => \R4_data[30]\, FCI => \sum3_6_cry_4\, 
        S => \sum3_6[5]\, Y => OPEN, FCO => \sum3_6_cry_5\);
    
    \SIG0[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[22]\, B => \R0_data[13]\, C => 
        \R0_data[2]\, Y => sum0_4);
    
    \next_reg_b[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(12), B => \R0_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[12]_net_1\);
    
    \next_reg_f[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(21), B => \R4_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[21]_net_1\);
    
    sum3_6_cry_27 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[27]\, B => \R4_data[1]\, C => 
        \R4_data[6]\, D => \R4_data[20]\, FCI => \sum3_6_cry_26\, 
        S => \sum3_6[27]\, Y => OPEN, FCO => \sum3_6_cry_27\);
    
    \next_reg_d[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(24), B => \R2_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[24]_net_1\);
    
    sum3_4_cry_13 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[13]\, B => m168_1_0, C => m168_1_1, D
         => Kt_addr(5), FCI => \sum3_4_cry_12\, S => \sum3_4[13]\, 
        Y => OPEN, FCO => \sum3_4_cry_13\);
    
    sum3_6_0_cry_10 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[10]\, B => \R4_data[10]\, C => 
        \R5_data[10]\, D => \R6_data[10]\, FCI => 
        \sum3_6_0_cry_9\, S => \sum3_6_0[10]\, Y => OPEN, FCO => 
        \sum3_6_0_cry_10\);
    
    \reg_h[13]\ : SLE
      port map(D => \next_reg_h[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[13]\);
    
    \reg_g[20]\ : SLE
      port map(D => \next_reg_g[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[20]\);
    
    sum3_6_0_cry_16 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[16]\, B => \R4_data[16]\, C => 
        \R5_data[16]\, D => \R6_data[16]\, FCI => 
        \sum3_6_0_cry_15\, S => \sum3_6_0[16]\, Y => OPEN, FCO
         => \sum3_6_0_cry_16\);
    
    \SIG0[30]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[20]\, B => \R0_data[11]\, C => 
        \R0_data[0]\, Y => \SIG0[30]_net_1\);
    
    sum3_6_0_cry_3 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[3]\, B => \R4_data[3]\, C => 
        \R5_data[3]\, D => \R6_data[3]\, FCI => \sum3_6_0_cry_2\, 
        S => \sum3_6_0[3]\, Y => OPEN, FCO => \sum3_6_0_cry_3\);
    
    \reg_a[14]\ : SLE
      port map(D => \next_reg_a[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[14]\);
    
    \reg_e[5]\ : SLE
      port map(D => \next_reg_e[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[5]\);
    
    \reg_f[27]\ : SLE
      port map(D => \next_reg_f[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[27]\);
    
    \reg_c[12]\ : SLE
      port map(D => \next_reg_c[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[12]\);
    
    \reg_f[15]\ : SLE
      port map(D => \next_reg_f[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[15]\);
    
    \reg_c[11]\ : SLE
      port map(D => \next_reg_c[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[11]\);
    
    sum3_4_cry_18 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[18]\, B => m215_am, C => m215_bm, D
         => Kt_addr(5), FCI => \sum3_4_cry_17\, S => \sum3_4[18]\, 
        Y => OPEN, FCO => \sum3_4_cry_18\);
    
    \SIG0[16]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[18]\, C => 
        \R0_data[6]\, Y => \SIG0[16]_net_1\);
    
    \reg_h[25]\ : SLE
      port map(D => \next_reg_h[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[25]\);
    
    sum3_6_cry_19 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[19]\, B => \R4_data[12]\, C => 
        \R4_data[25]\, D => \R4_data[30]\, FCI => \sum3_6_cry_18\, 
        S => \sum3_6[19]\, Y => OPEN, FCO => \sum3_6_cry_19\);
    
    \reg_b[2]\ : SLE
      port map(D => \next_reg_b[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[2]\);
    
    \reg_a[24]\ : SLE
      port map(D => \next_reg_a[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[24]\);
    
    sum3_cry_22 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[22]\, B => Wt_data(22), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_21\, S => 
        \sum3[22]\, Y => OPEN, FCO => \sum3_cry_22\);
    
    next_reg_e_cry_12_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[12]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(12), D => \R3_data[12]\, FCI => next_reg_e_cry_11, 
        S => \next_reg_e[12]\, Y => OPEN, FCO => 
        next_reg_e_cry_12);
    
    \next_reg_f[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[0]\, B => next_reg_H5_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_f[0]_net_1\);
    
    next_reg_a_cry_16_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[16]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[16]\, D => N0_data(16), FCI => next_reg_a_cry_15, S
         => \next_reg_a[16]\, Y => OPEN, FCO => next_reg_a_cry_16);
    
    \next_reg_g[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(28), B => \R5_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[28]_net_1\);
    
    sum3_6_cry_16 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[16]\, B => \R4_data[9]\, C => 
        \R4_data[22]\, D => \R4_data[27]\, FCI => \sum3_6_cry_15\, 
        S => \sum3_6[16]\, Y => OPEN, FCO => \sum3_6_cry_16\);
    
    \next_reg_d[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[1]\, B => N3_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[1]_net_1\);
    
    \next_reg_f[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(13), B => \R4_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[13]_net_1\);
    
    next_reg_e_cry_4_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[4]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(4), D => \R3_data[4]\, FCI => next_reg_e_cry_3, S
         => \next_reg_e[4]\, Y => OPEN, FCO => next_reg_e_cry_4);
    
    \reg_f[2]\ : SLE
      port map(D => \next_reg_f[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[2]\);
    
    \next_reg_h[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(16), B => \R6_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[16]_net_1\);
    
    sum0_4_cry_1 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[1]\, C => 
        \sum0_4_axb_1\, D => GND_net_1, FCI => \sum0_4_cry_0\, S
         => \sum0_4[1]\, Y => OPEN, FCO => \sum0_4_cry_1\);
    
    \next_reg_c[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(20), B => \R1_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[20]_net_1\);
    
    sum0_4_cry_15 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[15]\, C => 
        \sum0_4_axb_15\, D => GND_net_1, FCI => \sum0_4_cry_14\, 
        S => \sum0_4[15]\, Y => OPEN, FCO => \sum0_4_cry_15\);
    
    \next_reg_b[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[5]\, B => N1_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[5]_net_1\);
    
    \reg_h[14]\ : SLE
      port map(D => \next_reg_h[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[14]\);
    
    next_reg_e_cry_9_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[9]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(9), D => \R3_data[9]\, FCI => next_reg_e_cry_8, S
         => \next_reg_e[9]\, Y => OPEN, FCO => next_reg_e_cry_9);
    
    \reg_b[17]\ : SLE
      port map(D => \next_reg_b[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[17]\);
    
    \SIG0[29]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[19]\, C => 
        \R0_data[10]\, Y => \SIG0[29]_net_1\);
    
    next_reg_a_cry_21_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[21]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[21]\, D => N0_data(21), FCI => next_reg_a_cry_20, S
         => \next_reg_a[21]\, Y => OPEN, FCO => next_reg_a_cry_21);
    
    \reg_c[16]\ : SLE
      port map(D => \next_reg_c[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[16]\);
    
    sum0_4_cry_7 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[7]\, C => 
        \sum0_4_axb_7\, D => GND_net_1, FCI => \sum0_4_cry_6\, S
         => \sum0_4[7]\, Y => OPEN, FCO => \sum0_4_cry_7\);
    
    \reg_h[8]\ : SLE
      port map(D => \next_reg_h[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[8]\);
    
    next_reg_a_cry_4_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[4]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[4]\, D => N0_data(4), FCI => next_reg_a_cry_3, S
         => \next_reg_a[4]\, Y => OPEN, FCO => next_reg_a_cry_4);
    
    \reg_e[25]\ : SLE
      port map(D => \next_reg_e[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[25]\);
    
    \reg_a[8]\ : SLE
      port map(D => \next_reg_a[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[8]\);
    
    sum3_cry_14 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[14]\, B => Wt_data(14), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_13\, S => 
        \sum3[14]\, Y => OPEN, FCO => \sum3_cry_14\);
    
    \next_reg_c[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(11), B => \R1_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[11]_net_1\);
    
    sum3_cry_3 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[3]\, B => Wt_data(3), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_2\, S => \sum3[3]\, Y
         => OPEN, FCO => \sum3_cry_3\);
    
    sum0_4_cry_0_1007 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[20]\, C => 
        \R0_data[8]\, Y => \SIG0_0[18]\);
    
    next_reg_a_cry_28_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[28]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[28]\, D => N0_data(28), FCI => next_reg_a_cry_27, S
         => \next_reg_a[28]\, Y => OPEN, FCO => next_reg_a_cry_28);
    
    \next_reg_c[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(22), B => \R1_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[22]_net_1\);
    
    sum0_4_axb_18 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[18]\, B => \R1_data[18]\, C => 
        \R0_data[18]\, D => \SIG0[18]_net_1\, Y => 
        \sum0_4_axb_18\);
    
    \next_reg_h[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(8), B => \R6_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[8]_net_1\);
    
    \reg_f[30]\ : SLE
      port map(D => \next_reg_f[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[30]\);
    
    sum3_6_cry_24 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[24]\, B => \R4_data[3]\, C => 
        \R4_data[17]\, D => \R4_data[30]\, FCI => \sum3_6_cry_23\, 
        S => \sum3_6[24]\, Y => OPEN, FCO => \sum3_6_cry_24\);
    
    sum3_6_cry_12 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[12]\, B => \R4_data[5]\, C => 
        \R4_data[18]\, D => \R4_data[23]\, FCI => \sum3_6_cry_11\, 
        S => \sum3_6[12]\, Y => OPEN, FCO => \sum3_6_cry_12\);
    
    \reg_c[18]\ : SLE
      port map(D => \next_reg_c[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[18]\);
    
    next_reg_e_cry_5_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[5]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(5), D => \R3_data[5]\, FCI => next_reg_e_cry_4, S
         => \next_reg_e[5]\, Y => OPEN, FCO => next_reg_e_cry_5);
    
    sum3_6_0_s_31 : ARI1
      generic map(INIT => x"427D8")

      port map(A => \R7_data[31]\, B => \R4_data[31]\, C => 
        \R5_data[31]\, D => \R6_data[31]\, FCI => 
        \sum3_6_0_cry_30\, S => \sum3_6_0[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_e_cry_8_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[8]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(8), D => \R3_data[8]\, FCI => next_reg_e_cry_7, S
         => \next_reg_e[8]\, Y => OPEN, FCO => next_reg_e_cry_8);
    
    \next_reg_g[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[1]\, B => N6_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[1]_net_1\);
    
    \next_reg_g[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(13), B => \R5_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[13]_net_1\);
    
    \next_reg_g[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(26), B => \R5_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[26]_net_1\);
    
    \reg_b[6]\ : SLE
      port map(D => \next_reg_b[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[6]\);
    
    sum3_cry_16 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[16]\, B => Wt_data(16), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_15\, S => 
        \sum3[16]\, Y => OPEN, FCO => \sum3_cry_16\);
    
    \next_reg_d[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(27), B => \R2_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[27]_net_1\);
    
    sum3_6_cry_6 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[6]\, B => \R4_data[12]\, C => 
        \R4_data[17]\, D => \R4_data[31]\, FCI => \sum3_6_cry_5\, 
        S => \sum3_6[6]\, Y => OPEN, FCO => \sum3_6_cry_6\);
    
    next_reg_a_cry_11_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[11]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[11]\, D => N0_data(11), FCI => next_reg_a_cry_10, S
         => \next_reg_a[11]\, Y => OPEN, FCO => next_reg_a_cry_11);
    
    sum0_4_s_31 : ARI1
      generic map(INIT => x"46996")

      port map(A => \R0_data[21]\, B => \Maj[31]_net_1\, C => 
        \R0_data[1]\, D => \R0_data[12]\, FCI => \sum0_4_cry_30\, 
        S => \sum0_4[31]\, Y => OPEN, FCO => OPEN);
    
    \next_reg_d[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(25), B => \R2_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[25]_net_1\);
    
    \reg_f[10]\ : SLE
      port map(D => \next_reg_f[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[10]\);
    
    \reg_h[20]\ : SLE
      port map(D => \next_reg_h[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[20]\);
    
    \reg_d[12]\ : SLE
      port map(D => \next_reg_d[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[12]\);
    
    \next_reg_h[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[5]\, B => N7_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[5]_net_1\);
    
    sum0_4_cry_6 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[6]\, C => 
        \sum0_4_axb_6\, D => GND_net_1, FCI => \sum0_4_cry_5\, S
         => \sum0_4[6]\, Y => OPEN, FCO => \sum0_4_cry_6\);
    
    \reg_d[11]\ : SLE
      port map(D => \next_reg_d[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[11]\);
    
    \reg_c[2]\ : SLE
      port map(D => \next_reg_c[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[2]\);
    
    \next_reg_f[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(18), B => \R4_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[18]_net_1\);
    
    next_reg_a_cry_7_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[7]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[7]\, D => N0_data(7), FCI => next_reg_a_cry_6, S
         => \next_reg_a[7]\, Y => OPEN, FCO => next_reg_a_cry_7);
    
    \reg_d[25]\ : SLE
      port map(D => \next_reg_d[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[25]\);
    
    sum3_6_0_cry_22 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[22]\, B => \R4_data[22]\, C => 
        \R5_data[22]\, D => \R6_data[22]\, FCI => 
        \sum3_6_0_cry_21\, S => \sum3_6_0[22]\, Y => OPEN, FCO
         => \sum3_6_0_cry_22\);
    
    \reg_a[19]\ : SLE
      port map(D => \next_reg_a[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[19]\);
    
    sum3_4_cry_19 : ARI1
      generic map(INIT => x"53AC5")

      port map(A => \sum3_6[19]\, B => m219, C => m222_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_18\, S => \sum3_4[19]\, Y
         => OPEN, FCO => \sum3_4_cry_19\);
    
    next_reg_a_cry_18_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[18]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[18]\, D => N0_data(18), FCI => next_reg_a_cry_17, S
         => \next_reg_a[18]\, Y => OPEN, FCO => next_reg_a_cry_18);
    
    next_reg_e_cry_15_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[15]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(15), D => \R3_data[15]\, FCI => next_reg_e_cry_14, 
        S => \next_reg_e[15]\, Y => OPEN, FCO => 
        next_reg_e_cry_15);
    
    sum3_6_0_cry_14 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[14]\, B => \R4_data[14]\, C => 
        \R5_data[14]\, D => \R6_data[14]\, FCI => 
        \sum3_6_0_cry_13\, S => \sum3_6_0[14]\, Y => OPEN, FCO
         => \sum3_6_0_cry_14\);
    
    \next_reg_h[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(23), B => \R6_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[23]_net_1\);
    
    \reg_f[7]\ : SLE
      port map(D => \next_reg_f[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[7]\);
    
    \reg_a[29]\ : SLE
      port map(D => \next_reg_a[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[29]\);
    
    \next_reg_b[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(11), B => \R0_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[11]_net_1\);
    
    \reg_e[0]\ : SLE
      port map(D => next_reg_e_cry_0_0_Y, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[0]\);
    
    \SIG0[7]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[20]\, C => 
        \R0_data[9]\, Y => \SIG0[7]_net_1\);
    
    sum3_4_cry_16 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[16]\, B => m197_1_0, C => m197_1_1, D
         => Kt_addr(5), FCI => \sum3_4_cry_15\, S => \sum3_4[16]\, 
        Y => OPEN, FCO => \sum3_4_cry_16\);
    
    sum3_6_0_cry_11 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[11]\, B => \R4_data[11]\, C => 
        \R5_data[11]\, D => \R6_data[11]\, FCI => 
        \sum3_6_0_cry_10\, S => \sum3_6_0[11]\, Y => OPEN, FCO
         => \sum3_6_0_cry_11\);
    
    \next_reg_g[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[6]\, B => N6_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[6]_net_1\);
    
    \reg_e[1]\ : SLE
      port map(D => \next_reg_e[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[1]\);
    
    \SIG0[23]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[13]\, C => 
        \R0_data[4]\, Y => \SIG0[23]_net_1\);
    
    \reg_g[23]\ : SLE
      port map(D => \next_reg_g[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[23]\);
    
    sum3_6_0_cry_5 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[5]\, B => \R4_data[5]\, C => 
        \R5_data[5]\, D => \R6_data[5]\, FCI => \sum3_6_0_cry_4\, 
        S => \sum3_6_0[5]\, Y => OPEN, FCO => \sum3_6_0_cry_5\);
    
    sum3_4_cry_2 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[2]\, B => m49_am, C => m49_bm, D => 
        Kt_addr_5_rep1, FCI => \sum3_4_cry_1\, S => \sum3_4[2]\, 
        Y => OPEN, FCO => \sum3_4_cry_2\);
    
    sum3_4_cry_25 : ARI1
      generic map(INIT => x"5C53A")

      port map(A => \sum3_6[25]\, B => m273, C => m276_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_24\, S => \sum3_4[25]\, Y
         => OPEN, FCO => \sum3_4_cry_25\);
    
    \next_reg_d[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(19), B => \R2_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[19]_net_1\);
    
    \reg_d[16]\ : SLE
      port map(D => \next_reg_d[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[16]\);
    
    sum0_4_cry_27 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[27]\, C => 
        \sum0_4_axb_27\, D => GND_net_1, FCI => \sum0_4_cry_26\, 
        S => \sum0_4[27]\, Y => OPEN, FCO => \sum0_4_cry_27\);
    
    sum3_4_cry_30 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \sum3_6[30]\, B => m316, C => GND_net_1, D
         => GND_net_1, FCI => \sum3_4_cry_29\, S => \sum3_4[30]\, 
        Y => OPEN, FCO => \sum3_4_cry_30\);
    
    \reg_h[19]\ : SLE
      port map(D => \next_reg_h[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[19]\);
    
    \reg_e[20]\ : SLE
      port map(D => \next_reg_e[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[20]\);
    
    \reg_c[4]\ : SLE
      port map(D => \next_reg_c[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[4]\);
    
    sum0_4_cry_0_1025 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[22]\, B => \R0_data[13]\, C => 
        \R0_data[2]\, Y => sum0_4_0);
    
    sum0_4_axb_26 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[26]\, B => \R1_data[26]\, C => 
        \R0_data[26]\, D => \SIG0[26]_net_1\, Y => 
        \sum0_4_axb_26\);
    
    \reg_a[2]\ : SLE
      port map(D => \next_reg_a[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[2]\);
    
    sum0_4_cry_4 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[4]\, C => 
        \sum0_4_axb_4\, D => GND_net_1, FCI => \sum0_4_cry_3\, S
         => \sum0_4[4]\, Y => OPEN, FCO => \sum0_4_cry_4\);
    
    \next_reg_b[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[1]\, B => N1_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[1]_net_1\);
    
    sum3_cry_4 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[4]\, B => Wt_data(4), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_3\, S => \sum3[4]\, Y
         => OPEN, FCO => \sum3_cry_4\);
    
    sum0_4_axb_29 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[29]\, B => \R1_data[29]\, C => 
        \R0_data[29]\, D => \SIG0[29]_net_1\, Y => 
        \sum0_4_axb_29\);
    
    sum0_4_cry_0_1015 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[0]\, C => 
        \R0_data[12]\, Y => \SIG0_0[10]\);
    
    next_reg_e_cry_17_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[17]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(17), D => \R3_data[17]\, FCI => next_reg_e_cry_16, 
        S => \next_reg_e[17]\, Y => OPEN, FCO => 
        next_reg_e_cry_17);
    
    \next_reg_g[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(18), B => \R5_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[18]_net_1\);
    
    \next_reg_b[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(30), B => \R0_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[30]_net_1\);
    
    sum3_6_0_cry_27 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[27]\, B => \R4_data[27]\, C => 
        \R5_data[27]\, D => \R6_data[27]\, FCI => 
        \sum3_6_0_cry_26\, S => \sum3_6_0[27]\, Y => OPEN, FCO
         => \sum3_6_0_cry_27\);
    
    sum0_4_cry_8 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[8]\, C => 
        \sum0_4_axb_8\, D => GND_net_1, FCI => \sum0_4_cry_7\, S
         => \sum0_4[8]\, Y => OPEN, FCO => \sum0_4_cry_8\);
    
    \SIG0[4]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[17]\, C => 
        \R0_data[6]\, Y => \SIG0[4]_net_1\);
    
    \reg_d[18]\ : SLE
      port map(D => \next_reg_d[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[18]\);
    
    \next_reg_f[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(16), B => \R4_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[16]_net_1\);
    
    sum0_4_cry_3 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[3]\, C => 
        \sum0_4_axb_3\, D => GND_net_1, FCI => \sum0_4_cry_2\, S
         => \sum0_4[3]\, Y => OPEN, FCO => \sum0_4_cry_3\);
    
    \reg_g[5]\ : SLE
      port map(D => \next_reg_g[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[5]\);
    
    sum3_4_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \sum3_6[12]\, B => m157, C => GND_net_1, D
         => GND_net_1, FCI => \sum3_4_cry_11\, S => \sum3_4[12]\, 
        Y => OPEN, FCO => \sum3_4_cry_12\);
    
    \reg_g[24]\ : SLE
      port map(D => \next_reg_g[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[24]\);
    
    next_reg_a_cry_5_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[5]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[5]\, D => N0_data(5), FCI => next_reg_a_cry_4, S
         => \next_reg_a[5]\, Y => OPEN, FCO => next_reg_a_cry_5);
    
    sum3_cry_1 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[1]\, B => Wt_data(1), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_0\, S => \sum3[1]\, Y
         => OPEN, FCO => \sum3_cry_1\);
    
    \next_reg_b[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(23), B => \R0_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[23]_net_1\);
    
    sum3_6_0_cry_1 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[1]\, B => \R4_data[1]\, C => 
        \R5_data[1]\, D => \R6_data[1]\, FCI => \sum3_6_0_cry_0\, 
        S => \sum3_6_0[1]\, Y => OPEN, FCO => \sum3_6_0_cry_1\);
    
    sum3_cry_17 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[17]\, B => Wt_data(17), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_16\, S => 
        \sum3[17]\, Y => OPEN, FCO => \sum3_cry_17\);
    
    \SIG0[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[14]\, C => 
        \R0_data[3]\, Y => \SIG0[1]_net_1\);
    
    \next_reg_d[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(20), B => \R2_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[20]_net_1\);
    
    sum0_4_axb_21 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[21]\, B => \R1_data[21]\, C => 
        \R0_data[21]\, D => \SIG0[21]_net_1\, Y => 
        \sum0_4_axb_21\);
    
    \reg_a[17]\ : SLE
      port map(D => \next_reg_a[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[17]\);
    
    \SIG0[6]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[19]\, C => 
        \R0_data[8]\, Y => \SIG0[6]_net_1\);
    
    \next_reg_f[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(23), B => \R4_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[23]_net_1\);
    
    \reg_b[22]\ : SLE
      port map(D => \next_reg_b[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[22]\);
    
    \next_reg_h[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(28), B => \R6_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[28]_net_1\);
    
    \reg_d[20]\ : SLE
      port map(D => \next_reg_d[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[20]\);
    
    \reg_b[21]\ : SLE
      port map(D => \next_reg_b[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[21]\);
    
    \reg_f[0]\ : SLE
      port map(D => \next_reg_f[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[0]\);
    
    \reg_c[9]\ : SLE
      port map(D => \next_reg_c[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[9]\);
    
    \reg_a[27]\ : SLE
      port map(D => \next_reg_a[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[27]\);
    
    next_reg_a_cry_0_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => sum0_4_cry_0_Y_0, B => oregs_ce_i_a2_0_a2, C
         => sum3_cry_0_Y, D => next_reg_H0_cry_0_0_Y, FCI => 
        GND_net_1, S => OPEN, Y => next_reg_a_cry_0_0_Y, FCO => 
        next_reg_a_cry_0);
    
    \next_reg_c[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(21), B => \R1_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[21]_net_1\);
    
    sum3_cry_21 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[21]\, B => Wt_data(21), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_20\, S => 
        \sum3[21]\, Y => OPEN, FCO => \sum3_cry_21\);
    
    sum0_4_axb_30 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[30]\, B => \R1_data[30]\, C => 
        \R0_data[30]\, D => \SIG0[30]_net_1\, Y => 
        \sum0_4_axb_30\);
    
    \SIG0[8]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[10]\, C => 
        \R0_data[21]\, Y => \SIG0[8]_net_1\);
    
    \reg_g[31]\ : SLE
      port map(D => \next_reg_g[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[31]\);
    
    \reg_d[3]\ : SLE
      port map(D => \next_reg_d[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[3]\);
    
    \SIG0[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[22]\, C => 
        \R0_data[11]\, Y => \SIG0[9]_net_1\);
    
    \reg_e[30]\ : SLE
      port map(D => \next_reg_e[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[30]\);
    
    sum3_6_0_cry_9 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[9]\, B => \R4_data[9]\, C => 
        \R5_data[9]\, D => \R6_data[9]\, FCI => \sum3_6_0_cry_8\, 
        S => \sum3_6_0[9]\, Y => OPEN, FCO => \sum3_6_0_cry_9\);
    
    \reg_e[4]\ : SLE
      port map(D => \next_reg_e[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[4]\);
    
    next_reg_e_cry_22_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[22]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(22), D => \R3_data[22]\, FCI => next_reg_e_cry_21, 
        S => \next_reg_e[22]\, Y => OPEN, FCO => 
        next_reg_e_cry_22);
    
    \next_reg_d[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(22), B => \R2_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[22]_net_1\);
    
    \reg_h[17]\ : SLE
      port map(D => \next_reg_h[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[17]\);
    
    \next_reg_g[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(16), B => \R5_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[16]_net_1\);
    
    sum0_4_cry_24 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[24]\, C => 
        \sum0_4_axb_24\, D => GND_net_1, FCI => \sum0_4_cry_23\, 
        S => \sum0_4[24]\, Y => OPEN, FCO => \sum0_4_cry_24\);
    
    \SIG0[27]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[17]\, C => 
        \R0_data[8]\, Y => \SIG0[27]_net_1\);
    
    sum0_4_axb_22 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[22]\, B => \R1_data[22]\, C => 
        \R0_data[22]\, D => \SIG0[22]_net_1\, Y => 
        \sum0_4_axb_22\);
    
    sum3_cry_5 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[5]\, B => Wt_data(5), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_4\, S => \sum3[5]\, Y
         => OPEN, FCO => \sum3_cry_5\);
    
    \next_reg_c[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(9), B => \R1_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[9]_net_1\);
    
    \reg_f[13]\ : SLE
      port map(D => \next_reg_f[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[13]\);
    
    \reg_c[5]\ : SLE
      port map(D => \next_reg_c[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[5]\);
    
    \reg_b[26]\ : SLE
      port map(D => \next_reg_b[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[26]\);
    
    \reg_h[23]\ : SLE
      port map(D => \next_reg_h[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[23]\);
    
    \next_reg_f[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[1]\, B => N5_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[1]_net_1\);
    
    \reg_d[6]\ : SLE
      port map(D => \next_reg_d[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[6]\);
    
    sum0_4_axb_25 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[25]\, B => \R1_data[25]\, C => 
        \R0_data[25]\, D => \SIG0[25]_net_1\, Y => 
        \sum0_4_axb_25\);
    
    \next_reg_h[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[1]\, B => N7_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[1]_net_1\);
    
    sum0_4_cry_0_1000 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[15]\, C => 
        \R0_data[6]\, Y => \SIG0_0[25]\);
    
    sum3_6_cry_7 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[7]\, B => \R4_data[0]\, C => 
        \R4_data[13]\, D => \R4_data[18]\, FCI => \sum3_6_cry_6\, 
        S => \sum3_6[7]\, Y => OPEN, FCO => \sum3_6_cry_7\);
    
    \next_reg_b[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(28), B => \R0_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[28]_net_1\);
    
    sum3_6_cry_2 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[2]\, B => \R4_data[8]\, C => 
        \R4_data[13]\, D => \R4_data[27]\, FCI => \sum3_6_cry_1\, 
        S => \sum3_6[2]\, Y => OPEN, FCO => \sum3_6_cry_2\);
    
    \next_reg_h[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(26), B => \R6_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[26]_net_1\);
    
    sum3_6_cry_25 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[25]\, B => \R4_data[4]\, C => 
        \R4_data[18]\, D => \R4_data[31]\, FCI => \sum3_6_cry_24\, 
        S => \sum3_6[25]\, Y => OPEN, FCO => \sum3_6_cry_25\);
    
    \reg_d[4]\ : SLE
      port map(D => \next_reg_d[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[4]\);
    
    \reg_e[12]\ : SLE
      port map(D => \next_reg_e[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[12]\);
    
    \next_reg_c[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[6]\, B => N2_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[6]_net_1\);
    
    \reg_b[28]\ : SLE
      port map(D => \next_reg_b[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[28]\);
    
    \reg_e[11]\ : SLE
      port map(D => \next_reg_e[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[11]\);
    
    \next_reg_d[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(8), B => \R2_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[8]_net_1\);
    
    \next_reg_f[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(28), B => \R4_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[28]_net_1\);
    
    \next_reg_c[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(13), B => \R1_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[13]_net_1\);
    
    sum3_6_0_cry_29 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[29]\, B => \R4_data[29]\, C => 
        \R5_data[29]\, D => \R6_data[29]\, FCI => 
        \sum3_6_0_cry_28\, S => \sum3_6_0[29]\, Y => OPEN, FCO
         => \sum3_6_0_cry_29\);
    
    \reg_h[9]\ : SLE
      port map(D => \next_reg_h[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[9]\);
    
    \reg_f[14]\ : SLE
      port map(D => \next_reg_f[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[14]\);
    
    sum3_6_0_cry_15 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[15]\, B => \R4_data[15]\, C => 
        \R5_data[15]\, D => \R6_data[15]\, FCI => 
        \sum3_6_0_cry_14\, S => \sum3_6_0[15]\, Y => OPEN, FCO
         => \sum3_6_0_cry_15\);
    
    sum3_6_cry_17 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[17]\, B => \R4_data[10]\, C => 
        \R4_data[23]\, D => \R4_data[28]\, FCI => \sum3_6_cry_16\, 
        S => \sum3_6[17]\, Y => OPEN, FCO => \sum3_6_cry_17\);
    
    \reg_h[24]\ : SLE
      port map(D => \next_reg_h[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[24]\);
    
    \SIG0[20]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[10]\, B => \R0_data[1]\, C => 
        \R0_data[22]\, Y => \SIG0[20]_net_1\);
    
    \reg_g[29]\ : SLE
      port map(D => \next_reg_g[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[29]\);
    
    \reg_e[23]\ : SLE
      port map(D => \next_reg_e[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[23]\);
    
    sum0_4_cry_0_1016 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[22]\, C => 
        \R0_data[11]\, Y => \SIG0_0[9]\);
    
    \next_reg_g[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[5]\, B => N6_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[5]_net_1\);
    
    \reg_a[30]\ : SLE
      port map(D => \next_reg_a[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[30]\);
    
    \next_reg_f[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(8), B => \R4_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[8]_net_1\);
    
    \reg_b[31]\ : SLE
      port map(D => \next_reg_b[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[31]\);
    
    \next_reg_f[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(7), B => \R4_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[7]_net_1\);
    
    \next_reg_h[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(19), B => \R6_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[19]_net_1\);
    
    \next_reg_g[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[2]\, B => N6_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[2]_net_1\);
    
    \reg_d[31]\ : SLE
      port map(D => \next_reg_d[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[31]\);
    
    \reg_e[16]\ : SLE
      port map(D => \next_reg_e[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[16]\);
    
    \reg_c[7]\ : SLE
      port map(D => \next_reg_c[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[7]\);
    
    next_reg_a_cry_1_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[1]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[1]\, D => N0_data(1), FCI => next_reg_a_cry_0, S
         => \next_reg_a[1]\, Y => OPEN, FCO => next_reg_a_cry_1);
    
    next_reg_e_cry_0_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => sum3_cry_0_Y, B => oregs_ce_i_a2_0_a2, C => 
        next_reg_H4_cry_0_0_Y, D => \R3_data[0]\, FCI => 
        GND_net_1, S => OPEN, Y => next_reg_e_cry_0_0_Y, FCO => 
        next_reg_e_cry_0);
    
    \next_reg_d[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(14), B => \R2_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[14]_net_1\);
    
    \reg_f[5]\ : SLE
      port map(D => \next_reg_f[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[5]\);
    
    sum3_4_s_31 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \sum3_6[31]\, C => m325, D
         => GND_net_1, FCI => \sum3_4_cry_30\, S => \sum3_4[31]\, 
        Y => OPEN, FCO => OPEN);
    
    \next_reg_g[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(7), B => \R5_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[7]_net_1\);
    
    next_reg_e_cry_25_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[25]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(25), D => \R3_data[25]\, FCI => next_reg_e_cry_24, 
        S => \next_reg_e[25]\, Y => OPEN, FCO => 
        next_reg_e_cry_25);
    
    \next_reg_b[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(26), B => \R0_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[26]_net_1\);
    
    sum3_cry_9 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[9]\, B => Wt_data(9), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_8\, S => \sum3[9]\, Y
         => OPEN, FCO => \sum3_cry_9\);
    
    next_reg_e_cry_14_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[14]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(14), D => \R3_data[14]\, FCI => next_reg_e_cry_13, 
        S => \next_reg_e[14]\, Y => OPEN, FCO => 
        next_reg_e_cry_14);
    
    \reg_c[30]\ : SLE
      port map(D => \next_reg_c[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[30]\);
    
    sum0_4_cry_0_1001 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[14]\, C => 
        \R0_data[5]\, Y => \SIG0_0[24]\);
    
    \SIG0[28]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[18]\, C => 
        \R0_data[9]\, Y => \SIG0[28]_net_1\);
    
    \reg_e[24]\ : SLE
      port map(D => \next_reg_e[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[24]\);
    
    \reg_c[15]\ : SLE
      port map(D => \next_reg_c[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[15]\);
    
    \reg_h[31]\ : SLE
      port map(D => \next_reg_h[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[31]\);
    
    \next_reg_b[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(13), B => \R0_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[13]_net_1\);
    
    \reg_g[12]\ : SLE
      port map(D => \next_reg_g[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[12]\);
    
    \reg_e[18]\ : SLE
      port map(D => \next_reg_e[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[18]\);
    
    \reg_c[22]\ : SLE
      port map(D => \next_reg_c[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[22]\);
    
    \next_reg_f[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(26), B => \R4_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[26]_net_1\);
    
    \reg_g[11]\ : SLE
      port map(D => \next_reg_g[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[11]\);
    
    sum0_4_cry_11 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[11]\, C => 
        \sum0_4_axb_11\, D => GND_net_1, FCI => \sum0_4_cry_10\, 
        S => \sum0_4[11]\, Y => OPEN, FCO => \sum0_4_cry_11\);
    
    \reg_d[23]\ : SLE
      port map(D => \next_reg_d[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[23]\);
    
    \next_reg_b[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(31), B => \R0_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[31]_net_1\);
    
    \reg_c[21]\ : SLE
      port map(D => \next_reg_c[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[21]\);
    
    sum0_4_axb_3 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[3]\, B => \R1_data[3]\, C => 
        \R0_data[3]\, D => \SIG0[3]_net_1\, Y => \sum0_4_axb_3\);
    
    next_reg_a_cry_22_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[22]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[22]\, D => N0_data(22), FCI => next_reg_a_cry_21, S
         => \next_reg_a[22]\, Y => OPEN, FCO => next_reg_a_cry_22);
    
    \reg_b[0]\ : SLE
      port map(D => \next_reg_b[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[0]\);
    
    \next_reg_c[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(18), B => \R1_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[18]_net_1\);
    
    \next_reg_g[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(9), B => \R5_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[9]_net_1\);
    
    \reg_f[8]\ : SLE
      port map(D => \next_reg_f[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[8]\);
    
    next_reg_e_cry_19_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[19]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(19), D => \R3_data[19]\, FCI => next_reg_e_cry_18, 
        S => \next_reg_e[19]\, Y => OPEN, FCO => 
        next_reg_e_cry_19);
    
    sum0_4_cry_0_999 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[16]\, C => 
        \R0_data[7]\, Y => \SIG0_0[26]\);
    
    \next_reg_g[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(29), B => \R5_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[29]_net_1\);
    
    next_reg_e_cry_27_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[27]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(27), D => \R3_data[27]\, FCI => next_reg_e_cry_26, 
        S => \next_reg_e[27]\, Y => OPEN, FCO => 
        next_reg_e_cry_27);
    
    \next_reg_d[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(21), B => \R2_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[21]_net_1\);
    
    \SIG0[19]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[21]\, B => \R0_data[9]\, C => 
        \R0_data[0]\, Y => \SIG0[19]_net_1\);
    
    next_reg_e_cry_2_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[2]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(2), D => \R3_data[2]\, FCI => next_reg_e_cry_1, S
         => \next_reg_e[2]\, Y => OPEN, FCO => next_reg_e_cry_2);
    
    sum3_4_cry_8 : ARI1
      generic map(INIT => x"53AC5")

      port map(A => \sum3_6[8]\, B => m110_ns, C => m114, D => 
        Kt_addr(5), FCI => \sum3_4_cry_7\, S => \sum3_4[8]\, Y
         => OPEN, FCO => \sum3_4_cry_8\);
    
    \reg_g[27]\ : SLE
      port map(D => \next_reg_g[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[27]\);
    
    sum3_6_cry_14 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[14]\, B => \R4_data[7]\, C => 
        \R4_data[20]\, D => \R4_data[25]\, FCI => \sum3_6_cry_13\, 
        S => \sum3_6[14]\, Y => OPEN, FCO => \sum3_6_cry_14\);
    
    sum0_4_axb_16 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[16]\, B => \R1_data[16]\, C => 
        \R0_data[16]\, D => \SIG0[16]_net_1\, Y => 
        \sum0_4_axb_16\);
    
    \reg_g[16]\ : SLE
      port map(D => \next_reg_g[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[16]\);
    
    sum0_4_axb_19 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[19]\, B => \R1_data[19]\, C => 
        \R0_data[19]\, D => \SIG0[19]_net_1\, Y => 
        \sum0_4_axb_19\);
    
    \reg_c[26]\ : SLE
      port map(D => \next_reg_c[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[26]\);
    
    \reg_d[24]\ : SLE
      port map(D => \next_reg_d[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[24]\);
    
    sum3_4_cry_17 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[17]\, B => m207_1_0, C => m207_1_1, D
         => Kt_addr(5), FCI => \sum3_4_cry_16\, S => \sum3_4[17]\, 
        Y => OPEN, FCO => \sum3_4_cry_17\);
    
    \next_reg_g[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[3]\, B => N6_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[3]_net_1\);
    
    \reg_f[19]\ : SLE
      port map(D => \next_reg_f[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[19]\);
    
    next_reg_a_cry_12_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[12]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[12]\, D => N0_data(12), FCI => next_reg_a_cry_11, S
         => \next_reg_a[12]\, Y => OPEN, FCO => next_reg_a_cry_12);
    
    \reg_h[29]\ : SLE
      port map(D => \next_reg_h[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[29]\);
    
    \reg_f[22]\ : SLE
      port map(D => \next_reg_f[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[22]\);
    
    next_reg_a_cry_6_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[6]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[6]\, D => N0_data(6), FCI => next_reg_a_cry_5, S
         => \next_reg_a[6]\, Y => OPEN, FCO => next_reg_a_cry_6);
    
    \reg_f[21]\ : SLE
      port map(D => \next_reg_f[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[21]\);
    
    sum3_cry_12 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[12]\, B => Wt_data(12), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_11\, S => 
        \sum3[12]\, Y => OPEN, FCO => \sum3_cry_12\);
    
    \next_reg_c[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(30), B => \R1_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[30]_net_1\);
    
    \reg_g[18]\ : SLE
      port map(D => \next_reg_g[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[18]\);
    
    sum0_4_axb_8 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[8]\, B => \R1_data[8]\, C => 
        \R0_data[8]\, D => \SIG0[8]_net_1\, Y => \sum0_4_axb_8\);
    
    \reg_c[28]\ : SLE
      port map(D => \next_reg_c[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[28]\);
    
    sum3_6_0_cry_4 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[4]\, B => \R4_data[4]\, C => 
        \R5_data[4]\, D => \R6_data[4]\, FCI => \sum3_6_0_cry_3\, 
        S => \sum3_6_0[4]\, Y => OPEN, FCO => \sum3_6_0_cry_4\);
    
    \next_reg_b[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(18), B => \R0_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[18]_net_1\);
    
    next_reg_a_cry_8_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[8]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[8]\, D => N0_data(8), FCI => next_reg_a_cry_7, S
         => \next_reg_a[8]\, Y => OPEN, FCO => next_reg_a_cry_8);
    
    sum3_6_0_cry_18 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[18]\, B => \R4_data[18]\, C => 
        \R5_data[18]\, D => \R6_data[18]\, FCI => 
        \sum3_6_0_cry_17\, S => \sum3_6_0[18]\, Y => OPEN, FCO
         => \sum3_6_0_cry_18\);
    
    \next_reg_c[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(16), B => \R1_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[16]_net_1\);
    
    \next_reg_d[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(17), B => \R2_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[17]_net_1\);
    
    sum0_4_axb_11 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[11]\, B => \R1_data[11]\, C => 
        \R0_data[11]\, D => \SIG0[11]_net_1\, Y => 
        \sum0_4_axb_11\);
    
    sum0_4_cry_2 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[2]\, C => 
        \sum0_4_axb_2\, D => GND_net_1, FCI => \sum0_4_cry_1\, S
         => \sum0_4[2]\, Y => OPEN, FCO => \sum0_4_cry_2\);
    
    sum0_4_cry_25 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[25]\, C => 
        \sum0_4_axb_25\, D => GND_net_1, FCI => \sum0_4_cry_24\, 
        S => \sum0_4[25]\, Y => OPEN, FCO => \sum0_4_cry_25\);
    
    \next_reg_d[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(15), B => \R2_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[15]_net_1\);
    
    \reg_c[10]\ : SLE
      port map(D => \next_reg_c[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[10]\);
    
    \next_reg_c[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(23), B => \R1_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[23]_net_1\);
    
    \reg_d[15]\ : SLE
      port map(D => \next_reg_d[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[15]\);
    
    \reg_a[5]\ : SLE
      port map(D => \next_reg_a[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[5]\);
    
    \reg_b[1]\ : SLE
      port map(D => \next_reg_b[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[1]\);
    
    \reg_b[12]\ : SLE
      port map(D => \next_reg_b[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[12]\);
    
    \SIG0[2]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[24]\, B => \R0_data[15]\, C => 
        \R0_data[4]\, Y => \SIG0[2]_net_1\);
    
    sum0_4_axb_23 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[23]\, B => \R1_data[23]\, C => 
        \R0_data[23]\, D => \SIG0[23]_net_1\, Y => 
        \sum0_4_axb_23\);
    
    \next_reg_d[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(30), B => \R2_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[30]_net_1\);
    
    sum0_4_axb_5 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[5]\, B => \R1_data[5]\, C => 
        \R0_data[5]\, D => \SIG0[5]_net_1\, Y => \sum0_4_axb_5\);
    
    \reg_b[11]\ : SLE
      port map(D => \next_reg_b[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[11]\);
    
    sum0_4_cry_0_1023 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[24]\, B => \R0_data[15]\, C => 
        \R0_data[4]\, Y => \SIG0_0[2]\);
    
    \reg_f[26]\ : SLE
      port map(D => \next_reg_f[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[26]\);
    
    next_reg_e_cry_10_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[10]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(10), D => \R3_data[10]\, FCI => next_reg_e_cry_9, 
        S => \next_reg_e[10]\, Y => OPEN, FCO => 
        next_reg_e_cry_10);
    
    \reg_e[29]\ : SLE
      port map(D => \next_reg_e[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[29]\);
    
    \next_reg_b[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[2]\, B => N1_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[2]_net_1\);
    
    sum3_cry_8 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[8]\, B => Wt_data(8), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_7\, S => \sum3[8]\, Y
         => OPEN, FCO => \sum3_cry_8\);
    
    sum3_cry_23 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[23]\, B => Wt_data(23), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_22\, S => 
        \sum3[23]\, Y => OPEN, FCO => \sum3_cry_23\);
    
    sum0_4_cry_0_1013 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[14]\, C => 
        \R0_data[2]\, Y => \SIG0_0[12]\);
    
    sum0_4_axb_20 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[20]\, B => \R1_data[20]\, C => 
        \R0_data[20]\, D => \SIG0[20]_net_1\, Y => 
        \sum0_4_axb_20\);
    
    next_reg_a_cry_25_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[25]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[25]\, D => N0_data(25), FCI => next_reg_a_cry_24, S
         => \next_reg_a[25]\, Y => OPEN, FCO => next_reg_a_cry_25);
    
    \next_reg_f[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(19), B => \R4_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[19]_net_1\);
    
    sum3_4_cry_21 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[21]\, B => m235_ns, C => m239, D => 
        Kt_addr(5), FCI => \sum3_4_cry_20\, S => \sum3_4[21]\, Y
         => OPEN, FCO => \sum3_4_cry_21\);
    
    \Maj[31]\ : CFG3
      generic map(INIT => x"E8")

      port map(A => \R2_data[31]\, B => \R1_data[31]\, C => 
        \R0_data[31]\, Y => \Maj[31]_net_1\);
    
    \SIG0[13]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[15]\, C => 
        \R0_data[3]\, Y => \SIG0[13]_net_1\);
    
    sum0_4_axb_12 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[12]\, B => \R1_data[12]\, C => 
        \R0_data[12]\, D => \SIG0[12]_net_1\, Y => 
        \sum0_4_axb_12\);
    
    sum3_cry_6 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[6]\, B => Wt_data(6), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_5\, S => \sum3[6]\, Y
         => OPEN, FCO => \sum3_cry_6\);
    
    \reg_f[28]\ : SLE
      port map(D => \next_reg_f[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[28]\);
    
    sum0_4_cry_0_1018 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[20]\, C => 
        \R0_data[9]\, Y => \SIG0_0[7]\);
    
    \reg_f[17]\ : SLE
      port map(D => \next_reg_f[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[17]\);
    
    sum3_4_cry_14 : ARI1
      generic map(INIT => x"5C53A")

      port map(A => \sum3_6[14]\, B => m172_ns, C => m177, D => 
        Kt_addr(5), FCI => \sum3_4_cry_13\, S => \sum3_4[14]\, Y
         => OPEN, FCO => \sum3_4_cry_14\);
    
    \reg_h[27]\ : SLE
      port map(D => \next_reg_h[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[27]\);
    
    \reg_b[16]\ : SLE
      port map(D => \next_reg_b[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[16]\);
    
    sum0_4_axb_15 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[15]\, B => \R1_data[15]\, C => 
        \R0_data[15]\, D => \SIG0[15]_net_1\, Y => 
        \sum0_4_axb_15\);
    
    \next_reg_b[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(16), B => \R0_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[16]_net_1\);
    
    \next_reg_h[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(14), B => \R6_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[14]_net_1\);
    
    sum0_4_axb_9 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[9]\, B => \R1_data[9]\, C => 
        \R0_data[9]\, D => \SIG0[9]_net_1\, Y => \sum0_4_axb_9\);
    
    sum0_4_cry_0_1022 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[16]\, C => 
        \R0_data[5]\, Y => \SIG0_0[3]\);
    
    next_reg_a_cry_27_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[27]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[27]\, D => N0_data(27), FCI => next_reg_a_cry_26, S
         => \next_reg_a[27]\, Y => OPEN, FCO => next_reg_a_cry_27);
    
    next_reg_a_cry_15_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[15]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[15]\, D => N0_data(15), FCI => next_reg_a_cry_14, S
         => \next_reg_a[15]\, Y => OPEN, FCO => next_reg_a_cry_15);
    
    \reg_d[29]\ : SLE
      port map(D => \next_reg_d[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[29]\);
    
    sum0_4_cry_5 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[5]\, C => 
        \sum0_4_axb_5\, D => GND_net_1, FCI => \sum0_4_cry_4\, S
         => \sum0_4[5]\, Y => OPEN, FCO => \sum0_4_cry_5\);
    
    next_reg_e_cry_1_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[1]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(1), D => \R3_data[1]\, FCI => next_reg_e_cry_0, S
         => \next_reg_e[1]\, Y => OPEN, FCO => next_reg_e_cry_1);
    
    sum0_4_cry_0_1012 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[15]\, C => 
        \R0_data[3]\, Y => \SIG0_0[13]\);
    
    \reg_b[9]\ : SLE
      port map(D => \next_reg_b[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[9]\);
    
    \next_reg_c[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(28), B => \R1_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[28]_net_1\);
    
    \reg_b[18]\ : SLE
      port map(D => \next_reg_b[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[18]\);
    
    \next_reg_g[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(19), B => \R5_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[19]_net_1\);
    
    sum0_4_cry_10 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[10]\, C => 
        \sum0_4_axb_10\, D => GND_net_1, FCI => \sum0_4_cry_9\, S
         => \sum0_4[10]\, Y => OPEN, FCO => \sum0_4_cry_10\);
    
    sum3_6_0_cry_8 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[8]\, B => \R4_data[8]\, C => 
        \R5_data[8]\, D => \R6_data[8]\, FCI => \sum3_6_0_cry_7\, 
        S => \sum3_6_0[8]\, Y => OPEN, FCO => \sum3_6_0_cry_8\);
    
    \next_reg_c[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[0]\, B => next_reg_H2_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_c[0]_net_1\);
    
    \reg_d[7]\ : SLE
      port map(D => \next_reg_d[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[7]\);
    
    sum3_6_cry_0_992 : CFG4
      generic map(INIT => x"5A66")

      port map(A => \R7_data[0]\, B => \R6_data[0]\, C => 
        \R5_data[0]\, D => \R4_data[0]\, Y => sum3_6_0);
    
    \next_reg_d[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(10), B => \R2_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[10]_net_1\);
    
    \reg_d[10]\ : SLE
      port map(D => \next_reg_d[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[10]\);
    
    \SIG0[21]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[11]\, C => 
        \R0_data[2]\, Y => \SIG0[21]_net_1\);
    
    next_reg_e_cry_6_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[6]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(6), D => \R3_data[6]\, FCI => next_reg_e_cry_5, S
         => \next_reg_e[6]\, Y => OPEN, FCO => next_reg_e_cry_6);
    
    sum3_4_cry_9 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[9]\, B => m119_ns, C => m124, D => 
        Kt_addr(5), FCI => \sum3_4_cry_8\, S => \sum3_4[9]\, Y
         => OPEN, FCO => \sum3_4_cry_9\);
    
    \reg_e[27]\ : SLE
      port map(D => \next_reg_e[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[27]\);
    
    \reg_b[25]\ : SLE
      port map(D => \next_reg_b[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[25]\);
    
    \reg_g[3]\ : SLE
      port map(D => \next_reg_g[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[3]\);
    
    \next_reg_c[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[3]\, B => N2_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[3]_net_1\);
    
    next_reg_a_cry_17_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[17]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[17]\, D => N0_data(17), FCI => next_reg_a_cry_16, S
         => \next_reg_a[17]\, Y => OPEN, FCO => next_reg_a_cry_17);
    
    next_reg_e_cry_24_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[24]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(24), D => \R3_data[24]\, FCI => next_reg_e_cry_23, 
        S => \next_reg_e[24]\, Y => OPEN, FCO => 
        next_reg_e_cry_24);
    
    \next_reg_g[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(24), B => \R5_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[24]_net_1\);
    
    sum0_4_axb_0 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[0]\, B => \R1_data[0]\, C => 
        \R0_data[0]\, D => sum0_4, Y => \sum0_4[0]\);
    
    \next_reg_h[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(29), B => \R6_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[29]_net_1\);
    
    \reg_h[3]\ : SLE
      port map(D => \next_reg_h[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[3]\);
    
    next_reg_e_cry_13_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[13]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(13), D => \R3_data[13]\, FCI => next_reg_e_cry_12, 
        S => \next_reg_e[13]\, Y => OPEN, FCO => 
        next_reg_e_cry_13);
    
    sum0_4_cry_13 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[13]\, C => 
        \sum0_4_axb_13\, D => GND_net_1, FCI => \sum0_4_cry_12\, 
        S => \sum0_4[13]\, Y => OPEN, FCO => \sum0_4_cry_13\);
    
    sum0_4_axb_4 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[4]\, B => \R1_data[4]\, C => 
        \R0_data[4]\, D => \SIG0[4]_net_1\, Y => \sum0_4_axb_4\);
    
    sum0_4_cry_0_995 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[20]\, B => \R0_data[11]\, C => 
        \R0_data[0]\, Y => \SIG0_0[30]\);
    
    \reg_g[2]\ : SLE
      port map(D => \next_reg_g[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[2]\);
    
    \next_reg_d[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(12), B => \R2_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[12]_net_1\);
    
    sum3_s_31 : ARI1
      generic map(INIT => x"46600")

      port map(A => VCC_net_1, B => \sum3_4[31]\, C => 
        Wt_data(31), D => GND_net_1, FCI => \sum3_cry_30\, S => 
        \sum3[31]\, Y => OPEN, FCO => OPEN);
    
    sum3_6_0_cry_23 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[23]\, B => \R4_data[23]\, C => 
        \R5_data[23]\, D => \R6_data[23]\, FCI => 
        \sum3_6_0_cry_22\, S => \sum3_6_0[23]\, Y => OPEN, FCO
         => \sum3_6_0_cry_23\);
    
    sum3_6_cry_3 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[3]\, B => \R4_data[9]\, C => 
        \R4_data[14]\, D => \R4_data[28]\, FCI => \sum3_6_cry_2\, 
        S => \sum3_6[3]\, Y => OPEN, FCO => \sum3_6_cry_3\);
    
    sum3_6_0_cry_12 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[12]\, B => \R4_data[12]\, C => 
        \R5_data[12]\, D => \R6_data[12]\, FCI => 
        \sum3_6_0_cry_11\, S => \sum3_6_0[12]\, Y => OPEN, FCO
         => \sum3_6_0_cry_12\);
    
    \next_reg_f[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[2]\, B => N5_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[2]_net_1\);
    
    \SIG0[17]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[19]\, C => 
        \R0_data[7]\, Y => \SIG0[17]_net_1\);
    
    \reg_h[1]\ : SLE
      port map(D => \next_reg_h[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[1]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    sum3_6_cry_1 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[1]\, B => \R4_data[7]\, C => 
        \R4_data[12]\, D => \R4_data[26]\, FCI => \sum3_6_cry_0\, 
        S => \sum3_6[1]\, Y => OPEN, FCO => \sum3_6_cry_1\);
    
    \next_reg_d[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[5]\, B => N3_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[5]_net_1\);
    
    sum3_6_cry_15 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[15]\, B => \R4_data[8]\, C => 
        \R4_data[21]\, D => \R4_data[26]\, FCI => \sum3_6_cry_14\, 
        S => \sum3_6[15]\, Y => OPEN, FCO => \sum3_6_cry_15\);
    
    sum0_4_cry_18 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[18]\, C => 
        \sum0_4_axb_18\, D => GND_net_1, FCI => \sum0_4_cry_17\, 
        S => \sum0_4[18]\, Y => OPEN, FCO => \sum0_4_cry_18\);
    
    \reg_c[13]\ : SLE
      port map(D => \next_reg_c[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[13]\);
    
    \next_reg_c[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(26), B => \R1_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[26]_net_1\);
    
    next_reg_e_cry_29_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[29]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(29), D => \R3_data[29]\, FCI => next_reg_e_cry_28, 
        S => \next_reg_e[29]\, Y => OPEN, FCO => 
        next_reg_e_cry_29);
    
    \next_reg_h[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[2]\, B => N7_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[2]_net_1\);
    
    \next_reg_b[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(8), B => \R0_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[8]_net_1\);
    
    sum3_6_cry_21 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[21]\, B => \R4_data[0]\, C => 
        \R4_data[14]\, D => \R4_data[27]\, FCI => \sum3_6_cry_20\, 
        S => \sum3_6[21]\, Y => OPEN, FCO => \sum3_6_cry_21\);
    
    sum0_4_axb_2 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[2]\, B => \R1_data[2]\, C => 
        \R0_data[2]\, D => \SIG0[2]_net_1\, Y => \sum0_4_axb_2\);
    
    \reg_d[27]\ : SLE
      port map(D => \next_reg_d[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[27]\);
    
    sum0_4_axb_7 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[7]\, B => \R1_data[7]\, C => 
        \R0_data[7]\, D => \SIG0[7]_net_1\, Y => \sum0_4_axb_7\);
    
    \next_reg_d[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(23), B => \R2_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[23]_net_1\);
    
    \next_reg_c[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(31), B => \R1_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[31]_net_1\);
    
    \reg_a[12]\ : SLE
      port map(D => \next_reg_a[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[12]\);
    
    \next_reg_h[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(17), B => \R6_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[17]_net_1\);
    
    sum0_4_cry_0_997 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[18]\, C => 
        \R0_data[9]\, Y => \SIG0_0[28]\);
    
    sum0_4_cry_0_1024 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[14]\, C => 
        \R0_data[3]\, Y => \SIG0_0[1]\);
    
    \reg_a[11]\ : SLE
      port map(D => \next_reg_a[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[11]\);
    
    \next_reg_h[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[4]\, B => N7_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[4]_net_1\);
    
    \next_reg_h[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(15), B => \R6_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[15]_net_1\);
    
    sum0_4_cry_0_1014 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[13]\, B => \R0_data[1]\, C => 
        \R0_data[24]\, Y => \SIG0_0[11]\);
    
    sum3_6_cry_0 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => sum3_6_0, C => \sum3_6[0]\, D
         => GND_net_1, FCI => GND_net_1, S => OPEN, Y => 
        sum3_6_cry_0_Y, FCO => \sum3_6_cry_0\);
    
    \reg_e[15]\ : SLE
      port map(D => \next_reg_e[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[15]\);
    
    \reg_a[22]\ : SLE
      port map(D => \next_reg_a[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[22]\);
    
    \next_reg_b[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[4]\, B => N1_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[4]_net_1\);
    
    sum0_4_axb_24 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[24]\, B => \R1_data[24]\, C => 
        \R0_data[24]\, D => \SIG0[24]_net_1\, Y => 
        \sum0_4_axb_24\);
    
    \reg_a[21]\ : SLE
      port map(D => \next_reg_a[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[21]\);
    
    sum3_cry_20 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[20]\, B => Wt_data(20), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_19\, S => 
        \sum3[20]\, Y => OPEN, FCO => \sum3_cry_20\);
    
    sum3_cry_11 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[11]\, B => Wt_data(11), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_10\, S => 
        \sum3[11]\, Y => OPEN, FCO => \sum3_cry_11\);
    
    \next_reg_b[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(29), B => \R0_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[29]_net_1\);
    
    \next_reg_f[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[4]\, B => N5_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[4]_net_1\);
    
    \reg_e[7]\ : SLE
      port map(D => \next_reg_e[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[7]\);
    
    sum3_6_0_cry_17 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[17]\, B => \R4_data[17]\, C => 
        \R5_data[17]\, D => \R6_data[17]\, FCI => 
        \sum3_6_0_cry_16\, S => \sum3_6_0[17]\, Y => OPEN, FCO
         => \sum3_6_0_cry_17\);
    
    \reg_c[14]\ : SLE
      port map(D => \next_reg_c[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[14]\);
    
    \SIG0[10]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[0]\, C => 
        \R0_data[12]\, Y => \SIG0[10]_net_1\);
    
    next_reg_a_s_31 : ARI1
      generic map(INIT => x"47D28")

      port map(A => N0_data(31), B => oregs_ce_i_a2_0_a2, C => 
        \sum0_4[31]\, D => \sum3[31]\, FCI => next_reg_a_cry_30, 
        S => \next_reg_a[31]\, Y => OPEN, FCO => OPEN);
    
    \next_reg_d[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(31), B => \R2_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[31]_net_1\);
    
    \reg_b[20]\ : SLE
      port map(D => \next_reg_b[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[20]\);
    
    sum3_4_cry_20 : ARI1
      generic map(INIT => x"5C53A")

      port map(A => \sum3_6[20]\, B => m226_ns, C => m230, D => 
        Kt_addr(5), FCI => \sum3_4_cry_19\, S => \sum3_4[20]\, Y
         => OPEN, FCO => \sum3_4_cry_20\);
    
    \SIG0[24]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[14]\, C => 
        \R0_data[5]\, Y => \SIG0[24]_net_1\);
    
    \next_reg_f[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(29), B => \R4_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[29]_net_1\);
    
    \reg_h[12]\ : SLE
      port map(D => \next_reg_h[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[12]\);
    
    \next_reg_f[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(14), B => \R4_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[14]_net_1\);
    
    next_reg_e_cry_7_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[7]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(7), D => \R3_data[7]\, FCI => next_reg_e_cry_6, S
         => \next_reg_e[7]\, Y => OPEN, FCO => next_reg_e_cry_7);
    
    next_reg_a_cry_3_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[3]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[3]\, D => N0_data(3), FCI => next_reg_a_cry_2, S
         => \next_reg_a[3]\, Y => OPEN, FCO => next_reg_a_cry_3);
    
    \reg_h[11]\ : SLE
      port map(D => \next_reg_h[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[11]\);
    
    sum0_4_axb_27 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[27]\, B => \R1_data[27]\, C => 
        \R0_data[27]\, D => \SIG0[27]_net_1\, Y => 
        \sum0_4_axb_27\);
    
    \reg_a[16]\ : SLE
      port map(D => \next_reg_a[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[16]\);
    
    \reg_a[3]\ : SLE
      port map(D => \next_reg_a[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[3]\);
    
    \next_reg_d[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(9), B => \R2_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[9]_net_1\);
    
    \reg_g[30]\ : SLE
      port map(D => \next_reg_g[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[30]\);
    
    \reg_g[4]\ : SLE
      port map(D => \next_reg_g[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[4]\);
    
    sum3_4_cry_7 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[7]\, B => m104_am, C => m104_bm, D
         => Kt_addr_5_rep1, FCI => \sum3_4_cry_6\, S => 
        \sum3_4[7]\, Y => OPEN, FCO => \sum3_4_cry_7\);
    
    \next_reg_d[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[3]\, B => N3_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[3]_net_1\);
    
    \reg_a[26]\ : SLE
      port map(D => \next_reg_a[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[26]\);
    
    \next_reg_g[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(27), B => \R5_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[27]_net_1\);
    
    \next_reg_g[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(25), B => \R5_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[25]_net_1\);
    
    next_reg_e_cry_20_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[20]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(20), D => \R3_data[20]\, FCI => next_reg_e_cry_19, 
        S => \next_reg_e[20]\, Y => OPEN, FCO => 
        next_reg_e_cry_20);
    
    sum0_4_cry_0_1005 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[10]\, B => \R0_data[1]\, C => 
        \R0_data[22]\, Y => \SIG0_0[20]\);
    
    sum0_4_cry_30 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[30]\, C => 
        \sum0_4_axb_30\, D => GND_net_1, FCI => \sum0_4_cry_29\, 
        S => \sum0_4[30]\, Y => OPEN, FCO => \sum0_4_cry_30\);
    
    \next_reg_c[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[1]\, B => N2_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[1]_net_1\);
    
    sum3_4_cry_23 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[23]\, B => m254, C => m258_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_22\, S => \sum3_4[23]\, Y
         => OPEN, FCO => \sum3_4_cry_23\);
    
    sum0_4_cry_0_1019 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[19]\, C => 
        \R0_data[8]\, Y => \SIG0_0[6]\);
    
    \reg_a[7]\ : SLE
      port map(D => \next_reg_a[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[7]\);
    
    \SIG0[18]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[20]\, C => 
        \R0_data[8]\, Y => \SIG0[18]_net_1\);
    
    \reg_a[18]\ : SLE
      port map(D => \next_reg_a[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[18]\);
    
    \reg_e[6]\ : SLE
      port map(D => \next_reg_e[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[6]\);
    
    \next_reg_d[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(28), B => \R2_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[28]_net_1\);
    
    \reg_d[13]\ : SLE
      port map(D => \next_reg_d[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[13]\);
    
    next_reg_a_cry_24_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[24]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[24]\, D => N0_data(24), FCI => next_reg_a_cry_23, S
         => \next_reg_a[24]\, Y => OPEN, FCO => next_reg_a_cry_24);
    
    \reg_h[16]\ : SLE
      port map(D => \next_reg_h[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[16]\);
    
    sum3_4_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \sum3_6[1]\, B => m34, C => GND_net_1, D => 
        GND_net_1, FCI => \sum3_4_cry_0\, S => \sum3_4[1]\, Y => 
        OPEN, FCO => \sum3_4_cry_1\);
    
    sum0_4_axb_13 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[13]\, B => \R1_data[13]\, C => 
        \R0_data[13]\, D => \SIG0[13]_net_1\, Y => 
        \sum0_4_axb_13\);
    
    \reg_c[6]\ : SLE
      port map(D => \next_reg_c[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[6]\);
    
    sum3_4_cry_15 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_6[15]\, B => Kt_data_15, C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_4_cry_14\, S => \sum3_4[15]\, 
        Y => OPEN, FCO => \sum3_4_cry_15\);
    
    sum3_4_cry_0 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \Kt_data_0[0]\, C => 
        \sum3_4[0]\, D => GND_net_1, FCI => GND_net_1, S => OPEN, 
        Y => sum3_4_cry_0_Y, FCO => \sum3_4_cry_0\);
    
    \next_reg_f[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[3]\, B => N5_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[3]_net_1\);
    
    \reg_g[15]\ : SLE
      port map(D => \next_reg_g[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[15]\);
    
    sum0_4_cry_19 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[19]\, C => 
        \sum0_4_axb_19\, D => GND_net_1, FCI => \sum0_4_cry_18\, 
        S => \sum0_4[19]\, Y => OPEN, FCO => \sum0_4_cry_19\);
    
    \reg_a[28]\ : SLE
      port map(D => \next_reg_a[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[28]\);
    
    \reg_c[25]\ : SLE
      port map(D => \next_reg_c[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[25]\);
    
    sum0_4_axb_10 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[10]\, B => \R1_data[10]\, C => 
        \R0_data[10]\, D => \SIG0[10]_net_1\, Y => 
        \sum0_4_axb_10\);
    
    \reg_c[3]\ : SLE
      port map(D => \next_reg_c[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[3]\);
    
    sum3_4_cry_28 : ARI1
      generic map(INIT => x"53AC5")

      port map(A => \sum3_6[28]\, B => m296, C => m300_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_27\, S => \sum3_4[28]\, Y
         => OPEN, FCO => \sum3_4_cry_28\);
    
    sum3_6_0_cry_0 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[0]\, B => \R4_data[0]\, C => 
        \R5_data[0]\, D => \R6_data[0]\, FCI => GND_net_1, S => 
        OPEN, Y => sum3_6_0_cry_0_Y, FCO => \sum3_6_0_cry_0\);
    
    \next_reg_g[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(14), B => \R5_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[14]_net_1\);
    
    \SIG0[25]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[15]\, C => 
        \R0_data[6]\, Y => \SIG0[25]_net_1\);
    
    \next_reg_h[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[3]\, B => N7_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[3]_net_1\);
    
    \next_reg_b[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[6]\, B => N1_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[6]_net_1\);
    
    sum0_4_cry_16 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[16]\, C => 
        \sum0_4_axb_16\, D => GND_net_1, FCI => \sum0_4_cry_15\, 
        S => \sum0_4[16]\, Y => OPEN, FCO => \sum0_4_cry_16\);
    
    \next_reg_h[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(10), B => \R6_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[10]_net_1\);
    
    sum3_cry_29 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[29]\, B => Wt_data(29), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_28\, S => 
        \sum3[29]\, Y => OPEN, FCO => \sum3_cry_29\);
    
    \reg_e[10]\ : SLE
      port map(D => \next_reg_e[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[10]\);
    
    next_reg_e_s_31 : ARI1
      generic map(INIT => x"472D8")

      port map(A => \R3_data[31]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[31]\, D => N4_data(31), FCI => next_reg_e_cry_30, S
         => \next_reg_e[31]\, Y => OPEN, FCO => OPEN);
    
    sum3_cry_28 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[28]\, B => Wt_data(28), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_27\, S => 
        \sum3[28]\, Y => OPEN, FCO => \sum3_cry_28\);
    
    \reg_h[18]\ : SLE
      port map(D => \next_reg_h[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[18]\);
    
    next_reg_a_cry_29_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[29]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[29]\, D => N0_data(29), FCI => next_reg_a_cry_28, S
         => \next_reg_a[29]\, Y => OPEN, FCO => next_reg_a_cry_29);
    
    sum3_6_s_31 : ARI1
      generic map(INIT => x"46996")

      port map(A => \R4_data[24]\, B => \sum3_6_0[31]\, C => 
        \R4_data[5]\, D => \R4_data[10]\, FCI => \sum3_6_cry_30\, 
        S => \sum3_6[31]\, Y => OPEN, FCO => OPEN);
    
    \next_reg_d[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(11), B => \R2_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[11]_net_1\);
    
    \next_reg_c[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(19), B => \R1_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[19]_net_1\);
    
    \reg_c[1]\ : SLE
      port map(D => \next_reg_c[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[1]\);
    
    \next_reg_h[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(7), B => \R6_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[7]_net_1\);
    
    \reg_h[6]\ : SLE
      port map(D => \next_reg_h[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[6]\);
    
    \reg_d[14]\ : SLE
      port map(D => \next_reg_d[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[14]\);
    
    next_reg_a_cry_14_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[14]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[14]\, D => N0_data(14), FCI => next_reg_a_cry_13, S
         => \next_reg_a[14]\, Y => OPEN, FCO => next_reg_a_cry_14);
    
    next_reg_a_cry_2_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[2]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[2]\, D => N0_data(2), FCI => next_reg_a_cry_1, S
         => \next_reg_a[2]\, Y => OPEN, FCO => next_reg_a_cry_2);
    
    \reg_g[0]\ : SLE
      port map(D => \next_reg_g[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[0]\);
    
    \next_reg_h[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(24), B => \R6_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[24]_net_1\);
    
    \reg_h[2]\ : SLE
      port map(D => \next_reg_h[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[2]\);
    
    \reg_b[30]\ : SLE
      port map(D => \next_reg_b[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[30]\);
    
    \reg_c[19]\ : SLE
      port map(D => \next_reg_c[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[19]\);
    
    \next_reg_h[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(12), B => \R6_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[12]_net_1\);
    
    sum3_6_cry_9 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[9]\, B => \R4_data[2]\, C => 
        \R4_data[15]\, D => \R4_data[20]\, FCI => \sum3_6_cry_8\, 
        S => \sum3_6[9]\, Y => OPEN, FCO => \sum3_6_cry_9\);
    
    \next_reg_d[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(26), B => \R2_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[26]_net_1\);
    
    \reg_d[30]\ : SLE
      port map(D => \next_reg_d[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[30]\);
    
    sum3_6_0_cry_19 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[19]\, B => \R4_data[19]\, C => 
        \R5_data[19]\, D => \R6_data[19]\, FCI => 
        \sum3_6_0_cry_18\, S => \sum3_6_0[19]\, Y => OPEN, FCO
         => \sum3_6_0_cry_19\);
    
    \reg_f[25]\ : SLE
      port map(D => \next_reg_f[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[25]\);
    
    \next_reg_f[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(17), B => \R4_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[17]_net_1\);
    
    \next_reg_h[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[0]\, B => next_reg_H7_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_h[0]_net_1\);
    
    \next_reg_f[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(15), B => \R4_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[15]_net_1\);
    
    sum0_4_cry_21 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[21]\, C => 
        \sum0_4_axb_21\, D => GND_net_1, FCI => \sum0_4_cry_20\, 
        S => \sum0_4[21]\, Y => OPEN, FCO => \sum0_4_cry_21\);
    
    sum0_4_cry_12 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[12]\, C => 
        \sum0_4_axb_12\, D => GND_net_1, FCI => \sum0_4_cry_11\, 
        S => \sum0_4[12]\, Y => OPEN, FCO => \sum0_4_cry_12\);
    
    sum3_6_0_cry_20 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[20]\, B => \R4_data[20]\, C => 
        \R5_data[20]\, D => \R6_data[20]\, FCI => 
        \sum3_6_0_cry_19\, S => \sum3_6_0[20]\, Y => OPEN, FCO
         => \sum3_6_0_cry_20\);
    
    sum3_cry_0 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \Wt_data_0[0]\, C => 
        \sum3[0]\, D => GND_net_1, FCI => GND_net_1, S => OPEN, Y
         => sum3_cry_0_Y, FCO => \sum3_cry_0\);
    
    sum3_6_0_cry_26 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[26]\, B => \R4_data[26]\, C => 
        \R5_data[26]\, D => \R6_data[26]\, FCI => 
        \sum3_6_0_cry_25\, S => \sum3_6_0[26]\, Y => OPEN, FCO
         => \sum3_6_0_cry_26\);
    
    sum0_4_cry_9 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[9]\, C => 
        \sum0_4_axb_9\, D => GND_net_1, FCI => \sum0_4_cry_8\, S
         => \sum0_4[9]\, Y => OPEN, FCO => \sum0_4_cry_9\);
    
    next_reg_a_cry_19_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[19]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[19]\, D => N0_data(19), FCI => next_reg_a_cry_18, S
         => \next_reg_a[19]\, Y => OPEN, FCO => next_reg_a_cry_19);
    
    \reg_g[8]\ : SLE
      port map(D => \next_reg_g[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[8]\);
    
    \reg_d[1]\ : SLE
      port map(D => \next_reg_d[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[1]\);
    
    sum3_6_cry_20 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[20]\, B => \R4_data[13]\, C => 
        \R4_data[26]\, D => \R4_data[31]\, FCI => \sum3_6_cry_19\, 
        S => \sum3_6[20]\, Y => OPEN, FCO => \sum3_6_cry_20\);
    
    \next_reg_g[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(20), B => \R5_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[20]_net_1\);
    
    \next_reg_g[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(30), B => \R5_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[30]_net_1\);
    
    \reg_b[8]\ : SLE
      port map(D => \next_reg_b[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[8]\);
    
    next_reg_e_cry_23_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[23]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(23), D => \R3_data[23]\, FCI => next_reg_e_cry_22, 
        S => \next_reg_e[23]\, Y => OPEN, FCO => 
        next_reg_e_cry_23);
    
    \reg_h[30]\ : SLE
      port map(D => \next_reg_h[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[30]\);
    
    \next_reg_d[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[6]\, B => N3_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[6]_net_1\);
    
    \reg_g[10]\ : SLE
      port map(D => \next_reg_g[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[10]\);
    
    \reg_e[2]\ : SLE
      port map(D => \next_reg_e[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[2]\);
    
    \reg_c[20]\ : SLE
      port map(D => \next_reg_c[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[20]\);
    
    \next_reg_b[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(19), B => \R0_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[19]_net_1\);
    
    sum0_4_cry_0_1017 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[10]\, C => 
        \R0_data[21]\, Y => \SIG0_0[8]\);
    
    \reg_b[23]\ : SLE
      port map(D => \next_reg_b[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[23]\);
    
    \next_reg_f[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(30), B => \R4_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[30]_net_1\);
    
    \reg_g[22]\ : SLE
      port map(D => \next_reg_g[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[22]\);
    
    \reg_c[8]\ : SLE
      port map(D => \next_reg_c[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[8]\);
    
    \reg_b[15]\ : SLE
      port map(D => \next_reg_b[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[15]\);
    
    \reg_g[21]\ : SLE
      port map(D => \next_reg_g[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[21]\);
    
    \reg_h[7]\ : SLE
      port map(D => \next_reg_h[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[7]\);
    
    next_reg_a_cry_20_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[20]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[20]\, D => N0_data(20), FCI => next_reg_a_cry_19, S
         => \next_reg_a[20]\, Y => OPEN, FCO => next_reg_a_cry_20);
    
    sum0_4_cry_0_998 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[17]\, C => 
        \R0_data[8]\, Y => \SIG0_0[27]\);
    
    sum3_cry_25 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[25]\, B => Wt_data(25), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_24\, S => 
        \sum3[25]\, Y => OPEN, FCO => \sum3_cry_25\);
    
    \next_reg_g[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[4]\, B => N6_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[4]_net_1\);
    
    sum3_4_cry_29 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[29]\, B => m304, C => i3_mux_1, D => 
        Kt_addr(5), FCI => \sum3_4_cry_28\, S => \sum3_4[29]\, Y
         => OPEN, FCO => \sum3_4_cry_29\);
    
    sum3_6_cry_23 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[23]\, B => \R4_data[2]\, C => 
        \R4_data[16]\, D => \R4_data[29]\, FCI => \sum3_6_cry_22\, 
        S => \sum3_6[23]\, Y => OPEN, FCO => \sum3_6_cry_23\);
    
    \next_reg_g[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(22), B => \R5_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[22]_net_1\);
    
    \next_reg_b[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(24), B => \R0_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[24]_net_1\);
    
    \reg_e[3]\ : SLE
      port map(D => \next_reg_e[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[3]\);
    
    \SIG0[5]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[18]\, C => 
        \R0_data[7]\, Y => \SIG0[5]_net_1\);
    
    \next_reg_g[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(17), B => \R5_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[17]_net_1\);
    
    \next_reg_g[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(15), B => \R5_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[15]_net_1\);
    
    sum0_4_cry_0_1006 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[21]\, B => \R0_data[9]\, C => 
        \R0_data[0]\, Y => \SIG0_0[19]\);
    
    sum3_6_0_cry_7 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[7]\, B => \R4_data[7]\, C => 
        \R5_data[7]\, D => \R6_data[7]\, FCI => \sum3_6_0_cry_6\, 
        S => \sum3_6_0[7]\, Y => OPEN, FCO => \sum3_6_0_cry_7\);
    
    sum3_4_cry_26 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[26]\, B => m281_ns, C => m285, D => 
        Kt_addr(5), FCI => \sum3_4_cry_25\, S => \sum3_4[26]\, Y
         => OPEN, FCO => \sum3_4_cry_26\);
    
    \next_reg_f[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(24), B => \R4_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[24]_net_1\);
    
    \reg_f[6]\ : SLE
      port map(D => \next_reg_f[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[6]\);
    
    sum3_axb_0 : CFG2
      generic map(INIT => x"6")

      port map(A => sum3_4_cry_0_Y, B => Wt_data(0), Y => 
        \sum3[0]\);
    
    \next_reg_h[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(30), B => \R6_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[30]_net_1\);
    
    sum3_6_cry_28 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[28]\, B => \R4_data[2]\, C => 
        \R4_data[7]\, D => \R4_data[21]\, FCI => \sum3_6_cry_27\, 
        S => \sum3_6[28]\, Y => OPEN, FCO => \sum3_6_cry_28\);
    
    \reg_a[9]\ : SLE
      port map(D => \next_reg_a[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[9]\);
    
    \SIG0[3]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[16]\, C => 
        \R0_data[5]\, Y => \SIG0[3]_net_1\);
    
    \reg_c[17]\ : SLE
      port map(D => \next_reg_c[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[17]\);
    
    \reg_b[24]\ : SLE
      port map(D => \next_reg_b[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[24]\);
    
    sum0_4_axb_1 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[1]\, B => \R1_data[1]\, C => 
        \R0_data[1]\, D => \SIG0[1]_net_1\, Y => \sum0_4_axb_1\);
    
    \reg_g[26]\ : SLE
      port map(D => \next_reg_g[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[26]\);
    
    \reg_a[6]\ : SLE
      port map(D => \next_reg_a[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[6]\);
    
    \SIG0[22]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[24]\, B => \R0_data[3]\, C => 
        \R0_data[12]\, Y => \SIG0[22]_net_1\);
    
    \reg_d[19]\ : SLE
      port map(D => \next_reg_d[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[19]\);
    
    \reg_d[5]\ : SLE
      port map(D => \next_reg_d[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R3_data[5]\);
    
    \reg_a[4]\ : SLE
      port map(D => \next_reg_a[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[4]\);
    
    \reg_f[20]\ : SLE
      port map(D => \next_reg_f[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[20]\);
    
    next_reg_a_cry_10_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[10]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[10]\, D => N0_data(10), FCI => next_reg_a_cry_9, S
         => \next_reg_a[10]\, Y => OPEN, FCO => next_reg_a_cry_10);
    
    \next_reg_h[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(27), B => \R6_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[27]_net_1\);
    
    next_reg_e_cry_30_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[30]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(30), D => \R3_data[30]\, FCI => next_reg_e_cry_29, 
        S => \next_reg_e[30]\, Y => OPEN, FCO => 
        next_reg_e_cry_30);
    
    \reg_c[0]\ : SLE
      port map(D => \next_reg_c[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R2_data[0]\);
    
    \next_reg_h[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(25), B => \R6_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[25]_net_1\);
    
    \next_reg_d[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[4]\, B => N3_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[4]_net_1\);
    
    \next_reg_f[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(10), B => \R4_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[10]_net_1\);
    
    \reg_g[7]\ : SLE
      port map(D => \next_reg_g[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[7]\);
    
    sum0_4_axb_14 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[14]\, B => \R1_data[14]\, C => 
        \R0_data[14]\, D => \SIG0[14]_net_1\, Y => 
        \sum0_4_axb_14\);
    
    sum3_cry_13 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[13]\, B => Wt_data(13), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_12\, S => 
        \sum3[13]\, Y => OPEN, FCO => \sum3_cry_13\);
    
    \reg_e[13]\ : SLE
      port map(D => \next_reg_e[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R4_data[13]\);
    
    next_reg_a_cry_9_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[9]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[9]\, D => N0_data(9), FCI => next_reg_a_cry_8, S
         => \next_reg_a[9]\, Y => OPEN, FCO => next_reg_a_cry_9);
    
    next_reg_a_cry_30_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[30]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[30]\, D => N0_data(30), FCI => next_reg_a_cry_29, S
         => \next_reg_a[30]\, Y => OPEN, FCO => next_reg_a_cry_30);
    
    sum3_4_axb_0 : CFG2
      generic map(INIT => x"6")

      port map(A => Kt_data_0, B => sum3_6_cry_0_Y, Y => 
        \sum3_4[0]\);
    
    \reg_g[28]\ : SLE
      port map(D => \next_reg_g[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R6_data[28]\);
    
    next_reg_e_cry_16_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[16]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(16), D => \R3_data[16]\, FCI => next_reg_e_cry_15, 
        S => \next_reg_e[16]\, Y => OPEN, FCO => 
        next_reg_e_cry_16);
    
    \reg_h[5]\ : SLE
      port map(D => \next_reg_h[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R7_data[5]\);
    
    \next_reg_f[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[5]\, B => N5_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[5]_net_1\);
    
    sum3_4_cry_22 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[22]\, B => m250_am, C => m250_bm, D
         => Kt_addr(5), FCI => \sum3_4_cry_21\, S => \sum3_4[22]\, 
        Y => OPEN, FCO => \sum3_4_cry_22\);
    
    \SIG0[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[13]\, B => \R0_data[1]\, C => 
        \R0_data[24]\, Y => \SIG0[11]_net_1\);
    
    \reg_f[31]\ : SLE
      port map(D => \next_reg_f[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R5_data[31]\);
    
    \next_reg_c[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(29), B => \R1_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[29]_net_1\);
    
    \reg_b[10]\ : SLE
      port map(D => \next_reg_b[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R1_data[10]\);
    
    \reg_a[1]\ : SLE
      port map(D => \next_reg_a[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => core_ce_o_iv_i_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \R0_data[1]\);
    
    sum0_4_axb_17 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[17]\, B => \R1_data[17]\, C => 
        \R0_data[17]\, D => \SIG0[17]_net_1\, Y => 
        \sum0_4_axb_17\);
    
    sum3_4_cry_3 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[3]\, B => m62_am, C => m62_bm, D => 
        Kt_addr_5_rep1, FCI => \sum3_4_cry_2\, S => \sum3_4[3]\, 
        Y => OPEN, FCO => \sum3_4_cry_3\);
    
    \next_reg_f[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(12), B => \R4_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[12]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_regs is

    port( SHA256_BLOCK_0_H0_o          : out   std_logic_vector(31 downto 0);
          N0_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H1_o          : out   std_logic_vector(31 downto 0);
          N1_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H2_o          : out   std_logic_vector(31 downto 0);
          N2_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H3_o          : out   std_logic_vector(31 downto 0);
          N3_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H4_o          : out   std_logic_vector(31 downto 0);
          N4_data                      : out   std_logic_vector(31 downto 1);
          N5_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H5_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o          : out   std_logic_vector(31 downto 0);
          N6_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H7_o          : out   std_logic_vector(31 downto 0);
          N7_data                      : out   std_logic_vector(31 downto 1);
          hash_control_st_reg_i        : in    std_logic_vector(6 to 6);
          R0_data                      : in    std_logic_vector(31 downto 0);
          R1_data                      : in    std_logic_vector(31 downto 0);
          R2_data                      : in    std_logic_vector(31 downto 0);
          R3_data                      : in    std_logic_vector(31 downto 0);
          R4_data                      : in    std_logic_vector(31 downto 0);
          R5_data                      : in    std_logic_vector(31 downto 0);
          R6_data                      : in    std_logic_vector(31 downto 0);
          R7_data                      : in    std_logic_vector(31 downto 0);
          sha256_system_sb_0_FIC_0_CLK : in    std_logic;
          N_168_i_0                    : in    std_logic;
          next_reg_H0_cry_0_0_Y        : out   std_logic;
          next_reg_H1_cry_0_0_Y        : out   std_logic;
          next_reg_H2_cry_0_0_Y        : out   std_logic;
          next_reg_H3_cry_0_0_Y        : out   std_logic;
          next_reg_H4_cry_0_0_Y        : out   std_logic;
          next_reg_H5_cry_0_0_Y        : out   std_logic;
          next_reg_H6_cry_0_0_Y        : out   std_logic;
          next_reg_H7_cry_0_0_Y        : out   std_logic
        );

end sha256_regs;

architecture DEF_ARCH of sha256_regs is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \SHA256_BLOCK_0_H0_o[21]\, VCC_net_1, \N0_data[21]\, 
        GND_net_1, \SHA256_BLOCK_0_H0_o[22]\, \N0_data[22]\, 
        \SHA256_BLOCK_0_H0_o[23]\, \N0_data[23]\, 
        \SHA256_BLOCK_0_H0_o[24]\, \N0_data[24]\, 
        \SHA256_BLOCK_0_H0_o[25]\, \N0_data[25]\, 
        \SHA256_BLOCK_0_H0_o[26]\, \N0_data[26]\, 
        \SHA256_BLOCK_0_H0_o[27]\, \N0_data[27]\, 
        \SHA256_BLOCK_0_H0_o[28]\, \N0_data[28]\, 
        \SHA256_BLOCK_0_H0_o[29]\, \N0_data[29]\, 
        \SHA256_BLOCK_0_H0_o[30]\, \N0_data[30]\, 
        \SHA256_BLOCK_0_H0_o[31]\, \N0_data[31]\, 
        \SHA256_BLOCK_0_H0_o[6]\, \N0_data[6]\, 
        \SHA256_BLOCK_0_H0_o[7]\, \N0_data[7]\, 
        \SHA256_BLOCK_0_H0_o[8]\, \N0_data[8]\, 
        \SHA256_BLOCK_0_H0_o[9]\, \N0_data[9]\, 
        \SHA256_BLOCK_0_H0_o[10]\, \N0_data[10]\, 
        \SHA256_BLOCK_0_H0_o[11]\, \N0_data[11]\, 
        \SHA256_BLOCK_0_H0_o[12]\, \N0_data[12]\, 
        \SHA256_BLOCK_0_H0_o[13]\, \N0_data[13]\, 
        \SHA256_BLOCK_0_H0_o[14]\, \N0_data[14]\, 
        \SHA256_BLOCK_0_H0_o[15]\, \N0_data[15]\, 
        \SHA256_BLOCK_0_H0_o[16]\, \N0_data[16]\, 
        \SHA256_BLOCK_0_H0_o[17]\, \N0_data[17]\, 
        \SHA256_BLOCK_0_H0_o[18]\, \N0_data[18]\, 
        \SHA256_BLOCK_0_H0_o[19]\, \N0_data[19]\, 
        \SHA256_BLOCK_0_H0_o[20]\, \N0_data[20]\, 
        \SHA256_BLOCK_0_H1_o[23]\, \N1_data[23]\, 
        \SHA256_BLOCK_0_H1_o[24]\, \N1_data[24]\, 
        \SHA256_BLOCK_0_H1_o[25]\, \N1_data[25]\, 
        \SHA256_BLOCK_0_H1_o[26]\, \N1_data[26]\, 
        \SHA256_BLOCK_0_H1_o[27]\, \N1_data[27]\, 
        \SHA256_BLOCK_0_H1_o[28]\, \N1_data[28]\, 
        \SHA256_BLOCK_0_H1_o[29]\, \N1_data[29]\, 
        \SHA256_BLOCK_0_H1_o[30]\, \N1_data[30]\, 
        \SHA256_BLOCK_0_H1_o[31]\, \N1_data[31]\, 
        \SHA256_BLOCK_0_H0_o[0]\, \next_reg_H0_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H0_o[1]\, \N0_data[1]\, 
        \SHA256_BLOCK_0_H0_o[2]\, \N0_data[2]\, 
        \SHA256_BLOCK_0_H0_o[3]\, \N0_data[3]\, 
        \SHA256_BLOCK_0_H0_o[4]\, \N0_data[4]\, 
        \SHA256_BLOCK_0_H0_o[5]\, \N0_data[5]\, 
        \SHA256_BLOCK_0_H1_o[8]\, \N1_data[8]\, 
        \SHA256_BLOCK_0_H1_o[9]\, \N1_data[9]\, 
        \SHA256_BLOCK_0_H1_o[10]\, \N1_data[10]\, 
        \SHA256_BLOCK_0_H1_o[11]\, \N1_data[11]\, 
        \SHA256_BLOCK_0_H1_o[12]\, \N1_data[12]\, 
        \SHA256_BLOCK_0_H1_o[13]\, \N1_data[13]\, 
        \SHA256_BLOCK_0_H1_o[14]\, \N1_data[14]\, 
        \SHA256_BLOCK_0_H1_o[15]\, \N1_data[15]\, 
        \SHA256_BLOCK_0_H1_o[16]\, \N1_data[16]\, 
        \SHA256_BLOCK_0_H1_o[17]\, \N1_data[17]\, 
        \SHA256_BLOCK_0_H1_o[18]\, \N1_data[18]\, 
        \SHA256_BLOCK_0_H1_o[19]\, \N1_data[19]\, 
        \SHA256_BLOCK_0_H1_o[20]\, \N1_data[20]\, 
        \SHA256_BLOCK_0_H1_o[21]\, \N1_data[21]\, 
        \SHA256_BLOCK_0_H1_o[22]\, \N1_data[22]\, 
        \SHA256_BLOCK_0_H2_o[25]\, \N2_data[25]\, 
        \SHA256_BLOCK_0_H2_o[26]\, \N2_data[26]\, 
        \SHA256_BLOCK_0_H2_o[27]\, \N2_data[27]\, 
        \SHA256_BLOCK_0_H2_o[28]\, \N2_data[28]\, 
        \SHA256_BLOCK_0_H2_o[29]\, \N2_data[29]\, 
        \SHA256_BLOCK_0_H2_o[30]\, \N2_data[30]\, 
        \SHA256_BLOCK_0_H2_o[31]\, \N2_data[31]\, 
        \SHA256_BLOCK_0_H1_o[0]\, \next_reg_H1_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H1_o[1]\, \N1_data[1]\, 
        \SHA256_BLOCK_0_H1_o[2]\, \N1_data[2]\, 
        \SHA256_BLOCK_0_H1_o[3]\, \N1_data[3]\, 
        \SHA256_BLOCK_0_H1_o[4]\, \N1_data[4]\, 
        \SHA256_BLOCK_0_H1_o[5]\, \N1_data[5]\, 
        \SHA256_BLOCK_0_H1_o[6]\, \N1_data[6]\, 
        \SHA256_BLOCK_0_H1_o[7]\, \N1_data[7]\, 
        \SHA256_BLOCK_0_H2_o[10]\, \N2_data[10]\, 
        \SHA256_BLOCK_0_H2_o[11]\, \N2_data[11]\, 
        \SHA256_BLOCK_0_H2_o[12]\, \N2_data[12]\, 
        \SHA256_BLOCK_0_H2_o[13]\, \N2_data[13]\, 
        \SHA256_BLOCK_0_H2_o[14]\, \N2_data[14]\, 
        \SHA256_BLOCK_0_H2_o[15]\, \N2_data[15]\, 
        \SHA256_BLOCK_0_H2_o[16]\, \N2_data[16]\, 
        \SHA256_BLOCK_0_H2_o[17]\, \N2_data[17]\, 
        \SHA256_BLOCK_0_H2_o[18]\, \N2_data[18]\, 
        \SHA256_BLOCK_0_H2_o[19]\, \N2_data[19]\, 
        \SHA256_BLOCK_0_H2_o[20]\, \N2_data[20]\, 
        \SHA256_BLOCK_0_H2_o[21]\, \N2_data[21]\, 
        \SHA256_BLOCK_0_H2_o[22]\, \N2_data[22]\, 
        \SHA256_BLOCK_0_H2_o[23]\, \N2_data[23]\, 
        \SHA256_BLOCK_0_H2_o[24]\, \N2_data[24]\, 
        \SHA256_BLOCK_0_H3_o[27]\, \N3_data[27]\, 
        \SHA256_BLOCK_0_H3_o[28]\, \N3_data[28]\, 
        \SHA256_BLOCK_0_H3_o[29]\, \N3_data[29]\, 
        \SHA256_BLOCK_0_H3_o[30]\, \N3_data[30]\, 
        \SHA256_BLOCK_0_H3_o[31]\, \N3_data[31]\, 
        \SHA256_BLOCK_0_H2_o[0]\, \next_reg_H2_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H2_o[1]\, \N2_data[1]\, 
        \SHA256_BLOCK_0_H2_o[2]\, \N2_data[2]\, 
        \SHA256_BLOCK_0_H2_o[3]\, \N2_data[3]\, 
        \SHA256_BLOCK_0_H2_o[4]\, \N2_data[4]\, 
        \SHA256_BLOCK_0_H2_o[5]\, \N2_data[5]\, 
        \SHA256_BLOCK_0_H2_o[6]\, \N2_data[6]\, 
        \SHA256_BLOCK_0_H2_o[7]\, \N2_data[7]\, 
        \SHA256_BLOCK_0_H2_o[8]\, \N2_data[8]\, 
        \SHA256_BLOCK_0_H2_o[9]\, \N2_data[9]\, 
        \SHA256_BLOCK_0_H3_o[12]\, \N3_data[12]\, 
        \SHA256_BLOCK_0_H3_o[13]\, \N3_data[13]\, 
        \SHA256_BLOCK_0_H3_o[14]\, \N3_data[14]\, 
        \SHA256_BLOCK_0_H3_o[15]\, \N3_data[15]\, 
        \SHA256_BLOCK_0_H3_o[16]\, \N3_data[16]\, 
        \SHA256_BLOCK_0_H3_o[17]\, \N3_data[17]\, 
        \SHA256_BLOCK_0_H3_o[18]\, \N3_data[18]\, 
        \SHA256_BLOCK_0_H3_o[19]\, \N3_data[19]\, 
        \SHA256_BLOCK_0_H3_o[20]\, \N3_data[20]\, 
        \SHA256_BLOCK_0_H3_o[21]\, \N3_data[21]\, 
        \SHA256_BLOCK_0_H3_o[22]\, \N3_data[22]\, 
        \SHA256_BLOCK_0_H3_o[23]\, \N3_data[23]\, 
        \SHA256_BLOCK_0_H3_o[24]\, \N3_data[24]\, 
        \SHA256_BLOCK_0_H3_o[25]\, \N3_data[25]\, 
        \SHA256_BLOCK_0_H3_o[26]\, \N3_data[26]\, 
        \SHA256_BLOCK_0_H4_o[29]\, \N4_data[29]\, 
        \SHA256_BLOCK_0_H4_o[30]\, \N4_data[30]\, 
        \SHA256_BLOCK_0_H4_o[31]\, \N4_data[31]\, 
        \SHA256_BLOCK_0_H3_o[0]\, \next_reg_H3_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H3_o[1]\, \N3_data[1]\, 
        \SHA256_BLOCK_0_H3_o[2]\, \N3_data[2]\, 
        \SHA256_BLOCK_0_H3_o[3]\, \N3_data[3]\, 
        \SHA256_BLOCK_0_H3_o[4]\, \N3_data[4]\, 
        \SHA256_BLOCK_0_H3_o[5]\, \N3_data[5]\, 
        \SHA256_BLOCK_0_H3_o[6]\, \N3_data[6]\, 
        \SHA256_BLOCK_0_H3_o[7]\, \N3_data[7]\, 
        \SHA256_BLOCK_0_H3_o[8]\, \N3_data[8]\, 
        \SHA256_BLOCK_0_H3_o[9]\, \N3_data[9]\, 
        \SHA256_BLOCK_0_H3_o[10]\, \N3_data[10]\, 
        \SHA256_BLOCK_0_H3_o[11]\, \N3_data[11]\, 
        \SHA256_BLOCK_0_H4_o[14]\, \N4_data[14]\, 
        \SHA256_BLOCK_0_H4_o[15]\, \N4_data[15]\, 
        \SHA256_BLOCK_0_H4_o[16]\, \N4_data[16]\, 
        \SHA256_BLOCK_0_H4_o[17]\, \N4_data[17]\, 
        \SHA256_BLOCK_0_H4_o[18]\, \N4_data[18]\, 
        \SHA256_BLOCK_0_H4_o[19]\, \N4_data[19]\, 
        \SHA256_BLOCK_0_H4_o[20]\, \N4_data[20]\, 
        \SHA256_BLOCK_0_H4_o[21]\, \N4_data[21]\, 
        \SHA256_BLOCK_0_H4_o[22]\, \N4_data[22]\, 
        \SHA256_BLOCK_0_H4_o[23]\, \N4_data[23]\, 
        \SHA256_BLOCK_0_H4_o[24]\, \N4_data[24]\, 
        \SHA256_BLOCK_0_H4_o[25]\, \N4_data[25]\, 
        \SHA256_BLOCK_0_H4_o[26]\, \N4_data[26]\, 
        \SHA256_BLOCK_0_H4_o[27]\, \N4_data[27]\, 
        \SHA256_BLOCK_0_H4_o[28]\, \N4_data[28]\, 
        \SHA256_BLOCK_0_H5_o[31]\, \N5_data[31]\, 
        \SHA256_BLOCK_0_H4_o[0]\, \next_reg_H4_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H4_o[1]\, \N4_data[1]\, 
        \SHA256_BLOCK_0_H4_o[2]\, \N4_data[2]\, 
        \SHA256_BLOCK_0_H4_o[3]\, \N4_data[3]\, 
        \SHA256_BLOCK_0_H4_o[4]\, \N4_data[4]\, 
        \SHA256_BLOCK_0_H4_o[5]\, \N4_data[5]\, 
        \SHA256_BLOCK_0_H4_o[6]\, \N4_data[6]\, 
        \SHA256_BLOCK_0_H4_o[7]\, \N4_data[7]\, 
        \SHA256_BLOCK_0_H4_o[8]\, \N4_data[8]\, 
        \SHA256_BLOCK_0_H4_o[9]\, \N4_data[9]\, 
        \SHA256_BLOCK_0_H4_o[10]\, \N4_data[10]\, 
        \SHA256_BLOCK_0_H4_o[11]\, \N4_data[11]\, 
        \SHA256_BLOCK_0_H4_o[12]\, \N4_data[12]\, 
        \SHA256_BLOCK_0_H4_o[13]\, \N4_data[13]\, 
        \SHA256_BLOCK_0_H5_o[16]\, \N5_data[16]\, 
        \SHA256_BLOCK_0_H5_o[17]\, \N5_data[17]\, 
        \SHA256_BLOCK_0_H5_o[18]\, \N5_data[18]\, 
        \SHA256_BLOCK_0_H5_o[19]\, \N5_data[19]\, 
        \SHA256_BLOCK_0_H5_o[20]\, \N5_data[20]\, 
        \SHA256_BLOCK_0_H5_o[21]\, \N5_data[21]\, 
        \SHA256_BLOCK_0_H5_o[22]\, \N5_data[22]\, 
        \SHA256_BLOCK_0_H5_o[23]\, \N5_data[23]\, 
        \SHA256_BLOCK_0_H5_o[24]\, \N5_data[24]\, 
        \SHA256_BLOCK_0_H5_o[25]\, \N5_data[25]\, 
        \SHA256_BLOCK_0_H5_o[26]\, \N5_data[26]\, 
        \SHA256_BLOCK_0_H5_o[27]\, \N5_data[27]\, 
        \SHA256_BLOCK_0_H5_o[28]\, \N5_data[28]\, 
        \SHA256_BLOCK_0_H5_o[29]\, \N5_data[29]\, 
        \SHA256_BLOCK_0_H5_o[30]\, \N5_data[30]\, 
        \SHA256_BLOCK_0_H5_o[1]\, \N5_data[1]\, 
        \SHA256_BLOCK_0_H5_o[2]\, \N5_data[2]\, 
        \SHA256_BLOCK_0_H5_o[3]\, \N5_data[3]\, 
        \SHA256_BLOCK_0_H5_o[4]\, \N5_data[4]\, 
        \SHA256_BLOCK_0_H5_o[5]\, \N5_data[5]\, 
        \SHA256_BLOCK_0_H5_o[6]\, \N5_data[6]\, 
        \SHA256_BLOCK_0_H5_o[7]\, \N5_data[7]\, 
        \SHA256_BLOCK_0_H5_o[8]\, \N5_data[8]\, 
        \SHA256_BLOCK_0_H5_o[9]\, \N5_data[9]\, 
        \SHA256_BLOCK_0_H5_o[10]\, \N5_data[10]\, 
        \SHA256_BLOCK_0_H5_o[11]\, \N5_data[11]\, 
        \SHA256_BLOCK_0_H5_o[12]\, \N5_data[12]\, 
        \SHA256_BLOCK_0_H5_o[13]\, \N5_data[13]\, 
        \SHA256_BLOCK_0_H5_o[14]\, \N5_data[14]\, 
        \SHA256_BLOCK_0_H5_o[15]\, \N5_data[15]\, 
        \SHA256_BLOCK_0_H6_o[18]\, \N6_data[18]\, 
        \SHA256_BLOCK_0_H6_o[19]\, \N6_data[19]\, 
        \SHA256_BLOCK_0_H6_o[20]\, \N6_data[20]\, 
        \SHA256_BLOCK_0_H6_o[21]\, \N6_data[21]\, 
        \SHA256_BLOCK_0_H6_o[22]\, \N6_data[22]\, 
        \SHA256_BLOCK_0_H6_o[23]\, \N6_data[23]\, 
        \SHA256_BLOCK_0_H6_o[24]\, \N6_data[24]\, 
        \SHA256_BLOCK_0_H6_o[25]\, \N6_data[25]\, 
        \SHA256_BLOCK_0_H6_o[26]\, \N6_data[26]\, 
        \SHA256_BLOCK_0_H6_o[27]\, \N6_data[27]\, 
        \SHA256_BLOCK_0_H6_o[28]\, \N6_data[28]\, 
        \SHA256_BLOCK_0_H6_o[29]\, \N6_data[29]\, 
        \SHA256_BLOCK_0_H6_o[30]\, \N6_data[30]\, 
        \SHA256_BLOCK_0_H6_o[31]\, \N6_data[31]\, 
        \SHA256_BLOCK_0_H5_o[0]\, \next_reg_H5_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H6_o[3]\, \N6_data[3]\, 
        \SHA256_BLOCK_0_H6_o[4]\, \N6_data[4]\, 
        \SHA256_BLOCK_0_H6_o[5]\, \N6_data[5]\, 
        \SHA256_BLOCK_0_H6_o[6]\, \N6_data[6]\, 
        \SHA256_BLOCK_0_H6_o[7]\, \N6_data[7]\, 
        \SHA256_BLOCK_0_H6_o[8]\, \N6_data[8]\, 
        \SHA256_BLOCK_0_H6_o[9]\, \N6_data[9]\, 
        \SHA256_BLOCK_0_H6_o[10]\, \N6_data[10]\, 
        \SHA256_BLOCK_0_H6_o[11]\, \N6_data[11]\, 
        \SHA256_BLOCK_0_H6_o[12]\, \N6_data[12]\, 
        \SHA256_BLOCK_0_H6_o[13]\, \N6_data[13]\, 
        \SHA256_BLOCK_0_H6_o[14]\, \N6_data[14]\, 
        \SHA256_BLOCK_0_H6_o[15]\, \N6_data[15]\, 
        \SHA256_BLOCK_0_H6_o[16]\, \N6_data[16]\, 
        \SHA256_BLOCK_0_H6_o[17]\, \N6_data[17]\, 
        \SHA256_BLOCK_0_H7_o[20]\, \N7_data[20]\, 
        \SHA256_BLOCK_0_H7_o[21]\, \N7_data[21]\, 
        \SHA256_BLOCK_0_H7_o[22]\, \N7_data[22]\, 
        \SHA256_BLOCK_0_H7_o[23]\, \N7_data[23]\, 
        \SHA256_BLOCK_0_H7_o[24]\, \N7_data[24]\, 
        \SHA256_BLOCK_0_H7_o[25]\, \N7_data[25]\, 
        \SHA256_BLOCK_0_H7_o[26]\, \N7_data[26]\, 
        \SHA256_BLOCK_0_H7_o[27]\, \N7_data[27]\, 
        \SHA256_BLOCK_0_H7_o[28]\, \N7_data[28]\, 
        \SHA256_BLOCK_0_H7_o[29]\, \N7_data[29]\, 
        \SHA256_BLOCK_0_H7_o[30]\, \N7_data[30]\, 
        \SHA256_BLOCK_0_H7_o[31]\, \N7_data[31]\, 
        \SHA256_BLOCK_0_H6_o[0]\, \next_reg_H6_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H6_o[1]\, \N6_data[1]\, 
        \SHA256_BLOCK_0_H6_o[2]\, \N6_data[2]\, 
        \SHA256_BLOCK_0_H7_o[5]\, \N7_data[5]\, 
        \SHA256_BLOCK_0_H7_o[6]\, \N7_data[6]\, 
        \SHA256_BLOCK_0_H7_o[7]\, \N7_data[7]\, 
        \SHA256_BLOCK_0_H7_o[8]\, \N7_data[8]\, 
        \SHA256_BLOCK_0_H7_o[9]\, \N7_data[9]\, 
        \SHA256_BLOCK_0_H7_o[10]\, \N7_data[10]\, 
        \SHA256_BLOCK_0_H7_o[11]\, \N7_data[11]\, 
        \SHA256_BLOCK_0_H7_o[12]\, \N7_data[12]\, 
        \SHA256_BLOCK_0_H7_o[13]\, \N7_data[13]\, 
        \SHA256_BLOCK_0_H7_o[14]\, \N7_data[14]\, 
        \SHA256_BLOCK_0_H7_o[15]\, \N7_data[15]\, 
        \SHA256_BLOCK_0_H7_o[16]\, \N7_data[16]\, 
        \SHA256_BLOCK_0_H7_o[17]\, \N7_data[17]\, 
        \SHA256_BLOCK_0_H7_o[18]\, \N7_data[18]\, 
        \SHA256_BLOCK_0_H7_o[19]\, \N7_data[19]\, 
        \SHA256_BLOCK_0_H7_o[0]\, \next_reg_H7_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H7_o[1]\, \N7_data[1]\, 
        \SHA256_BLOCK_0_H7_o[2]\, \N7_data[2]\, 
        \SHA256_BLOCK_0_H7_o[3]\, \N7_data[3]\, 
        \SHA256_BLOCK_0_H7_o[4]\, \N7_data[4]\, next_reg_H0_cry_0, 
        next_reg_H0_cry_1, next_reg_H0_cry_2, next_reg_H0_cry_3, 
        next_reg_H0_cry_4, next_reg_H0_cry_5, next_reg_H0_cry_6, 
        next_reg_H0_cry_7, next_reg_H0_cry_8, next_reg_H0_cry_9, 
        next_reg_H0_cry_10, next_reg_H0_cry_11, 
        next_reg_H0_cry_12, next_reg_H0_cry_13, 
        next_reg_H0_cry_14, next_reg_H0_cry_15, 
        next_reg_H0_cry_16, next_reg_H0_cry_17, 
        next_reg_H0_cry_18, next_reg_H0_cry_19, 
        next_reg_H0_cry_20, next_reg_H0_cry_21, 
        next_reg_H0_cry_22, next_reg_H0_cry_23, 
        next_reg_H0_cry_24, next_reg_H0_cry_25, 
        next_reg_H0_cry_26, next_reg_H0_cry_27, 
        next_reg_H0_cry_28, next_reg_H0_cry_29, 
        next_reg_H0_cry_30, next_reg_H1_cry_0, next_reg_H1_cry_1, 
        next_reg_H1_cry_2, next_reg_H1_cry_3, next_reg_H1_cry_4, 
        next_reg_H1_cry_5, next_reg_H1_cry_6, next_reg_H1_cry_7, 
        next_reg_H1_cry_8, next_reg_H1_cry_9, next_reg_H1_cry_10, 
        next_reg_H1_cry_11, next_reg_H1_cry_12, 
        next_reg_H1_cry_13, next_reg_H1_cry_14, 
        next_reg_H1_cry_15, next_reg_H1_cry_16, 
        next_reg_H1_cry_17, next_reg_H1_cry_18, 
        next_reg_H1_cry_19, next_reg_H1_cry_20, 
        next_reg_H1_cry_21, next_reg_H1_cry_22, 
        next_reg_H1_cry_23, next_reg_H1_cry_24, 
        next_reg_H1_cry_25, next_reg_H1_cry_26, 
        next_reg_H1_cry_27, next_reg_H1_cry_28, 
        next_reg_H1_cry_29, next_reg_H1_cry_30, next_reg_H2_cry_0, 
        next_reg_H2_cry_1, next_reg_H2_cry_2, next_reg_H2_cry_3, 
        next_reg_H2_cry_4, next_reg_H2_cry_5, next_reg_H2_cry_6, 
        next_reg_H2_cry_7, next_reg_H2_cry_8, next_reg_H2_cry_9, 
        next_reg_H2_cry_10, next_reg_H2_cry_11, 
        next_reg_H2_cry_12, next_reg_H2_cry_13, 
        next_reg_H2_cry_14, next_reg_H2_cry_15, 
        next_reg_H2_cry_16, next_reg_H2_cry_17, 
        next_reg_H2_cry_18, next_reg_H2_cry_19, 
        next_reg_H2_cry_20, next_reg_H2_cry_21, 
        next_reg_H2_cry_22, next_reg_H2_cry_23, 
        next_reg_H2_cry_24, next_reg_H2_cry_25, 
        next_reg_H2_cry_26, next_reg_H2_cry_27, 
        next_reg_H2_cry_28, next_reg_H2_cry_29, 
        next_reg_H2_cry_30, next_reg_H3_cry_0, next_reg_H3_cry_1, 
        next_reg_H3_cry_2, next_reg_H3_cry_3, next_reg_H3_cry_4, 
        next_reg_H3_cry_5, next_reg_H3_cry_6, next_reg_H3_cry_7, 
        next_reg_H3_cry_8, next_reg_H3_cry_9, next_reg_H3_cry_10, 
        next_reg_H3_cry_11, next_reg_H3_cry_12, 
        next_reg_H3_cry_13, next_reg_H3_cry_14, 
        next_reg_H3_cry_15, next_reg_H3_cry_16, 
        next_reg_H3_cry_17, next_reg_H3_cry_18, 
        next_reg_H3_cry_19, next_reg_H3_cry_20, 
        next_reg_H3_cry_21, next_reg_H3_cry_22, 
        next_reg_H3_cry_23, next_reg_H3_cry_24, 
        next_reg_H3_cry_25, next_reg_H3_cry_26, 
        next_reg_H3_cry_27, next_reg_H3_cry_28, 
        next_reg_H3_cry_29, next_reg_H3_cry_30, next_reg_H4_cry_0, 
        next_reg_H4_cry_1, next_reg_H4_cry_2, next_reg_H4_cry_3, 
        next_reg_H4_cry_4, next_reg_H4_cry_5, next_reg_H4_cry_6, 
        next_reg_H4_cry_7, next_reg_H4_cry_8, next_reg_H4_cry_9, 
        next_reg_H4_cry_10, next_reg_H4_cry_11, 
        next_reg_H4_cry_12, next_reg_H4_cry_13, 
        next_reg_H4_cry_14, next_reg_H4_cry_15, 
        next_reg_H4_cry_16, next_reg_H4_cry_17, 
        next_reg_H4_cry_18, next_reg_H4_cry_19, 
        next_reg_H4_cry_20, next_reg_H4_cry_21, 
        next_reg_H4_cry_22, next_reg_H4_cry_23, 
        next_reg_H4_cry_24, next_reg_H4_cry_25, 
        next_reg_H4_cry_26, next_reg_H4_cry_27, 
        next_reg_H4_cry_28, next_reg_H4_cry_29, 
        next_reg_H4_cry_30, next_reg_H5_cry_0, next_reg_H5_cry_1, 
        next_reg_H5_cry_2, next_reg_H5_cry_3, next_reg_H5_cry_4, 
        next_reg_H5_cry_5, next_reg_H5_cry_6, next_reg_H5_cry_7, 
        next_reg_H5_cry_8, next_reg_H5_cry_9, next_reg_H5_cry_10, 
        next_reg_H5_cry_11, next_reg_H5_cry_12, 
        next_reg_H5_cry_13, next_reg_H5_cry_14, 
        next_reg_H5_cry_15, next_reg_H5_cry_16, 
        next_reg_H5_cry_17, next_reg_H5_cry_18, 
        next_reg_H5_cry_19, next_reg_H5_cry_20, 
        next_reg_H5_cry_21, next_reg_H5_cry_22, 
        next_reg_H5_cry_23, next_reg_H5_cry_24, 
        next_reg_H5_cry_25, next_reg_H5_cry_26, 
        next_reg_H5_cry_27, next_reg_H5_cry_28, 
        next_reg_H5_cry_29, next_reg_H5_cry_30, next_reg_H6_cry_0, 
        next_reg_H6_cry_1, next_reg_H6_cry_2, next_reg_H6_cry_3, 
        next_reg_H6_cry_4, next_reg_H6_cry_5, next_reg_H6_cry_6, 
        next_reg_H6_cry_7, next_reg_H6_cry_8, next_reg_H6_cry_9, 
        next_reg_H6_cry_10, next_reg_H6_cry_11, 
        next_reg_H6_cry_12, next_reg_H6_cry_13, 
        next_reg_H6_cry_14, next_reg_H6_cry_15, 
        next_reg_H6_cry_16, next_reg_H6_cry_17, 
        next_reg_H6_cry_18, next_reg_H6_cry_19, 
        next_reg_H6_cry_20, next_reg_H6_cry_21, 
        next_reg_H6_cry_22, next_reg_H6_cry_23, 
        next_reg_H6_cry_24, next_reg_H6_cry_25, 
        next_reg_H6_cry_26, next_reg_H6_cry_27, 
        next_reg_H6_cry_28, next_reg_H6_cry_29, 
        next_reg_H6_cry_30, next_reg_H7_cry_0, next_reg_H7_cry_1, 
        next_reg_H7_cry_2, next_reg_H7_cry_3, next_reg_H7_cry_4, 
        next_reg_H7_cry_5, next_reg_H7_cry_6, next_reg_H7_cry_7, 
        next_reg_H7_cry_8, next_reg_H7_cry_9, next_reg_H7_cry_10, 
        next_reg_H7_cry_11, next_reg_H7_cry_12, 
        next_reg_H7_cry_13, next_reg_H7_cry_14, 
        next_reg_H7_cry_15, next_reg_H7_cry_16, 
        next_reg_H7_cry_17, next_reg_H7_cry_18, 
        next_reg_H7_cry_19, next_reg_H7_cry_20, 
        next_reg_H7_cry_21, next_reg_H7_cry_22, 
        next_reg_H7_cry_23, next_reg_H7_cry_24, 
        next_reg_H7_cry_25, next_reg_H7_cry_26, 
        next_reg_H7_cry_27, next_reg_H7_cry_28, 
        next_reg_H7_cry_29, next_reg_H7_cry_30 : std_logic;

begin 

    SHA256_BLOCK_0_H0_o(31) <= \SHA256_BLOCK_0_H0_o[31]\;
    SHA256_BLOCK_0_H0_o(30) <= \SHA256_BLOCK_0_H0_o[30]\;
    SHA256_BLOCK_0_H0_o(29) <= \SHA256_BLOCK_0_H0_o[29]\;
    SHA256_BLOCK_0_H0_o(28) <= \SHA256_BLOCK_0_H0_o[28]\;
    SHA256_BLOCK_0_H0_o(27) <= \SHA256_BLOCK_0_H0_o[27]\;
    SHA256_BLOCK_0_H0_o(26) <= \SHA256_BLOCK_0_H0_o[26]\;
    SHA256_BLOCK_0_H0_o(25) <= \SHA256_BLOCK_0_H0_o[25]\;
    SHA256_BLOCK_0_H0_o(24) <= \SHA256_BLOCK_0_H0_o[24]\;
    SHA256_BLOCK_0_H0_o(23) <= \SHA256_BLOCK_0_H0_o[23]\;
    SHA256_BLOCK_0_H0_o(22) <= \SHA256_BLOCK_0_H0_o[22]\;
    SHA256_BLOCK_0_H0_o(21) <= \SHA256_BLOCK_0_H0_o[21]\;
    SHA256_BLOCK_0_H0_o(20) <= \SHA256_BLOCK_0_H0_o[20]\;
    SHA256_BLOCK_0_H0_o(19) <= \SHA256_BLOCK_0_H0_o[19]\;
    SHA256_BLOCK_0_H0_o(18) <= \SHA256_BLOCK_0_H0_o[18]\;
    SHA256_BLOCK_0_H0_o(17) <= \SHA256_BLOCK_0_H0_o[17]\;
    SHA256_BLOCK_0_H0_o(16) <= \SHA256_BLOCK_0_H0_o[16]\;
    SHA256_BLOCK_0_H0_o(15) <= \SHA256_BLOCK_0_H0_o[15]\;
    SHA256_BLOCK_0_H0_o(14) <= \SHA256_BLOCK_0_H0_o[14]\;
    SHA256_BLOCK_0_H0_o(13) <= \SHA256_BLOCK_0_H0_o[13]\;
    SHA256_BLOCK_0_H0_o(12) <= \SHA256_BLOCK_0_H0_o[12]\;
    SHA256_BLOCK_0_H0_o(11) <= \SHA256_BLOCK_0_H0_o[11]\;
    SHA256_BLOCK_0_H0_o(10) <= \SHA256_BLOCK_0_H0_o[10]\;
    SHA256_BLOCK_0_H0_o(9) <= \SHA256_BLOCK_0_H0_o[9]\;
    SHA256_BLOCK_0_H0_o(8) <= \SHA256_BLOCK_0_H0_o[8]\;
    SHA256_BLOCK_0_H0_o(7) <= \SHA256_BLOCK_0_H0_o[7]\;
    SHA256_BLOCK_0_H0_o(6) <= \SHA256_BLOCK_0_H0_o[6]\;
    SHA256_BLOCK_0_H0_o(5) <= \SHA256_BLOCK_0_H0_o[5]\;
    SHA256_BLOCK_0_H0_o(4) <= \SHA256_BLOCK_0_H0_o[4]\;
    SHA256_BLOCK_0_H0_o(3) <= \SHA256_BLOCK_0_H0_o[3]\;
    SHA256_BLOCK_0_H0_o(2) <= \SHA256_BLOCK_0_H0_o[2]\;
    SHA256_BLOCK_0_H0_o(1) <= \SHA256_BLOCK_0_H0_o[1]\;
    SHA256_BLOCK_0_H0_o(0) <= \SHA256_BLOCK_0_H0_o[0]\;
    N0_data(31) <= \N0_data[31]\;
    N0_data(30) <= \N0_data[30]\;
    N0_data(29) <= \N0_data[29]\;
    N0_data(28) <= \N0_data[28]\;
    N0_data(27) <= \N0_data[27]\;
    N0_data(26) <= \N0_data[26]\;
    N0_data(25) <= \N0_data[25]\;
    N0_data(24) <= \N0_data[24]\;
    N0_data(23) <= \N0_data[23]\;
    N0_data(22) <= \N0_data[22]\;
    N0_data(21) <= \N0_data[21]\;
    N0_data(20) <= \N0_data[20]\;
    N0_data(19) <= \N0_data[19]\;
    N0_data(18) <= \N0_data[18]\;
    N0_data(17) <= \N0_data[17]\;
    N0_data(16) <= \N0_data[16]\;
    N0_data(15) <= \N0_data[15]\;
    N0_data(14) <= \N0_data[14]\;
    N0_data(13) <= \N0_data[13]\;
    N0_data(12) <= \N0_data[12]\;
    N0_data(11) <= \N0_data[11]\;
    N0_data(10) <= \N0_data[10]\;
    N0_data(9) <= \N0_data[9]\;
    N0_data(8) <= \N0_data[8]\;
    N0_data(7) <= \N0_data[7]\;
    N0_data(6) <= \N0_data[6]\;
    N0_data(5) <= \N0_data[5]\;
    N0_data(4) <= \N0_data[4]\;
    N0_data(3) <= \N0_data[3]\;
    N0_data(2) <= \N0_data[2]\;
    N0_data(1) <= \N0_data[1]\;
    SHA256_BLOCK_0_H1_o(31) <= \SHA256_BLOCK_0_H1_o[31]\;
    SHA256_BLOCK_0_H1_o(30) <= \SHA256_BLOCK_0_H1_o[30]\;
    SHA256_BLOCK_0_H1_o(29) <= \SHA256_BLOCK_0_H1_o[29]\;
    SHA256_BLOCK_0_H1_o(28) <= \SHA256_BLOCK_0_H1_o[28]\;
    SHA256_BLOCK_0_H1_o(27) <= \SHA256_BLOCK_0_H1_o[27]\;
    SHA256_BLOCK_0_H1_o(26) <= \SHA256_BLOCK_0_H1_o[26]\;
    SHA256_BLOCK_0_H1_o(25) <= \SHA256_BLOCK_0_H1_o[25]\;
    SHA256_BLOCK_0_H1_o(24) <= \SHA256_BLOCK_0_H1_o[24]\;
    SHA256_BLOCK_0_H1_o(23) <= \SHA256_BLOCK_0_H1_o[23]\;
    SHA256_BLOCK_0_H1_o(22) <= \SHA256_BLOCK_0_H1_o[22]\;
    SHA256_BLOCK_0_H1_o(21) <= \SHA256_BLOCK_0_H1_o[21]\;
    SHA256_BLOCK_0_H1_o(20) <= \SHA256_BLOCK_0_H1_o[20]\;
    SHA256_BLOCK_0_H1_o(19) <= \SHA256_BLOCK_0_H1_o[19]\;
    SHA256_BLOCK_0_H1_o(18) <= \SHA256_BLOCK_0_H1_o[18]\;
    SHA256_BLOCK_0_H1_o(17) <= \SHA256_BLOCK_0_H1_o[17]\;
    SHA256_BLOCK_0_H1_o(16) <= \SHA256_BLOCK_0_H1_o[16]\;
    SHA256_BLOCK_0_H1_o(15) <= \SHA256_BLOCK_0_H1_o[15]\;
    SHA256_BLOCK_0_H1_o(14) <= \SHA256_BLOCK_0_H1_o[14]\;
    SHA256_BLOCK_0_H1_o(13) <= \SHA256_BLOCK_0_H1_o[13]\;
    SHA256_BLOCK_0_H1_o(12) <= \SHA256_BLOCK_0_H1_o[12]\;
    SHA256_BLOCK_0_H1_o(11) <= \SHA256_BLOCK_0_H1_o[11]\;
    SHA256_BLOCK_0_H1_o(10) <= \SHA256_BLOCK_0_H1_o[10]\;
    SHA256_BLOCK_0_H1_o(9) <= \SHA256_BLOCK_0_H1_o[9]\;
    SHA256_BLOCK_0_H1_o(8) <= \SHA256_BLOCK_0_H1_o[8]\;
    SHA256_BLOCK_0_H1_o(7) <= \SHA256_BLOCK_0_H1_o[7]\;
    SHA256_BLOCK_0_H1_o(6) <= \SHA256_BLOCK_0_H1_o[6]\;
    SHA256_BLOCK_0_H1_o(5) <= \SHA256_BLOCK_0_H1_o[5]\;
    SHA256_BLOCK_0_H1_o(4) <= \SHA256_BLOCK_0_H1_o[4]\;
    SHA256_BLOCK_0_H1_o(3) <= \SHA256_BLOCK_0_H1_o[3]\;
    SHA256_BLOCK_0_H1_o(2) <= \SHA256_BLOCK_0_H1_o[2]\;
    SHA256_BLOCK_0_H1_o(1) <= \SHA256_BLOCK_0_H1_o[1]\;
    SHA256_BLOCK_0_H1_o(0) <= \SHA256_BLOCK_0_H1_o[0]\;
    N1_data(31) <= \N1_data[31]\;
    N1_data(30) <= \N1_data[30]\;
    N1_data(29) <= \N1_data[29]\;
    N1_data(28) <= \N1_data[28]\;
    N1_data(27) <= \N1_data[27]\;
    N1_data(26) <= \N1_data[26]\;
    N1_data(25) <= \N1_data[25]\;
    N1_data(24) <= \N1_data[24]\;
    N1_data(23) <= \N1_data[23]\;
    N1_data(22) <= \N1_data[22]\;
    N1_data(21) <= \N1_data[21]\;
    N1_data(20) <= \N1_data[20]\;
    N1_data(19) <= \N1_data[19]\;
    N1_data(18) <= \N1_data[18]\;
    N1_data(17) <= \N1_data[17]\;
    N1_data(16) <= \N1_data[16]\;
    N1_data(15) <= \N1_data[15]\;
    N1_data(14) <= \N1_data[14]\;
    N1_data(13) <= \N1_data[13]\;
    N1_data(12) <= \N1_data[12]\;
    N1_data(11) <= \N1_data[11]\;
    N1_data(10) <= \N1_data[10]\;
    N1_data(9) <= \N1_data[9]\;
    N1_data(8) <= \N1_data[8]\;
    N1_data(7) <= \N1_data[7]\;
    N1_data(6) <= \N1_data[6]\;
    N1_data(5) <= \N1_data[5]\;
    N1_data(4) <= \N1_data[4]\;
    N1_data(3) <= \N1_data[3]\;
    N1_data(2) <= \N1_data[2]\;
    N1_data(1) <= \N1_data[1]\;
    SHA256_BLOCK_0_H2_o(31) <= \SHA256_BLOCK_0_H2_o[31]\;
    SHA256_BLOCK_0_H2_o(30) <= \SHA256_BLOCK_0_H2_o[30]\;
    SHA256_BLOCK_0_H2_o(29) <= \SHA256_BLOCK_0_H2_o[29]\;
    SHA256_BLOCK_0_H2_o(28) <= \SHA256_BLOCK_0_H2_o[28]\;
    SHA256_BLOCK_0_H2_o(27) <= \SHA256_BLOCK_0_H2_o[27]\;
    SHA256_BLOCK_0_H2_o(26) <= \SHA256_BLOCK_0_H2_o[26]\;
    SHA256_BLOCK_0_H2_o(25) <= \SHA256_BLOCK_0_H2_o[25]\;
    SHA256_BLOCK_0_H2_o(24) <= \SHA256_BLOCK_0_H2_o[24]\;
    SHA256_BLOCK_0_H2_o(23) <= \SHA256_BLOCK_0_H2_o[23]\;
    SHA256_BLOCK_0_H2_o(22) <= \SHA256_BLOCK_0_H2_o[22]\;
    SHA256_BLOCK_0_H2_o(21) <= \SHA256_BLOCK_0_H2_o[21]\;
    SHA256_BLOCK_0_H2_o(20) <= \SHA256_BLOCK_0_H2_o[20]\;
    SHA256_BLOCK_0_H2_o(19) <= \SHA256_BLOCK_0_H2_o[19]\;
    SHA256_BLOCK_0_H2_o(18) <= \SHA256_BLOCK_0_H2_o[18]\;
    SHA256_BLOCK_0_H2_o(17) <= \SHA256_BLOCK_0_H2_o[17]\;
    SHA256_BLOCK_0_H2_o(16) <= \SHA256_BLOCK_0_H2_o[16]\;
    SHA256_BLOCK_0_H2_o(15) <= \SHA256_BLOCK_0_H2_o[15]\;
    SHA256_BLOCK_0_H2_o(14) <= \SHA256_BLOCK_0_H2_o[14]\;
    SHA256_BLOCK_0_H2_o(13) <= \SHA256_BLOCK_0_H2_o[13]\;
    SHA256_BLOCK_0_H2_o(12) <= \SHA256_BLOCK_0_H2_o[12]\;
    SHA256_BLOCK_0_H2_o(11) <= \SHA256_BLOCK_0_H2_o[11]\;
    SHA256_BLOCK_0_H2_o(10) <= \SHA256_BLOCK_0_H2_o[10]\;
    SHA256_BLOCK_0_H2_o(9) <= \SHA256_BLOCK_0_H2_o[9]\;
    SHA256_BLOCK_0_H2_o(8) <= \SHA256_BLOCK_0_H2_o[8]\;
    SHA256_BLOCK_0_H2_o(7) <= \SHA256_BLOCK_0_H2_o[7]\;
    SHA256_BLOCK_0_H2_o(6) <= \SHA256_BLOCK_0_H2_o[6]\;
    SHA256_BLOCK_0_H2_o(5) <= \SHA256_BLOCK_0_H2_o[5]\;
    SHA256_BLOCK_0_H2_o(4) <= \SHA256_BLOCK_0_H2_o[4]\;
    SHA256_BLOCK_0_H2_o(3) <= \SHA256_BLOCK_0_H2_o[3]\;
    SHA256_BLOCK_0_H2_o(2) <= \SHA256_BLOCK_0_H2_o[2]\;
    SHA256_BLOCK_0_H2_o(1) <= \SHA256_BLOCK_0_H2_o[1]\;
    SHA256_BLOCK_0_H2_o(0) <= \SHA256_BLOCK_0_H2_o[0]\;
    N2_data(31) <= \N2_data[31]\;
    N2_data(30) <= \N2_data[30]\;
    N2_data(29) <= \N2_data[29]\;
    N2_data(28) <= \N2_data[28]\;
    N2_data(27) <= \N2_data[27]\;
    N2_data(26) <= \N2_data[26]\;
    N2_data(25) <= \N2_data[25]\;
    N2_data(24) <= \N2_data[24]\;
    N2_data(23) <= \N2_data[23]\;
    N2_data(22) <= \N2_data[22]\;
    N2_data(21) <= \N2_data[21]\;
    N2_data(20) <= \N2_data[20]\;
    N2_data(19) <= \N2_data[19]\;
    N2_data(18) <= \N2_data[18]\;
    N2_data(17) <= \N2_data[17]\;
    N2_data(16) <= \N2_data[16]\;
    N2_data(15) <= \N2_data[15]\;
    N2_data(14) <= \N2_data[14]\;
    N2_data(13) <= \N2_data[13]\;
    N2_data(12) <= \N2_data[12]\;
    N2_data(11) <= \N2_data[11]\;
    N2_data(10) <= \N2_data[10]\;
    N2_data(9) <= \N2_data[9]\;
    N2_data(8) <= \N2_data[8]\;
    N2_data(7) <= \N2_data[7]\;
    N2_data(6) <= \N2_data[6]\;
    N2_data(5) <= \N2_data[5]\;
    N2_data(4) <= \N2_data[4]\;
    N2_data(3) <= \N2_data[3]\;
    N2_data(2) <= \N2_data[2]\;
    N2_data(1) <= \N2_data[1]\;
    SHA256_BLOCK_0_H3_o(31) <= \SHA256_BLOCK_0_H3_o[31]\;
    SHA256_BLOCK_0_H3_o(30) <= \SHA256_BLOCK_0_H3_o[30]\;
    SHA256_BLOCK_0_H3_o(29) <= \SHA256_BLOCK_0_H3_o[29]\;
    SHA256_BLOCK_0_H3_o(28) <= \SHA256_BLOCK_0_H3_o[28]\;
    SHA256_BLOCK_0_H3_o(27) <= \SHA256_BLOCK_0_H3_o[27]\;
    SHA256_BLOCK_0_H3_o(26) <= \SHA256_BLOCK_0_H3_o[26]\;
    SHA256_BLOCK_0_H3_o(25) <= \SHA256_BLOCK_0_H3_o[25]\;
    SHA256_BLOCK_0_H3_o(24) <= \SHA256_BLOCK_0_H3_o[24]\;
    SHA256_BLOCK_0_H3_o(23) <= \SHA256_BLOCK_0_H3_o[23]\;
    SHA256_BLOCK_0_H3_o(22) <= \SHA256_BLOCK_0_H3_o[22]\;
    SHA256_BLOCK_0_H3_o(21) <= \SHA256_BLOCK_0_H3_o[21]\;
    SHA256_BLOCK_0_H3_o(20) <= \SHA256_BLOCK_0_H3_o[20]\;
    SHA256_BLOCK_0_H3_o(19) <= \SHA256_BLOCK_0_H3_o[19]\;
    SHA256_BLOCK_0_H3_o(18) <= \SHA256_BLOCK_0_H3_o[18]\;
    SHA256_BLOCK_0_H3_o(17) <= \SHA256_BLOCK_0_H3_o[17]\;
    SHA256_BLOCK_0_H3_o(16) <= \SHA256_BLOCK_0_H3_o[16]\;
    SHA256_BLOCK_0_H3_o(15) <= \SHA256_BLOCK_0_H3_o[15]\;
    SHA256_BLOCK_0_H3_o(14) <= \SHA256_BLOCK_0_H3_o[14]\;
    SHA256_BLOCK_0_H3_o(13) <= \SHA256_BLOCK_0_H3_o[13]\;
    SHA256_BLOCK_0_H3_o(12) <= \SHA256_BLOCK_0_H3_o[12]\;
    SHA256_BLOCK_0_H3_o(11) <= \SHA256_BLOCK_0_H3_o[11]\;
    SHA256_BLOCK_0_H3_o(10) <= \SHA256_BLOCK_0_H3_o[10]\;
    SHA256_BLOCK_0_H3_o(9) <= \SHA256_BLOCK_0_H3_o[9]\;
    SHA256_BLOCK_0_H3_o(8) <= \SHA256_BLOCK_0_H3_o[8]\;
    SHA256_BLOCK_0_H3_o(7) <= \SHA256_BLOCK_0_H3_o[7]\;
    SHA256_BLOCK_0_H3_o(6) <= \SHA256_BLOCK_0_H3_o[6]\;
    SHA256_BLOCK_0_H3_o(5) <= \SHA256_BLOCK_0_H3_o[5]\;
    SHA256_BLOCK_0_H3_o(4) <= \SHA256_BLOCK_0_H3_o[4]\;
    SHA256_BLOCK_0_H3_o(3) <= \SHA256_BLOCK_0_H3_o[3]\;
    SHA256_BLOCK_0_H3_o(2) <= \SHA256_BLOCK_0_H3_o[2]\;
    SHA256_BLOCK_0_H3_o(1) <= \SHA256_BLOCK_0_H3_o[1]\;
    SHA256_BLOCK_0_H3_o(0) <= \SHA256_BLOCK_0_H3_o[0]\;
    N3_data(31) <= \N3_data[31]\;
    N3_data(30) <= \N3_data[30]\;
    N3_data(29) <= \N3_data[29]\;
    N3_data(28) <= \N3_data[28]\;
    N3_data(27) <= \N3_data[27]\;
    N3_data(26) <= \N3_data[26]\;
    N3_data(25) <= \N3_data[25]\;
    N3_data(24) <= \N3_data[24]\;
    N3_data(23) <= \N3_data[23]\;
    N3_data(22) <= \N3_data[22]\;
    N3_data(21) <= \N3_data[21]\;
    N3_data(20) <= \N3_data[20]\;
    N3_data(19) <= \N3_data[19]\;
    N3_data(18) <= \N3_data[18]\;
    N3_data(17) <= \N3_data[17]\;
    N3_data(16) <= \N3_data[16]\;
    N3_data(15) <= \N3_data[15]\;
    N3_data(14) <= \N3_data[14]\;
    N3_data(13) <= \N3_data[13]\;
    N3_data(12) <= \N3_data[12]\;
    N3_data(11) <= \N3_data[11]\;
    N3_data(10) <= \N3_data[10]\;
    N3_data(9) <= \N3_data[9]\;
    N3_data(8) <= \N3_data[8]\;
    N3_data(7) <= \N3_data[7]\;
    N3_data(6) <= \N3_data[6]\;
    N3_data(5) <= \N3_data[5]\;
    N3_data(4) <= \N3_data[4]\;
    N3_data(3) <= \N3_data[3]\;
    N3_data(2) <= \N3_data[2]\;
    N3_data(1) <= \N3_data[1]\;
    SHA256_BLOCK_0_H4_o(31) <= \SHA256_BLOCK_0_H4_o[31]\;
    SHA256_BLOCK_0_H4_o(30) <= \SHA256_BLOCK_0_H4_o[30]\;
    SHA256_BLOCK_0_H4_o(29) <= \SHA256_BLOCK_0_H4_o[29]\;
    SHA256_BLOCK_0_H4_o(28) <= \SHA256_BLOCK_0_H4_o[28]\;
    SHA256_BLOCK_0_H4_o(27) <= \SHA256_BLOCK_0_H4_o[27]\;
    SHA256_BLOCK_0_H4_o(26) <= \SHA256_BLOCK_0_H4_o[26]\;
    SHA256_BLOCK_0_H4_o(25) <= \SHA256_BLOCK_0_H4_o[25]\;
    SHA256_BLOCK_0_H4_o(24) <= \SHA256_BLOCK_0_H4_o[24]\;
    SHA256_BLOCK_0_H4_o(23) <= \SHA256_BLOCK_0_H4_o[23]\;
    SHA256_BLOCK_0_H4_o(22) <= \SHA256_BLOCK_0_H4_o[22]\;
    SHA256_BLOCK_0_H4_o(21) <= \SHA256_BLOCK_0_H4_o[21]\;
    SHA256_BLOCK_0_H4_o(20) <= \SHA256_BLOCK_0_H4_o[20]\;
    SHA256_BLOCK_0_H4_o(19) <= \SHA256_BLOCK_0_H4_o[19]\;
    SHA256_BLOCK_0_H4_o(18) <= \SHA256_BLOCK_0_H4_o[18]\;
    SHA256_BLOCK_0_H4_o(17) <= \SHA256_BLOCK_0_H4_o[17]\;
    SHA256_BLOCK_0_H4_o(16) <= \SHA256_BLOCK_0_H4_o[16]\;
    SHA256_BLOCK_0_H4_o(15) <= \SHA256_BLOCK_0_H4_o[15]\;
    SHA256_BLOCK_0_H4_o(14) <= \SHA256_BLOCK_0_H4_o[14]\;
    SHA256_BLOCK_0_H4_o(13) <= \SHA256_BLOCK_0_H4_o[13]\;
    SHA256_BLOCK_0_H4_o(12) <= \SHA256_BLOCK_0_H4_o[12]\;
    SHA256_BLOCK_0_H4_o(11) <= \SHA256_BLOCK_0_H4_o[11]\;
    SHA256_BLOCK_0_H4_o(10) <= \SHA256_BLOCK_0_H4_o[10]\;
    SHA256_BLOCK_0_H4_o(9) <= \SHA256_BLOCK_0_H4_o[9]\;
    SHA256_BLOCK_0_H4_o(8) <= \SHA256_BLOCK_0_H4_o[8]\;
    SHA256_BLOCK_0_H4_o(7) <= \SHA256_BLOCK_0_H4_o[7]\;
    SHA256_BLOCK_0_H4_o(6) <= \SHA256_BLOCK_0_H4_o[6]\;
    SHA256_BLOCK_0_H4_o(5) <= \SHA256_BLOCK_0_H4_o[5]\;
    SHA256_BLOCK_0_H4_o(4) <= \SHA256_BLOCK_0_H4_o[4]\;
    SHA256_BLOCK_0_H4_o(3) <= \SHA256_BLOCK_0_H4_o[3]\;
    SHA256_BLOCK_0_H4_o(2) <= \SHA256_BLOCK_0_H4_o[2]\;
    SHA256_BLOCK_0_H4_o(1) <= \SHA256_BLOCK_0_H4_o[1]\;
    SHA256_BLOCK_0_H4_o(0) <= \SHA256_BLOCK_0_H4_o[0]\;
    N4_data(31) <= \N4_data[31]\;
    N4_data(30) <= \N4_data[30]\;
    N4_data(29) <= \N4_data[29]\;
    N4_data(28) <= \N4_data[28]\;
    N4_data(27) <= \N4_data[27]\;
    N4_data(26) <= \N4_data[26]\;
    N4_data(25) <= \N4_data[25]\;
    N4_data(24) <= \N4_data[24]\;
    N4_data(23) <= \N4_data[23]\;
    N4_data(22) <= \N4_data[22]\;
    N4_data(21) <= \N4_data[21]\;
    N4_data(20) <= \N4_data[20]\;
    N4_data(19) <= \N4_data[19]\;
    N4_data(18) <= \N4_data[18]\;
    N4_data(17) <= \N4_data[17]\;
    N4_data(16) <= \N4_data[16]\;
    N4_data(15) <= \N4_data[15]\;
    N4_data(14) <= \N4_data[14]\;
    N4_data(13) <= \N4_data[13]\;
    N4_data(12) <= \N4_data[12]\;
    N4_data(11) <= \N4_data[11]\;
    N4_data(10) <= \N4_data[10]\;
    N4_data(9) <= \N4_data[9]\;
    N4_data(8) <= \N4_data[8]\;
    N4_data(7) <= \N4_data[7]\;
    N4_data(6) <= \N4_data[6]\;
    N4_data(5) <= \N4_data[5]\;
    N4_data(4) <= \N4_data[4]\;
    N4_data(3) <= \N4_data[3]\;
    N4_data(2) <= \N4_data[2]\;
    N4_data(1) <= \N4_data[1]\;
    N5_data(31) <= \N5_data[31]\;
    N5_data(30) <= \N5_data[30]\;
    N5_data(29) <= \N5_data[29]\;
    N5_data(28) <= \N5_data[28]\;
    N5_data(27) <= \N5_data[27]\;
    N5_data(26) <= \N5_data[26]\;
    N5_data(25) <= \N5_data[25]\;
    N5_data(24) <= \N5_data[24]\;
    N5_data(23) <= \N5_data[23]\;
    N5_data(22) <= \N5_data[22]\;
    N5_data(21) <= \N5_data[21]\;
    N5_data(20) <= \N5_data[20]\;
    N5_data(19) <= \N5_data[19]\;
    N5_data(18) <= \N5_data[18]\;
    N5_data(17) <= \N5_data[17]\;
    N5_data(16) <= \N5_data[16]\;
    N5_data(15) <= \N5_data[15]\;
    N5_data(14) <= \N5_data[14]\;
    N5_data(13) <= \N5_data[13]\;
    N5_data(12) <= \N5_data[12]\;
    N5_data(11) <= \N5_data[11]\;
    N5_data(10) <= \N5_data[10]\;
    N5_data(9) <= \N5_data[9]\;
    N5_data(8) <= \N5_data[8]\;
    N5_data(7) <= \N5_data[7]\;
    N5_data(6) <= \N5_data[6]\;
    N5_data(5) <= \N5_data[5]\;
    N5_data(4) <= \N5_data[4]\;
    N5_data(3) <= \N5_data[3]\;
    N5_data(2) <= \N5_data[2]\;
    N5_data(1) <= \N5_data[1]\;
    SHA256_BLOCK_0_H5_o(31) <= \SHA256_BLOCK_0_H5_o[31]\;
    SHA256_BLOCK_0_H5_o(30) <= \SHA256_BLOCK_0_H5_o[30]\;
    SHA256_BLOCK_0_H5_o(29) <= \SHA256_BLOCK_0_H5_o[29]\;
    SHA256_BLOCK_0_H5_o(28) <= \SHA256_BLOCK_0_H5_o[28]\;
    SHA256_BLOCK_0_H5_o(27) <= \SHA256_BLOCK_0_H5_o[27]\;
    SHA256_BLOCK_0_H5_o(26) <= \SHA256_BLOCK_0_H5_o[26]\;
    SHA256_BLOCK_0_H5_o(25) <= \SHA256_BLOCK_0_H5_o[25]\;
    SHA256_BLOCK_0_H5_o(24) <= \SHA256_BLOCK_0_H5_o[24]\;
    SHA256_BLOCK_0_H5_o(23) <= \SHA256_BLOCK_0_H5_o[23]\;
    SHA256_BLOCK_0_H5_o(22) <= \SHA256_BLOCK_0_H5_o[22]\;
    SHA256_BLOCK_0_H5_o(21) <= \SHA256_BLOCK_0_H5_o[21]\;
    SHA256_BLOCK_0_H5_o(20) <= \SHA256_BLOCK_0_H5_o[20]\;
    SHA256_BLOCK_0_H5_o(19) <= \SHA256_BLOCK_0_H5_o[19]\;
    SHA256_BLOCK_0_H5_o(18) <= \SHA256_BLOCK_0_H5_o[18]\;
    SHA256_BLOCK_0_H5_o(17) <= \SHA256_BLOCK_0_H5_o[17]\;
    SHA256_BLOCK_0_H5_o(16) <= \SHA256_BLOCK_0_H5_o[16]\;
    SHA256_BLOCK_0_H5_o(15) <= \SHA256_BLOCK_0_H5_o[15]\;
    SHA256_BLOCK_0_H5_o(14) <= \SHA256_BLOCK_0_H5_o[14]\;
    SHA256_BLOCK_0_H5_o(13) <= \SHA256_BLOCK_0_H5_o[13]\;
    SHA256_BLOCK_0_H5_o(12) <= \SHA256_BLOCK_0_H5_o[12]\;
    SHA256_BLOCK_0_H5_o(11) <= \SHA256_BLOCK_0_H5_o[11]\;
    SHA256_BLOCK_0_H5_o(10) <= \SHA256_BLOCK_0_H5_o[10]\;
    SHA256_BLOCK_0_H5_o(9) <= \SHA256_BLOCK_0_H5_o[9]\;
    SHA256_BLOCK_0_H5_o(8) <= \SHA256_BLOCK_0_H5_o[8]\;
    SHA256_BLOCK_0_H5_o(7) <= \SHA256_BLOCK_0_H5_o[7]\;
    SHA256_BLOCK_0_H5_o(6) <= \SHA256_BLOCK_0_H5_o[6]\;
    SHA256_BLOCK_0_H5_o(5) <= \SHA256_BLOCK_0_H5_o[5]\;
    SHA256_BLOCK_0_H5_o(4) <= \SHA256_BLOCK_0_H5_o[4]\;
    SHA256_BLOCK_0_H5_o(3) <= \SHA256_BLOCK_0_H5_o[3]\;
    SHA256_BLOCK_0_H5_o(2) <= \SHA256_BLOCK_0_H5_o[2]\;
    SHA256_BLOCK_0_H5_o(1) <= \SHA256_BLOCK_0_H5_o[1]\;
    SHA256_BLOCK_0_H5_o(0) <= \SHA256_BLOCK_0_H5_o[0]\;
    SHA256_BLOCK_0_H6_o(31) <= \SHA256_BLOCK_0_H6_o[31]\;
    SHA256_BLOCK_0_H6_o(30) <= \SHA256_BLOCK_0_H6_o[30]\;
    SHA256_BLOCK_0_H6_o(29) <= \SHA256_BLOCK_0_H6_o[29]\;
    SHA256_BLOCK_0_H6_o(28) <= \SHA256_BLOCK_0_H6_o[28]\;
    SHA256_BLOCK_0_H6_o(27) <= \SHA256_BLOCK_0_H6_o[27]\;
    SHA256_BLOCK_0_H6_o(26) <= \SHA256_BLOCK_0_H6_o[26]\;
    SHA256_BLOCK_0_H6_o(25) <= \SHA256_BLOCK_0_H6_o[25]\;
    SHA256_BLOCK_0_H6_o(24) <= \SHA256_BLOCK_0_H6_o[24]\;
    SHA256_BLOCK_0_H6_o(23) <= \SHA256_BLOCK_0_H6_o[23]\;
    SHA256_BLOCK_0_H6_o(22) <= \SHA256_BLOCK_0_H6_o[22]\;
    SHA256_BLOCK_0_H6_o(21) <= \SHA256_BLOCK_0_H6_o[21]\;
    SHA256_BLOCK_0_H6_o(20) <= \SHA256_BLOCK_0_H6_o[20]\;
    SHA256_BLOCK_0_H6_o(19) <= \SHA256_BLOCK_0_H6_o[19]\;
    SHA256_BLOCK_0_H6_o(18) <= \SHA256_BLOCK_0_H6_o[18]\;
    SHA256_BLOCK_0_H6_o(17) <= \SHA256_BLOCK_0_H6_o[17]\;
    SHA256_BLOCK_0_H6_o(16) <= \SHA256_BLOCK_0_H6_o[16]\;
    SHA256_BLOCK_0_H6_o(15) <= \SHA256_BLOCK_0_H6_o[15]\;
    SHA256_BLOCK_0_H6_o(14) <= \SHA256_BLOCK_0_H6_o[14]\;
    SHA256_BLOCK_0_H6_o(13) <= \SHA256_BLOCK_0_H6_o[13]\;
    SHA256_BLOCK_0_H6_o(12) <= \SHA256_BLOCK_0_H6_o[12]\;
    SHA256_BLOCK_0_H6_o(11) <= \SHA256_BLOCK_0_H6_o[11]\;
    SHA256_BLOCK_0_H6_o(10) <= \SHA256_BLOCK_0_H6_o[10]\;
    SHA256_BLOCK_0_H6_o(9) <= \SHA256_BLOCK_0_H6_o[9]\;
    SHA256_BLOCK_0_H6_o(8) <= \SHA256_BLOCK_0_H6_o[8]\;
    SHA256_BLOCK_0_H6_o(7) <= \SHA256_BLOCK_0_H6_o[7]\;
    SHA256_BLOCK_0_H6_o(6) <= \SHA256_BLOCK_0_H6_o[6]\;
    SHA256_BLOCK_0_H6_o(5) <= \SHA256_BLOCK_0_H6_o[5]\;
    SHA256_BLOCK_0_H6_o(4) <= \SHA256_BLOCK_0_H6_o[4]\;
    SHA256_BLOCK_0_H6_o(3) <= \SHA256_BLOCK_0_H6_o[3]\;
    SHA256_BLOCK_0_H6_o(2) <= \SHA256_BLOCK_0_H6_o[2]\;
    SHA256_BLOCK_0_H6_o(1) <= \SHA256_BLOCK_0_H6_o[1]\;
    SHA256_BLOCK_0_H6_o(0) <= \SHA256_BLOCK_0_H6_o[0]\;
    N6_data(31) <= \N6_data[31]\;
    N6_data(30) <= \N6_data[30]\;
    N6_data(29) <= \N6_data[29]\;
    N6_data(28) <= \N6_data[28]\;
    N6_data(27) <= \N6_data[27]\;
    N6_data(26) <= \N6_data[26]\;
    N6_data(25) <= \N6_data[25]\;
    N6_data(24) <= \N6_data[24]\;
    N6_data(23) <= \N6_data[23]\;
    N6_data(22) <= \N6_data[22]\;
    N6_data(21) <= \N6_data[21]\;
    N6_data(20) <= \N6_data[20]\;
    N6_data(19) <= \N6_data[19]\;
    N6_data(18) <= \N6_data[18]\;
    N6_data(17) <= \N6_data[17]\;
    N6_data(16) <= \N6_data[16]\;
    N6_data(15) <= \N6_data[15]\;
    N6_data(14) <= \N6_data[14]\;
    N6_data(13) <= \N6_data[13]\;
    N6_data(12) <= \N6_data[12]\;
    N6_data(11) <= \N6_data[11]\;
    N6_data(10) <= \N6_data[10]\;
    N6_data(9) <= \N6_data[9]\;
    N6_data(8) <= \N6_data[8]\;
    N6_data(7) <= \N6_data[7]\;
    N6_data(6) <= \N6_data[6]\;
    N6_data(5) <= \N6_data[5]\;
    N6_data(4) <= \N6_data[4]\;
    N6_data(3) <= \N6_data[3]\;
    N6_data(2) <= \N6_data[2]\;
    N6_data(1) <= \N6_data[1]\;
    SHA256_BLOCK_0_H7_o(31) <= \SHA256_BLOCK_0_H7_o[31]\;
    SHA256_BLOCK_0_H7_o(30) <= \SHA256_BLOCK_0_H7_o[30]\;
    SHA256_BLOCK_0_H7_o(29) <= \SHA256_BLOCK_0_H7_o[29]\;
    SHA256_BLOCK_0_H7_o(28) <= \SHA256_BLOCK_0_H7_o[28]\;
    SHA256_BLOCK_0_H7_o(27) <= \SHA256_BLOCK_0_H7_o[27]\;
    SHA256_BLOCK_0_H7_o(26) <= \SHA256_BLOCK_0_H7_o[26]\;
    SHA256_BLOCK_0_H7_o(25) <= \SHA256_BLOCK_0_H7_o[25]\;
    SHA256_BLOCK_0_H7_o(24) <= \SHA256_BLOCK_0_H7_o[24]\;
    SHA256_BLOCK_0_H7_o(23) <= \SHA256_BLOCK_0_H7_o[23]\;
    SHA256_BLOCK_0_H7_o(22) <= \SHA256_BLOCK_0_H7_o[22]\;
    SHA256_BLOCK_0_H7_o(21) <= \SHA256_BLOCK_0_H7_o[21]\;
    SHA256_BLOCK_0_H7_o(20) <= \SHA256_BLOCK_0_H7_o[20]\;
    SHA256_BLOCK_0_H7_o(19) <= \SHA256_BLOCK_0_H7_o[19]\;
    SHA256_BLOCK_0_H7_o(18) <= \SHA256_BLOCK_0_H7_o[18]\;
    SHA256_BLOCK_0_H7_o(17) <= \SHA256_BLOCK_0_H7_o[17]\;
    SHA256_BLOCK_0_H7_o(16) <= \SHA256_BLOCK_0_H7_o[16]\;
    SHA256_BLOCK_0_H7_o(15) <= \SHA256_BLOCK_0_H7_o[15]\;
    SHA256_BLOCK_0_H7_o(14) <= \SHA256_BLOCK_0_H7_o[14]\;
    SHA256_BLOCK_0_H7_o(13) <= \SHA256_BLOCK_0_H7_o[13]\;
    SHA256_BLOCK_0_H7_o(12) <= \SHA256_BLOCK_0_H7_o[12]\;
    SHA256_BLOCK_0_H7_o(11) <= \SHA256_BLOCK_0_H7_o[11]\;
    SHA256_BLOCK_0_H7_o(10) <= \SHA256_BLOCK_0_H7_o[10]\;
    SHA256_BLOCK_0_H7_o(9) <= \SHA256_BLOCK_0_H7_o[9]\;
    SHA256_BLOCK_0_H7_o(8) <= \SHA256_BLOCK_0_H7_o[8]\;
    SHA256_BLOCK_0_H7_o(7) <= \SHA256_BLOCK_0_H7_o[7]\;
    SHA256_BLOCK_0_H7_o(6) <= \SHA256_BLOCK_0_H7_o[6]\;
    SHA256_BLOCK_0_H7_o(5) <= \SHA256_BLOCK_0_H7_o[5]\;
    SHA256_BLOCK_0_H7_o(4) <= \SHA256_BLOCK_0_H7_o[4]\;
    SHA256_BLOCK_0_H7_o(3) <= \SHA256_BLOCK_0_H7_o[3]\;
    SHA256_BLOCK_0_H7_o(2) <= \SHA256_BLOCK_0_H7_o[2]\;
    SHA256_BLOCK_0_H7_o(1) <= \SHA256_BLOCK_0_H7_o[1]\;
    SHA256_BLOCK_0_H7_o(0) <= \SHA256_BLOCK_0_H7_o[0]\;
    N7_data(31) <= \N7_data[31]\;
    N7_data(30) <= \N7_data[30]\;
    N7_data(29) <= \N7_data[29]\;
    N7_data(28) <= \N7_data[28]\;
    N7_data(27) <= \N7_data[27]\;
    N7_data(26) <= \N7_data[26]\;
    N7_data(25) <= \N7_data[25]\;
    N7_data(24) <= \N7_data[24]\;
    N7_data(23) <= \N7_data[23]\;
    N7_data(22) <= \N7_data[22]\;
    N7_data(21) <= \N7_data[21]\;
    N7_data(20) <= \N7_data[20]\;
    N7_data(19) <= \N7_data[19]\;
    N7_data(18) <= \N7_data[18]\;
    N7_data(17) <= \N7_data[17]\;
    N7_data(16) <= \N7_data[16]\;
    N7_data(15) <= \N7_data[15]\;
    N7_data(14) <= \N7_data[14]\;
    N7_data(13) <= \N7_data[13]\;
    N7_data(12) <= \N7_data[12]\;
    N7_data(11) <= \N7_data[11]\;
    N7_data(10) <= \N7_data[10]\;
    N7_data(9) <= \N7_data[9]\;
    N7_data(8) <= \N7_data[8]\;
    N7_data(7) <= \N7_data[7]\;
    N7_data(6) <= \N7_data[6]\;
    N7_data(5) <= \N7_data[5]\;
    N7_data(4) <= \N7_data[4]\;
    N7_data(3) <= \N7_data[3]\;
    N7_data(2) <= \N7_data[2]\;
    N7_data(1) <= \N7_data[1]\;
    next_reg_H0_cry_0_0_Y <= \next_reg_H0_cry_0_0_Y\;
    next_reg_H1_cry_0_0_Y <= \next_reg_H1_cry_0_0_Y\;
    next_reg_H2_cry_0_0_Y <= \next_reg_H2_cry_0_0_Y\;
    next_reg_H3_cry_0_0_Y <= \next_reg_H3_cry_0_0_Y\;
    next_reg_H4_cry_0_0_Y <= \next_reg_H4_cry_0_0_Y\;
    next_reg_H5_cry_0_0_Y <= \next_reg_H5_cry_0_0_Y\;
    next_reg_H6_cry_0_0_Y <= \next_reg_H6_cry_0_0_Y\;
    next_reg_H7_cry_0_0_Y <= \next_reg_H7_cry_0_0_Y\;

    \reg_H7[31]\ : SLE
      port map(D => \N7_data[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[31]\);
    
    next_reg_H2_cry_21_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[21]\, B => 
        hash_control_st_reg_i(6), C => R2_data(21), D => 
        GND_net_1, FCI => next_reg_H2_cry_20, S => \N2_data[21]\, 
        Y => OPEN, FCO => next_reg_H2_cry_21);
    
    \reg_H4[12]\ : SLE
      port map(D => \N4_data[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[12]\);
    
    next_reg_H1_cry_8_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[8]\, B => 
        hash_control_st_reg_i(6), C => R1_data(8), D => GND_net_1, 
        FCI => next_reg_H1_cry_7, S => \N1_data[8]\, Y => OPEN, 
        FCO => next_reg_H1_cry_8);
    
    \reg_H3[4]\ : SLE
      port map(D => \N3_data[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[4]\);
    
    next_reg_H7_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[14]\, B => 
        hash_control_st_reg_i(6), C => R7_data(14), D => 
        GND_net_1, FCI => next_reg_H7_cry_13, S => \N7_data[14]\, 
        Y => OPEN, FCO => next_reg_H7_cry_14);
    
    \reg_H4[17]\ : SLE
      port map(D => \N4_data[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[17]\);
    
    next_reg_H4_cry_22_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[22]\, B => 
        hash_control_st_reg_i(6), C => R4_data(22), D => 
        GND_net_1, FCI => next_reg_H4_cry_21, S => \N4_data[22]\, 
        Y => OPEN, FCO => next_reg_H4_cry_22);
    
    \reg_H1[2]\ : SLE
      port map(D => \N1_data[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[2]\);
    
    next_reg_H7_cry_25_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[25]\, B => 
        hash_control_st_reg_i(6), C => R7_data(25), D => 
        GND_net_1, FCI => next_reg_H7_cry_24, S => \N7_data[25]\, 
        Y => OPEN, FCO => next_reg_H7_cry_25);
    
    next_reg_H4_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[20]\, B => 
        hash_control_st_reg_i(6), C => R4_data(20), D => 
        GND_net_1, FCI => next_reg_H4_cry_19, S => \N4_data[20]\, 
        Y => OPEN, FCO => next_reg_H4_cry_20);
    
    \reg_H6[5]\ : SLE
      port map(D => \N6_data[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[5]\);
    
    next_reg_H0_cry_11_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[11]\, B => 
        hash_control_st_reg_i(6), C => R0_data(11), D => 
        GND_net_1, FCI => next_reg_H0_cry_10, S => \N0_data[11]\, 
        Y => OPEN, FCO => next_reg_H0_cry_11);
    
    \reg_H1[5]\ : SLE
      port map(D => \N1_data[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[5]\);
    
    next_reg_H5_cry_25_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[25]\, B => 
        hash_control_st_reg_i(6), C => R5_data(25), D => 
        GND_net_1, FCI => next_reg_H5_cry_24, S => \N5_data[25]\, 
        Y => OPEN, FCO => next_reg_H5_cry_25);
    
    \reg_H5[12]\ : SLE
      port map(D => \N5_data[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[12]\);
    
    \reg_H3[20]\ : SLE
      port map(D => \N3_data[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[20]\);
    
    next_reg_H5_s_31 : ARI1
      generic map(INIT => x"47D00")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R5_data(31), D => \SHA256_BLOCK_0_H5_o[31]\, FCI => 
        next_reg_H5_cry_30, S => \N5_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    \reg_H0[16]\ : SLE
      port map(D => \N0_data[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[16]\);
    
    next_reg_H3_cry_11_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[11]\, B => 
        hash_control_st_reg_i(6), C => R3_data(11), D => 
        GND_net_1, FCI => next_reg_H3_cry_10, S => \N3_data[11]\, 
        Y => OPEN, FCO => next_reg_H3_cry_11);
    
    \reg_H5[17]\ : SLE
      port map(D => \N5_data[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[17]\);
    
    next_reg_H5_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[14]\, B => 
        hash_control_st_reg_i(6), C => R5_data(14), D => 
        GND_net_1, FCI => next_reg_H5_cry_13, S => \N5_data[14]\, 
        Y => OPEN, FCO => next_reg_H5_cry_14);
    
    next_reg_H1_cry_13_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[13]\, B => 
        hash_control_st_reg_i(6), C => R1_data(13), D => 
        GND_net_1, FCI => next_reg_H1_cry_12, S => \N1_data[13]\, 
        Y => OPEN, FCO => next_reg_H1_cry_13);
    
    \reg_H3[30]\ : SLE
      port map(D => \N3_data[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[30]\);
    
    next_reg_H3_cry_29_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[29]\, B => 
        hash_control_st_reg_i(6), C => R3_data(29), D => 
        GND_net_1, FCI => next_reg_H3_cry_28, S => \N3_data[29]\, 
        Y => OPEN, FCO => next_reg_H3_cry_29);
    
    \reg_H1[8]\ : SLE
      port map(D => \N1_data[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[8]\);
    
    next_reg_H7_cry_4_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[4]\, B => 
        hash_control_st_reg_i(6), C => R7_data(4), D => GND_net_1, 
        FCI => next_reg_H7_cry_3, S => \N7_data[4]\, Y => OPEN, 
        FCO => next_reg_H7_cry_4);
    
    \reg_H5[22]\ : SLE
      port map(D => \N5_data[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[22]\);
    
    next_reg_H6_cry_18_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[18]\, B => 
        hash_control_st_reg_i(6), C => R6_data(18), D => 
        GND_net_1, FCI => next_reg_H6_cry_17, S => \N6_data[18]\, 
        Y => OPEN, FCO => next_reg_H6_cry_18);
    
    \reg_H1[4]\ : SLE
      port map(D => \N1_data[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[4]\);
    
    \reg_H1[21]\ : SLE
      port map(D => \N1_data[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[21]\);
    
    next_reg_H5_cry_9_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[9]\, B => 
        hash_control_st_reg_i(6), C => R5_data(9), D => GND_net_1, 
        FCI => next_reg_H5_cry_8, S => \N5_data[9]\, Y => OPEN, 
        FCO => next_reg_H5_cry_9);
    
    next_reg_H2_cry_0_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[0]\, B => 
        hash_control_st_reg_i(6), C => R2_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H2_cry_0_0_Y\, 
        FCO => next_reg_H2_cry_0);
    
    next_reg_H6_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[24]\, B => 
        hash_control_st_reg_i(6), C => R6_data(24), D => 
        GND_net_1, FCI => next_reg_H6_cry_23, S => \N6_data[24]\, 
        Y => OPEN, FCO => next_reg_H6_cry_24);
    
    \reg_H7[28]\ : SLE
      port map(D => \N7_data[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[28]\);
    
    \reg_H5[31]\ : SLE
      port map(D => \N5_data[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[31]\);
    
    \reg_H5[27]\ : SLE
      port map(D => \N5_data[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[27]\);
    
    next_reg_H7_cry_30_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[30]\, B => 
        hash_control_st_reg_i(6), C => R7_data(30), D => 
        GND_net_1, FCI => next_reg_H7_cry_29, S => \N7_data[30]\, 
        Y => OPEN, FCO => next_reg_H7_cry_30);
    
    \reg_H7[0]\ : SLE
      port map(D => \next_reg_H7_cry_0_0_Y\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[0]\);
    
    \reg_H6[20]\ : SLE
      port map(D => \N6_data[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[20]\);
    
    next_reg_H2_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[15]\, B => 
        hash_control_st_reg_i(6), C => R2_data(15), D => 
        GND_net_1, FCI => next_reg_H2_cry_14, S => \N2_data[15]\, 
        Y => OPEN, FCO => next_reg_H2_cry_15);
    
    \reg_H6[6]\ : SLE
      port map(D => \N6_data[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[6]\);
    
    next_reg_H6_cry_4_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[4]\, B => 
        hash_control_st_reg_i(6), C => R6_data(4), D => GND_net_1, 
        FCI => next_reg_H6_cry_3, S => \N6_data[4]\, Y => OPEN, 
        FCO => next_reg_H6_cry_4);
    
    \reg_H4[7]\ : SLE
      port map(D => \N4_data[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[7]\);
    
    \reg_H4[13]\ : SLE
      port map(D => \N4_data[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[13]\);
    
    next_reg_H4_cry_13_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[13]\, B => 
        hash_control_st_reg_i(6), C => R4_data(13), D => 
        GND_net_1, FCI => next_reg_H4_cry_12, S => \N4_data[13]\, 
        Y => OPEN, FCO => next_reg_H4_cry_13);
    
    next_reg_H0_cry_9_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[9]\, B => 
        hash_control_st_reg_i(6), C => R0_data(9), D => GND_net_1, 
        FCI => next_reg_H0_cry_8, S => \N0_data[9]\, Y => OPEN, 
        FCO => next_reg_H0_cry_9);
    
    \reg_H4[14]\ : SLE
      port map(D => \N4_data[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[14]\);
    
    \reg_H2[9]\ : SLE
      port map(D => \N2_data[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[9]\);
    
    next_reg_H1_cry_25_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[25]\, B => 
        hash_control_st_reg_i(6), C => R1_data(25), D => 
        GND_net_1, FCI => next_reg_H1_cry_24, S => \N1_data[25]\, 
        Y => OPEN, FCO => next_reg_H1_cry_25);
    
    \reg_H2[22]\ : SLE
      port map(D => \N2_data[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[22]\);
    
    \reg_H3[29]\ : SLE
      port map(D => \N3_data[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[29]\);
    
    \reg_H7[25]\ : SLE
      port map(D => \N7_data[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[25]\);
    
    \reg_H0[20]\ : SLE
      port map(D => \N0_data[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[20]\);
    
    \reg_H4[4]\ : SLE
      port map(D => \N4_data[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[4]\);
    
    \reg_H2[27]\ : SLE
      port map(D => \N2_data[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[27]\);
    
    next_reg_H6_cry_30_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[30]\, B => 
        hash_control_st_reg_i(6), C => R6_data(30), D => 
        GND_net_1, FCI => next_reg_H6_cry_29, S => \N6_data[30]\, 
        Y => OPEN, FCO => next_reg_H6_cry_30);
    
    \reg_H1[26]\ : SLE
      port map(D => \N1_data[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[26]\);
    
    next_reg_H7_cry_2_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[2]\, B => 
        hash_control_st_reg_i(6), C => R7_data(2), D => GND_net_1, 
        FCI => next_reg_H7_cry_1, S => \N7_data[2]\, Y => OPEN, 
        FCO => next_reg_H7_cry_2);
    
    next_reg_H3_cry_2_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[2]\, B => 
        hash_control_st_reg_i(6), C => R3_data(2), D => GND_net_1, 
        FCI => next_reg_H3_cry_1, S => \N3_data[2]\, Y => OPEN, 
        FCO => next_reg_H3_cry_2);
    
    next_reg_H0_cry_6_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[6]\, B => 
        hash_control_st_reg_i(6), C => R0_data(6), D => GND_net_1, 
        FCI => next_reg_H0_cry_5, S => \N0_data[6]\, Y => OPEN, 
        FCO => next_reg_H0_cry_6);
    
    next_reg_H7_cry_18_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[18]\, B => 
        hash_control_st_reg_i(6), C => R7_data(18), D => 
        GND_net_1, FCI => next_reg_H7_cry_17, S => \N7_data[18]\, 
        Y => OPEN, FCO => next_reg_H7_cry_18);
    
    next_reg_H6_cry_11_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[11]\, B => 
        hash_control_st_reg_i(6), C => R6_data(11), D => 
        GND_net_1, FCI => next_reg_H6_cry_10, S => \N6_data[11]\, 
        Y => OPEN, FCO => next_reg_H6_cry_11);
    
    next_reg_H3_cry_9_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[9]\, B => 
        hash_control_st_reg_i(6), C => R3_data(9), D => GND_net_1, 
        FCI => next_reg_H3_cry_8, S => \N3_data[9]\, Y => OPEN, 
        FCO => next_reg_H3_cry_9);
    
    \reg_H5[13]\ : SLE
      port map(D => \N5_data[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[13]\);
    
    \reg_H0[1]\ : SLE
      port map(D => \N0_data[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[1]\);
    
    \reg_H5[14]\ : SLE
      port map(D => \N5_data[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[14]\);
    
    \reg_H4[2]\ : SLE
      port map(D => \N4_data[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[2]\);
    
    next_reg_H2_cry_25_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[25]\, B => 
        hash_control_st_reg_i(6), C => R2_data(25), D => 
        GND_net_1, FCI => next_reg_H2_cry_24, S => \N2_data[25]\, 
        Y => OPEN, FCO => next_reg_H2_cry_25);
    
    \reg_H3[8]\ : SLE
      port map(D => \N3_data[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[8]\);
    
    \reg_H6[29]\ : SLE
      port map(D => \N6_data[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[29]\);
    
    \reg_H5[23]\ : SLE
      port map(D => \N5_data[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[23]\);
    
    \reg_H0[12]\ : SLE
      port map(D => \N0_data[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[12]\);
    
    \reg_H5[24]\ : SLE
      port map(D => \N5_data[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[24]\);
    
    next_reg_H5_cry_2_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[2]\, B => 
        hash_control_st_reg_i(6), C => R5_data(2), D => GND_net_1, 
        FCI => next_reg_H5_cry_1, S => \N5_data[2]\, Y => OPEN, 
        FCO => next_reg_H5_cry_2);
    
    next_reg_H0_cry_26_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[26]\, B => 
        hash_control_st_reg_i(6), C => R0_data(26), D => 
        GND_net_1, FCI => next_reg_H0_cry_25, S => \N0_data[26]\, 
        Y => OPEN, FCO => next_reg_H0_cry_26);
    
    next_reg_H0_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[15]\, B => 
        hash_control_st_reg_i(6), C => R0_data(15), D => 
        GND_net_1, FCI => next_reg_H0_cry_14, S => \N0_data[15]\, 
        Y => OPEN, FCO => next_reg_H0_cry_15);
    
    \reg_H7[18]\ : SLE
      port map(D => \N7_data[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[18]\);
    
    \reg_H0[17]\ : SLE
      port map(D => \N0_data[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[17]\);
    
    next_reg_H1_cry_30_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[30]\, B => 
        hash_control_st_reg_i(6), C => R1_data(30), D => 
        GND_net_1, FCI => next_reg_H1_cry_29, S => \N1_data[30]\, 
        Y => OPEN, FCO => next_reg_H1_cry_30);
    
    next_reg_H1_cry_17_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[17]\, B => 
        hash_control_st_reg_i(6), C => R1_data(17), D => 
        GND_net_1, FCI => next_reg_H1_cry_16, S => \N1_data[17]\, 
        Y => OPEN, FCO => next_reg_H1_cry_17);
    
    \reg_H1[1]\ : SLE
      port map(D => \N1_data[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[1]\);
    
    \reg_H1[18]\ : SLE
      port map(D => \N1_data[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[18]\);
    
    next_reg_H5_cry_18_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[18]\, B => 
        hash_control_st_reg_i(6), C => R5_data(18), D => 
        GND_net_1, FCI => next_reg_H5_cry_17, S => \N5_data[18]\, 
        Y => OPEN, FCO => next_reg_H5_cry_18);
    
    next_reg_H3_cry_22_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[22]\, B => 
        hash_control_st_reg_i(6), C => R3_data(22), D => 
        GND_net_1, FCI => next_reg_H3_cry_21, S => \N3_data[22]\, 
        Y => OPEN, FCO => next_reg_H3_cry_22);
    
    next_reg_H7_cry_3_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[3]\, B => 
        hash_control_st_reg_i(6), C => R7_data(3), D => GND_net_1, 
        FCI => next_reg_H7_cry_2, S => \N7_data[3]\, Y => OPEN, 
        FCO => next_reg_H7_cry_3);
    
    next_reg_H3_cry_8_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[8]\, B => 
        hash_control_st_reg_i(6), C => R3_data(8), D => GND_net_1, 
        FCI => next_reg_H3_cry_7, S => \N3_data[8]\, Y => OPEN, 
        FCO => next_reg_H3_cry_8);
    
    next_reg_H3_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[15]\, B => 
        hash_control_st_reg_i(6), C => R3_data(15), D => 
        GND_net_1, FCI => next_reg_H3_cry_14, S => \N3_data[15]\, 
        Y => OPEN, FCO => next_reg_H3_cry_15);
    
    \reg_H0[29]\ : SLE
      port map(D => \N0_data[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[29]\);
    
    next_reg_H4_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[23]\, B => 
        hash_control_st_reg_i(6), C => R4_data(23), D => 
        GND_net_1, FCI => next_reg_H4_cry_22, S => \N4_data[23]\, 
        Y => OPEN, FCO => next_reg_H4_cry_23);
    
    next_reg_H3_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[20]\, B => 
        hash_control_st_reg_i(6), C => R3_data(20), D => 
        GND_net_1, FCI => next_reg_H3_cry_19, S => \N3_data[20]\, 
        Y => OPEN, FCO => next_reg_H3_cry_20);
    
    next_reg_H7_cry_11_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[11]\, B => 
        hash_control_st_reg_i(6), C => R7_data(11), D => 
        GND_net_1, FCI => next_reg_H7_cry_10, S => \N7_data[11]\, 
        Y => OPEN, FCO => next_reg_H7_cry_11);
    
    next_reg_H6_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[28]\, B => 
        hash_control_st_reg_i(6), C => R6_data(28), D => 
        GND_net_1, FCI => next_reg_H6_cry_27, S => \N6_data[28]\, 
        Y => OPEN, FCO => next_reg_H6_cry_28);
    
    \reg_H4[30]\ : SLE
      port map(D => \N4_data[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[30]\);
    
    next_reg_H6_cry_7_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[7]\, B => 
        hash_control_st_reg_i(6), C => R6_data(7), D => GND_net_1, 
        FCI => next_reg_H6_cry_6, S => \N6_data[7]\, Y => OPEN, 
        FCO => next_reg_H6_cry_7);
    
    \reg_H2[23]\ : SLE
      port map(D => \N2_data[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[23]\);
    
    next_reg_H7_cry_26_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[26]\, B => 
        hash_control_st_reg_i(6), C => R7_data(26), D => 
        GND_net_1, FCI => next_reg_H7_cry_25, S => \N7_data[26]\, 
        Y => OPEN, FCO => next_reg_H7_cry_26);
    
    \reg_H2[24]\ : SLE
      port map(D => \N2_data[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[24]\);
    
    \reg_H7[21]\ : SLE
      port map(D => \N7_data[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[21]\);
    
    next_reg_H5_cry_26_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[26]\, B => 
        hash_control_st_reg_i(6), C => R5_data(26), D => 
        GND_net_1, FCI => next_reg_H5_cry_25, S => \N5_data[26]\, 
        Y => OPEN, FCO => next_reg_H5_cry_26);
    
    \reg_H7[15]\ : SLE
      port map(D => \N7_data[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[15]\);
    
    next_reg_H4_cry_17_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[17]\, B => 
        hash_control_st_reg_i(6), C => R4_data(17), D => 
        GND_net_1, FCI => next_reg_H4_cry_16, S => \N4_data[17]\, 
        Y => OPEN, FCO => next_reg_H4_cry_17);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \reg_H5[9]\ : SLE
      port map(D => \N5_data[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[9]\);
    
    \reg_H1[15]\ : SLE
      port map(D => \N1_data[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[15]\);
    
    \reg_H6[9]\ : SLE
      port map(D => \N6_data[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[9]\);
    
    \reg_H6[8]\ : SLE
      port map(D => \N6_data[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[8]\);
    
    \reg_H5[0]\ : SLE
      port map(D => \next_reg_H5_cry_0_0_Y\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[0]\);
    
    \reg_H3[3]\ : SLE
      port map(D => \N3_data[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[3]\);
    
    \reg_H2[18]\ : SLE
      port map(D => \N2_data[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[18]\);
    
    \reg_H1[22]\ : SLE
      port map(D => \N1_data[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[22]\);
    
    \reg_H6[2]\ : SLE
      port map(D => \N6_data[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[2]\);
    
    \reg_H6[18]\ : SLE
      port map(D => \N6_data[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[18]\);
    
    next_reg_H5_cry_3_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[3]\, B => 
        hash_control_st_reg_i(6), C => R5_data(3), D => GND_net_1, 
        FCI => next_reg_H5_cry_2, S => \N5_data[3]\, Y => OPEN, 
        FCO => next_reg_H5_cry_3);
    
    next_reg_H0_cry_29_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[29]\, B => 
        hash_control_st_reg_i(6), C => R0_data(29), D => 
        GND_net_1, FCI => next_reg_H0_cry_28, S => \N0_data[29]\, 
        Y => OPEN, FCO => next_reg_H0_cry_29);
    
    \reg_H0[2]\ : SLE
      port map(D => \N0_data[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[2]\);
    
    next_reg_H5_cry_11_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[11]\, B => 
        hash_control_st_reg_i(6), C => R5_data(11), D => 
        GND_net_1, FCI => next_reg_H5_cry_10, S => \N5_data[11]\, 
        Y => OPEN, FCO => next_reg_H5_cry_11);
    
    \reg_H3[0]\ : SLE
      port map(D => \next_reg_H3_cry_0_0_Y\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[0]\);
    
    \reg_H1[27]\ : SLE
      port map(D => \N1_data[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[27]\);
    
    next_reg_H0_cry_30_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[30]\, B => 
        hash_control_st_reg_i(6), C => R0_data(30), D => 
        GND_net_1, FCI => next_reg_H0_cry_29, S => \N0_data[30]\, 
        Y => OPEN, FCO => next_reg_H0_cry_30);
    
    \reg_H4[28]\ : SLE
      port map(D => \N4_data[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[28]\);
    
    next_reg_H1_cry_14_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[14]\, B => 
        hash_control_st_reg_i(6), C => R1_data(14), D => 
        GND_net_1, FCI => next_reg_H1_cry_13, S => \N1_data[14]\, 
        Y => OPEN, FCO => next_reg_H1_cry_14);
    
    \reg_H0[13]\ : SLE
      port map(D => \N0_data[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[13]\);
    
    \reg_H0[14]\ : SLE
      port map(D => \N0_data[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[14]\);
    
    next_reg_H2_cry_2_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[2]\, B => 
        hash_control_st_reg_i(6), C => R2_data(2), D => GND_net_1, 
        FCI => next_reg_H2_cry_1, S => \N2_data[2]\, Y => OPEN, 
        FCO => next_reg_H2_cry_2);
    
    \reg_H7[26]\ : SLE
      port map(D => \N7_data[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[26]\);
    
    next_reg_H6_cry_21_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[21]\, B => 
        hash_control_st_reg_i(6), C => R6_data(21), D => 
        GND_net_1, FCI => next_reg_H6_cry_20, S => \N6_data[21]\, 
        Y => OPEN, FCO => next_reg_H6_cry_21);
    
    next_reg_H2_cry_16_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[16]\, B => 
        hash_control_st_reg_i(6), C => R2_data(16), D => 
        GND_net_1, FCI => next_reg_H2_cry_15, S => \N2_data[16]\, 
        Y => OPEN, FCO => next_reg_H2_cry_16);
    
    next_reg_H6_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[15]\, B => 
        hash_control_st_reg_i(6), C => R6_data(15), D => 
        GND_net_1, FCI => next_reg_H6_cry_14, S => \N6_data[15]\, 
        Y => OPEN, FCO => next_reg_H6_cry_15);
    
    \reg_H4[10]\ : SLE
      port map(D => \N4_data[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[10]\);
    
    \reg_H0[8]\ : SLE
      port map(D => \N0_data[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[8]\);
    
    \reg_H7[4]\ : SLE
      port map(D => \N7_data[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[4]\);
    
    \reg_H2[15]\ : SLE
      port map(D => \N2_data[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[15]\);
    
    \reg_H6[15]\ : SLE
      port map(D => \N6_data[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[15]\);
    
    next_reg_H7_cry_29_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[29]\, B => 
        hash_control_st_reg_i(6), C => R7_data(29), D => 
        GND_net_1, FCI => next_reg_H7_cry_28, S => \N7_data[29]\, 
        Y => OPEN, FCO => next_reg_H7_cry_29);
    
    next_reg_H1_cry_26_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[26]\, B => 
        hash_control_st_reg_i(6), C => R1_data(26), D => 
        GND_net_1, FCI => next_reg_H1_cry_25, S => \N1_data[26]\, 
        Y => OPEN, FCO => next_reg_H1_cry_26);
    
    next_reg_H5_cry_29_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[29]\, B => 
        hash_control_st_reg_i(6), C => R5_data(29), D => 
        GND_net_1, FCI => next_reg_H5_cry_28, S => \N5_data[29]\, 
        Y => OPEN, FCO => next_reg_H5_cry_29);
    
    next_reg_H1_s_31 : ARI1
      generic map(INIT => x"47D00")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R1_data(31), D => \SHA256_BLOCK_0_H1_o[31]\, FCI => 
        next_reg_H1_cry_30, S => \N1_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    \reg_H4[25]\ : SLE
      port map(D => \N4_data[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[25]\);
    
    next_reg_H4_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[14]\, B => 
        hash_control_st_reg_i(6), C => R4_data(14), D => 
        GND_net_1, FCI => next_reg_H4_cry_13, S => \N4_data[14]\, 
        Y => OPEN, FCO => next_reg_H4_cry_14);
    
    next_reg_H0_cry_5_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[5]\, B => 
        hash_control_st_reg_i(6), C => R0_data(5), D => GND_net_1, 
        FCI => next_reg_H0_cry_4, S => \N0_data[5]\, Y => OPEN, 
        FCO => next_reg_H0_cry_5);
    
    next_reg_H2_cry_5_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[5]\, B => 
        hash_control_st_reg_i(6), C => R2_data(5), D => GND_net_1, 
        FCI => next_reg_H2_cry_4, S => \N2_data[5]\, Y => OPEN, 
        FCO => next_reg_H2_cry_5);
    
    \reg_H2[0]\ : SLE
      port map(D => \next_reg_H2_cry_0_0_Y\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[0]\);
    
    \reg_H7[11]\ : SLE
      port map(D => \N7_data[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[11]\);
    
    next_reg_H6_cry_8_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[8]\, B => 
        hash_control_st_reg_i(6), C => R6_data(8), D => GND_net_1, 
        FCI => next_reg_H6_cry_7, S => \N6_data[8]\, Y => OPEN, 
        FCO => next_reg_H6_cry_8);
    
    next_reg_H4_cry_27_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[27]\, B => 
        hash_control_st_reg_i(6), C => R4_data(27), D => 
        GND_net_1, FCI => next_reg_H4_cry_26, S => \N4_data[27]\, 
        Y => OPEN, FCO => next_reg_H4_cry_27);
    
    \reg_H4[0]\ : SLE
      port map(D => \next_reg_H4_cry_0_0_Y\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[0]\);
    
    \reg_H1[11]\ : SLE
      port map(D => \N1_data[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[11]\);
    
    \reg_H6[31]\ : SLE
      port map(D => \N6_data[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[31]\);
    
    \reg_H5[10]\ : SLE
      port map(D => \N5_data[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[10]\);
    
    \reg_H6[1]\ : SLE
      port map(D => \N6_data[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[1]\);
    
    \reg_H2[30]\ : SLE
      port map(D => \N2_data[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[30]\);
    
    next_reg_H6_cry_2_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[2]\, B => 
        hash_control_st_reg_i(6), C => R6_data(2), D => GND_net_1, 
        FCI => next_reg_H6_cry_1, S => \N6_data[2]\, Y => OPEN, 
        FCO => next_reg_H6_cry_2);
    
    next_reg_H2_cry_26_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[26]\, B => 
        hash_control_st_reg_i(6), C => R2_data(26), D => 
        GND_net_1, FCI => next_reg_H2_cry_25, S => \N2_data[26]\, 
        Y => OPEN, FCO => next_reg_H2_cry_26);
    
    \reg_H7[7]\ : SLE
      port map(D => \N7_data[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[7]\);
    
    \reg_H0[31]\ : SLE
      port map(D => \N0_data[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[31]\);
    
    \reg_H1[23]\ : SLE
      port map(D => \N1_data[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[23]\);
    
    \reg_H1[24]\ : SLE
      port map(D => \N1_data[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[24]\);
    
    next_reg_H7_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[15]\, B => 
        hash_control_st_reg_i(6), C => R7_data(15), D => 
        GND_net_1, FCI => next_reg_H7_cry_14, S => \N7_data[15]\, 
        Y => OPEN, FCO => next_reg_H7_cry_15);
    
    \reg_H5[20]\ : SLE
      port map(D => \N5_data[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[20]\);
    
    \reg_H4[8]\ : SLE
      port map(D => \N4_data[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[8]\);
    
    next_reg_H2_cry_19_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[19]\, B => 
        hash_control_st_reg_i(6), C => R2_data(19), D => 
        GND_net_1, FCI => next_reg_H2_cry_18, S => \N2_data[19]\, 
        Y => OPEN, FCO => next_reg_H2_cry_19);
    
    \reg_H7[5]\ : SLE
      port map(D => \N7_data[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[5]\);
    
    next_reg_H0_cry_16_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[16]\, B => 
        hash_control_st_reg_i(6), C => R0_data(16), D => 
        GND_net_1, FCI => next_reg_H0_cry_15, S => \N0_data[16]\, 
        Y => OPEN, FCO => next_reg_H0_cry_16);
    
    \reg_H4[19]\ : SLE
      port map(D => \N4_data[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[19]\);
    
    \reg_H0[4]\ : SLE
      port map(D => \N0_data[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[4]\);
    
    next_reg_H5_cry_0_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[0]\, B => 
        hash_control_st_reg_i(6), C => R5_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H5_cry_0_0_Y\, 
        FCO => next_reg_H5_cry_0);
    
    next_reg_H1_cry_6_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[6]\, B => 
        hash_control_st_reg_i(6), C => R1_data(6), D => GND_net_1, 
        FCI => next_reg_H1_cry_5, S => \N1_data[6]\, Y => OPEN, 
        FCO => next_reg_H1_cry_6);
    
    next_reg_H1_cry_1_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[1]\, B => 
        hash_control_st_reg_i(6), C => R1_data(1), D => GND_net_1, 
        FCI => next_reg_H1_cry_0, S => \N1_data[1]\, Y => OPEN, 
        FCO => next_reg_H1_cry_1);
    
    \reg_H7[16]\ : SLE
      port map(D => \N7_data[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[16]\);
    
    next_reg_H3_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[23]\, B => 
        hash_control_st_reg_i(6), C => R3_data(23), D => 
        GND_net_1, FCI => next_reg_H3_cry_22, S => \N3_data[23]\, 
        Y => OPEN, FCO => next_reg_H3_cry_23);
    
    \reg_H1[16]\ : SLE
      port map(D => \N1_data[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[16]\);
    
    next_reg_H3_cry_6_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[6]\, B => 
        hash_control_st_reg_i(6), C => R3_data(6), D => GND_net_1, 
        FCI => next_reg_H3_cry_5, S => \N3_data[6]\, Y => OPEN, 
        FCO => next_reg_H3_cry_6);
    
    next_reg_H1_cry_29_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[29]\, B => 
        hash_control_st_reg_i(6), C => R1_data(29), D => 
        GND_net_1, FCI => next_reg_H1_cry_28, S => \N1_data[29]\, 
        Y => OPEN, FCO => next_reg_H1_cry_29);
    
    next_reg_H0_cry_22_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[22]\, B => 
        hash_control_st_reg_i(6), C => R0_data(22), D => 
        GND_net_1, FCI => next_reg_H0_cry_21, S => \N0_data[22]\, 
        Y => OPEN, FCO => next_reg_H0_cry_22);
    
    next_reg_H3_cry_16_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[16]\, B => 
        hash_control_st_reg_i(6), C => R3_data(16), D => 
        GND_net_1, FCI => next_reg_H3_cry_15, S => \N3_data[16]\, 
        Y => OPEN, FCO => next_reg_H3_cry_16);
    
    \reg_H2[11]\ : SLE
      port map(D => \N2_data[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[11]\);
    
    \reg_H6[3]\ : SLE
      port map(D => \N6_data[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[3]\);
    
    \reg_H6[11]\ : SLE
      port map(D => \N6_data[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[11]\);
    
    next_reg_H1_cry_18_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[18]\, B => 
        hash_control_st_reg_i(6), C => R1_data(18), D => 
        GND_net_1, FCI => next_reg_H1_cry_17, S => \N1_data[18]\, 
        Y => OPEN, FCO => next_reg_H1_cry_18);
    
    next_reg_H0_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[20]\, B => 
        hash_control_st_reg_i(6), C => R0_data(20), D => 
        GND_net_1, FCI => next_reg_H0_cry_19, S => \N0_data[20]\, 
        Y => OPEN, FCO => next_reg_H0_cry_20);
    
    \reg_H7[22]\ : SLE
      port map(D => \N7_data[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[22]\);
    
    \reg_H3[7]\ : SLE
      port map(D => \N3_data[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[7]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \reg_H2[20]\ : SLE
      port map(D => \N2_data[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[20]\);
    
    next_reg_H5_cry_15_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[15]\, B => 
        hash_control_st_reg_i(6), C => R5_data(15), D => 
        GND_net_1, FCI => next_reg_H5_cry_14, S => \N5_data[15]\, 
        Y => OPEN, FCO => next_reg_H5_cry_15);
    
    \reg_H4[21]\ : SLE
      port map(D => \N4_data[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[21]\);
    
    next_reg_H4_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[24]\, B => 
        hash_control_st_reg_i(6), C => R4_data(24), D => 
        GND_net_1, FCI => next_reg_H4_cry_23, S => \N4_data[24]\, 
        Y => OPEN, FCO => next_reg_H4_cry_24);
    
    \reg_H7[27]\ : SLE
      port map(D => \N7_data[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[27]\);
    
    \reg_H5[19]\ : SLE
      port map(D => \N5_data[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[19]\);
    
    next_reg_H1_cry_2_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[2]\, B => 
        hash_control_st_reg_i(6), C => R1_data(2), D => GND_net_1, 
        FCI => next_reg_H1_cry_1, S => \N1_data[2]\, Y => OPEN, 
        FCO => next_reg_H1_cry_2);
    
    \reg_H1[31]\ : SLE
      port map(D => \N1_data[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[31]\);
    
    next_reg_H2_cry_29_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[29]\, B => 
        hash_control_st_reg_i(6), C => R2_data(29), D => 
        GND_net_1, FCI => next_reg_H2_cry_28, S => \N2_data[29]\, 
        Y => OPEN, FCO => next_reg_H2_cry_29);
    
    next_reg_H6_cry_25_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[25]\, B => 
        hash_control_st_reg_i(6), C => R6_data(25), D => 
        GND_net_1, FCI => next_reg_H6_cry_24, S => \N6_data[25]\, 
        Y => OPEN, FCO => next_reg_H6_cry_25);
    
    \reg_H3[18]\ : SLE
      port map(D => \N3_data[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[18]\);
    
    next_reg_H7_cry_22_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[22]\, B => 
        hash_control_st_reg_i(6), C => R7_data(22), D => 
        GND_net_1, FCI => next_reg_H7_cry_21, S => \N7_data[22]\, 
        Y => OPEN, FCO => next_reg_H7_cry_22);
    
    next_reg_H2_cry_4_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[4]\, B => 
        hash_control_st_reg_i(6), C => R2_data(4), D => GND_net_1, 
        FCI => next_reg_H2_cry_3, S => \N2_data[4]\, Y => OPEN, 
        FCO => next_reg_H2_cry_4);
    
    \reg_H5[29]\ : SLE
      port map(D => \N5_data[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[29]\);
    
    next_reg_H5_cry_22_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[22]\, B => 
        hash_control_st_reg_i(6), C => R5_data(22), D => 
        GND_net_1, FCI => next_reg_H5_cry_21, S => \N5_data[22]\, 
        Y => OPEN, FCO => next_reg_H5_cry_22);
    
    next_reg_H3_cry_5_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[5]\, B => 
        hash_control_st_reg_i(6), C => R3_data(5), D => GND_net_1, 
        FCI => next_reg_H3_cry_4, S => \N3_data[5]\, Y => OPEN, 
        FCO => next_reg_H3_cry_5);
    
    next_reg_H7_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[20]\, B => 
        hash_control_st_reg_i(6), C => R7_data(20), D => 
        GND_net_1, FCI => next_reg_H7_cry_19, S => \N7_data[20]\, 
        Y => OPEN, FCO => next_reg_H7_cry_20);
    
    next_reg_H4_cry_18_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[18]\, B => 
        hash_control_st_reg_i(6), C => R4_data(18), D => 
        GND_net_1, FCI => next_reg_H4_cry_17, S => \N4_data[18]\, 
        Y => OPEN, FCO => next_reg_H4_cry_18);
    
    next_reg_H0_cry_4_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[4]\, B => 
        hash_control_st_reg_i(6), C => R0_data(4), D => GND_net_1, 
        FCI => next_reg_H0_cry_3, S => \N0_data[4]\, Y => OPEN, 
        FCO => next_reg_H0_cry_4);
    
    \reg_H1[3]\ : SLE
      port map(D => \N1_data[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[3]\);
    
    next_reg_H7_cry_5_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[5]\, B => 
        hash_control_st_reg_i(6), C => R7_data(5), D => GND_net_1, 
        FCI => next_reg_H7_cry_4, S => \N7_data[5]\, Y => OPEN, 
        FCO => next_reg_H7_cry_5);
    
    \reg_H5[6]\ : SLE
      port map(D => \N5_data[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[6]\);
    
    next_reg_H5_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[20]\, B => 
        hash_control_st_reg_i(6), C => R5_data(20), D => 
        GND_net_1, FCI => next_reg_H5_cry_19, S => \N5_data[20]\, 
        Y => OPEN, FCO => next_reg_H5_cry_20);
    
    \reg_H2[16]\ : SLE
      port map(D => \N2_data[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[16]\);
    
    next_reg_H4_cry_9_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[9]\, B => 
        hash_control_st_reg_i(6), C => R4_data(9), D => GND_net_1, 
        FCI => next_reg_H4_cry_8, S => \N4_data[9]\, Y => OPEN, 
        FCO => next_reg_H4_cry_9);
    
    next_reg_H0_cry_19_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[19]\, B => 
        hash_control_st_reg_i(6), C => R0_data(19), D => 
        GND_net_1, FCI => next_reg_H0_cry_18, S => \N0_data[19]\, 
        Y => OPEN, FCO => next_reg_H0_cry_19);
    
    \reg_H6[16]\ : SLE
      port map(D => \N6_data[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[16]\);
    
    \reg_H1[6]\ : SLE
      port map(D => \N1_data[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[6]\);
    
    \reg_H0[10]\ : SLE
      port map(D => \N0_data[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[10]\);
    
    next_reg_H2_cry_9_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[9]\, B => 
        hash_control_st_reg_i(6), C => R2_data(9), D => GND_net_1, 
        FCI => next_reg_H2_cry_8, S => \N2_data[9]\, Y => OPEN, 
        FCO => next_reg_H2_cry_9);
    
    \reg_H7[30]\ : SLE
      port map(D => \N7_data[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[30]\);
    
    \reg_H6[4]\ : SLE
      port map(D => \N6_data[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[4]\);
    
    \reg_H4[26]\ : SLE
      port map(D => \N4_data[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[26]\);
    
    next_reg_H7_s_31 : ARI1
      generic map(INIT => x"42800")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R7_data(31), D => \SHA256_BLOCK_0_H7_o[31]\, FCI => 
        next_reg_H7_cry_30, S => \N7_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_H1_cry_11_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[11]\, B => 
        hash_control_st_reg_i(6), C => R1_data(11), D => 
        GND_net_1, FCI => next_reg_H1_cry_10, S => \N1_data[11]\, 
        Y => OPEN, FCO => next_reg_H1_cry_11);
    
    \reg_H4[5]\ : SLE
      port map(D => \N4_data[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[5]\);
    
    \reg_H3[15]\ : SLE
      port map(D => \N3_data[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[15]\);
    
    next_reg_H5_cry_8_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[8]\, B => 
        hash_control_st_reg_i(6), C => R5_data(8), D => GND_net_1, 
        FCI => next_reg_H5_cry_7, S => \N5_data[8]\, Y => OPEN, 
        FCO => next_reg_H5_cry_8);
    
    next_reg_H3_cry_19_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[19]\, B => 
        hash_control_st_reg_i(6), C => R3_data(19), D => 
        GND_net_1, FCI => next_reg_H3_cry_18, S => \N3_data[19]\, 
        Y => OPEN, FCO => next_reg_H3_cry_19);
    
    next_reg_H6_cry_16_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[16]\, B => 
        hash_control_st_reg_i(6), C => R6_data(16), D => 
        GND_net_1, FCI => next_reg_H6_cry_15, S => \N6_data[16]\, 
        Y => OPEN, FCO => next_reg_H6_cry_16);
    
    \reg_H2[29]\ : SLE
      port map(D => \N2_data[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[29]\);
    
    next_reg_H4_cry_4_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[4]\, B => 
        hash_control_st_reg_i(6), C => R4_data(4), D => GND_net_1, 
        FCI => next_reg_H4_cry_3, S => \N4_data[4]\, Y => OPEN, 
        FCO => next_reg_H4_cry_4);
    
    \reg_H3[6]\ : SLE
      port map(D => \N3_data[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[6]\);
    
    next_reg_H0_cry_7_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[7]\, B => 
        hash_control_st_reg_i(6), C => R0_data(7), D => GND_net_1, 
        FCI => next_reg_H0_cry_6, S => \N0_data[7]\, Y => OPEN, 
        FCO => next_reg_H0_cry_7);
    
    next_reg_H2_cry_8_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[8]\, B => 
        hash_control_st_reg_i(6), C => R2_data(8), D => GND_net_1, 
        FCI => next_reg_H2_cry_7, S => \N2_data[8]\, Y => OPEN, 
        FCO => next_reg_H2_cry_8);
    
    next_reg_H2_cry_12_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[12]\, B => 
        hash_control_st_reg_i(6), C => R2_data(12), D => 
        GND_net_1, FCI => next_reg_H2_cry_11, S => \N2_data[12]\, 
        Y => OPEN, FCO => next_reg_H2_cry_12);
    
    \reg_H7[23]\ : SLE
      port map(D => \N7_data[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[23]\);
    
    \reg_H7[12]\ : SLE
      port map(D => \N7_data[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[12]\);
    
    \reg_H4[1]\ : SLE
      port map(D => \N4_data[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[1]\);
    
    \reg_H0[6]\ : SLE
      port map(D => \N0_data[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[6]\);
    
    \reg_H7[24]\ : SLE
      port map(D => \N7_data[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[24]\);
    
    next_reg_H3_cry_27_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[27]\, B => 
        hash_control_st_reg_i(6), C => R3_data(27), D => 
        GND_net_1, FCI => next_reg_H3_cry_26, S => \N3_data[27]\, 
        Y => OPEN, FCO => next_reg_H3_cry_27);
    
    \reg_H1[12]\ : SLE
      port map(D => \N1_data[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[12]\);
    
    next_reg_H2_cry_10_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[10]\, B => 
        hash_control_st_reg_i(6), C => R2_data(10), D => 
        GND_net_1, FCI => next_reg_H2_cry_9, S => \N2_data[10]\, 
        Y => OPEN, FCO => next_reg_H2_cry_10);
    
    \reg_H7[17]\ : SLE
      port map(D => \N7_data[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[17]\);
    
    next_reg_H4_cry_11_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[11]\, B => 
        hash_control_st_reg_i(6), C => R4_data(11), D => 
        GND_net_1, FCI => next_reg_H4_cry_10, S => \N4_data[11]\, 
        Y => OPEN, FCO => next_reg_H4_cry_11);
    
    \reg_H1[17]\ : SLE
      port map(D => \N1_data[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[17]\);
    
    next_reg_H1_cry_22_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[22]\, B => 
        hash_control_st_reg_i(6), C => R1_data(22), D => 
        GND_net_1, FCI => next_reg_H1_cry_21, S => \N1_data[22]\, 
        Y => OPEN, FCO => next_reg_H1_cry_22);
    
    next_reg_H1_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[20]\, B => 
        hash_control_st_reg_i(6), C => R1_data(20), D => 
        GND_net_1, FCI => next_reg_H1_cry_19, S => \N1_data[20]\, 
        Y => OPEN, FCO => next_reg_H1_cry_20);
    
    next_reg_H4_cry_0_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[0]\, B => 
        hash_control_st_reg_i(6), C => R4_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H4_cry_0_0_Y\, 
        FCO => next_reg_H4_cry_0);
    
    next_reg_H3_cry_1_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[1]\, B => 
        hash_control_st_reg_i(6), C => R3_data(1), D => GND_net_1, 
        FCI => next_reg_H3_cry_0, S => \N3_data[1]\, Y => OPEN, 
        FCO => next_reg_H3_cry_1);
    
    \reg_H3[2]\ : SLE
      port map(D => \N3_data[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[2]\);
    
    \reg_H0[19]\ : SLE
      port map(D => \N0_data[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[19]\);
    
    next_reg_H4_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[28]\, B => 
        hash_control_st_reg_i(6), C => R4_data(28), D => 
        GND_net_1, FCI => next_reg_H4_cry_27, S => \N4_data[28]\, 
        Y => OPEN, FCO => next_reg_H4_cry_28);
    
    \reg_H1[20]\ : SLE
      port map(D => \N1_data[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[20]\);
    
    \reg_H5[30]\ : SLE
      port map(D => \N5_data[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[30]\);
    
    next_reg_H7_cry_16_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[16]\, B => 
        hash_control_st_reg_i(6), C => R7_data(16), D => 
        GND_net_1, FCI => next_reg_H7_cry_15, S => \N7_data[16]\, 
        Y => OPEN, FCO => next_reg_H7_cry_16);
    
    next_reg_H4_cry_1_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[1]\, B => 
        hash_control_st_reg_i(6), C => R4_data(1), D => GND_net_1, 
        FCI => next_reg_H4_cry_0, S => \N4_data[1]\, Y => OPEN, 
        FCO => next_reg_H4_cry_1);
    
    next_reg_H2_cry_22_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[22]\, B => 
        hash_control_st_reg_i(6), C => R2_data(22), D => 
        GND_net_1, FCI => next_reg_H2_cry_21, S => \N2_data[22]\, 
        Y => OPEN, FCO => next_reg_H2_cry_22);
    
    next_reg_H6_cry_19_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[19]\, B => 
        hash_control_st_reg_i(6), C => R6_data(19), D => 
        GND_net_1, FCI => next_reg_H6_cry_18, S => \N6_data[19]\, 
        Y => OPEN, FCO => next_reg_H6_cry_19);
    
    next_reg_H2_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[20]\, B => 
        hash_control_st_reg_i(6), C => R2_data(20), D => 
        GND_net_1, FCI => next_reg_H2_cry_19, S => \N2_data[20]\, 
        Y => OPEN, FCO => next_reg_H2_cry_20);
    
    \reg_H3[11]\ : SLE
      port map(D => \N3_data[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[11]\);
    
    \reg_H2[12]\ : SLE
      port map(D => \N2_data[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[12]\);
    
    \reg_H6[12]\ : SLE
      port map(D => \N6_data[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[12]\);
    
    next_reg_H0_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[23]\, B => 
        hash_control_st_reg_i(6), C => R0_data(23), D => 
        GND_net_1, FCI => next_reg_H0_cry_22, S => \N0_data[23]\, 
        Y => OPEN, FCO => next_reg_H0_cry_23);
    
    \reg_H2[17]\ : SLE
      port map(D => \N2_data[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[17]\);
    
    next_reg_H0_cry_12_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[12]\, B => 
        hash_control_st_reg_i(6), C => R0_data(12), D => 
        GND_net_1, FCI => next_reg_H0_cry_11, S => \N0_data[12]\, 
        Y => OPEN, FCO => next_reg_H0_cry_12);
    
    \reg_H6[17]\ : SLE
      port map(D => \N6_data[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[17]\);
    
    \reg_H4[22]\ : SLE
      port map(D => \N4_data[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[22]\);
    
    \reg_H3[28]\ : SLE
      port map(D => \N3_data[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[28]\);
    
    next_reg_H3_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[24]\, B => 
        hash_control_st_reg_i(6), C => R3_data(24), D => 
        GND_net_1, FCI => next_reg_H3_cry_23, S => \N3_data[24]\, 
        Y => OPEN, FCO => next_reg_H3_cry_24);
    
    next_reg_H0_cry_10_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[10]\, B => 
        hash_control_st_reg_i(6), C => R0_data(10), D => 
        GND_net_1, FCI => next_reg_H0_cry_9, S => \N0_data[10]\, 
        Y => OPEN, FCO => next_reg_H0_cry_10);
    
    next_reg_H5_cry_1_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[1]\, B => 
        hash_control_st_reg_i(6), C => R5_data(1), D => GND_net_1, 
        FCI => next_reg_H5_cry_0, S => \N5_data[1]\, Y => OPEN, 
        FCO => next_reg_H5_cry_1);
    
    \reg_H4[27]\ : SLE
      port map(D => \N4_data[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[27]\);
    
    next_reg_H5_cry_16_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[16]\, B => 
        hash_control_st_reg_i(6), C => R5_data(16), D => 
        GND_net_1, FCI => next_reg_H5_cry_15, S => \N5_data[16]\, 
        Y => OPEN, FCO => next_reg_H5_cry_16);
    
    \reg_H7[13]\ : SLE
      port map(D => \N7_data[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[13]\);
    
    \reg_H7[14]\ : SLE
      port map(D => \N7_data[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[14]\);
    
    \reg_H1[13]\ : SLE
      port map(D => \N1_data[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[13]\);
    
    next_reg_H3_cry_12_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[12]\, B => 
        hash_control_st_reg_i(6), C => R3_data(12), D => 
        GND_net_1, FCI => next_reg_H3_cry_11, S => \N3_data[12]\, 
        Y => OPEN, FCO => next_reg_H3_cry_12);
    
    \reg_H1[14]\ : SLE
      port map(D => \N1_data[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[14]\);
    
    next_reg_H7_cry_8_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[8]\, B => 
        hash_control_st_reg_i(6), C => R7_data(8), D => GND_net_1, 
        FCI => next_reg_H7_cry_7, S => \N7_data[8]\, Y => OPEN, 
        FCO => next_reg_H7_cry_8);
    
    next_reg_H5_cry_4_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[4]\, B => 
        hash_control_st_reg_i(6), C => R5_data(4), D => GND_net_1, 
        FCI => next_reg_H5_cry_3, S => \N5_data[4]\, Y => OPEN, 
        FCO => next_reg_H5_cry_4);
    
    next_reg_H4_cry_21_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[21]\, B => 
        hash_control_st_reg_i(6), C => R4_data(21), D => 
        GND_net_1, FCI => next_reg_H4_cry_20, S => \N4_data[21]\, 
        Y => OPEN, FCO => next_reg_H4_cry_21);
    
    \reg_H1[0]\ : SLE
      port map(D => \next_reg_H1_cry_0_0_Y\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[0]\);
    
    next_reg_H3_cry_10_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[10]\, B => 
        hash_control_st_reg_i(6), C => R3_data(10), D => 
        GND_net_1, FCI => next_reg_H3_cry_9, S => \N3_data[10]\, 
        Y => OPEN, FCO => next_reg_H3_cry_10);
    
    next_reg_H1_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[15]\, B => 
        hash_control_st_reg_i(6), C => R1_data(15), D => 
        GND_net_1, FCI => next_reg_H1_cry_14, S => \N1_data[15]\, 
        Y => OPEN, FCO => next_reg_H1_cry_15);
    
    \reg_H1[29]\ : SLE
      port map(D => \N1_data[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[29]\);
    
    next_reg_H7_cry_23_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[23]\, B => 
        hash_control_st_reg_i(6), C => R7_data(23), D => 
        GND_net_1, FCI => next_reg_H7_cry_22, S => \N7_data[23]\, 
        Y => OPEN, FCO => next_reg_H7_cry_23);
    
    next_reg_H6_cry_26_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[26]\, B => 
        hash_control_st_reg_i(6), C => R6_data(26), D => 
        GND_net_1, FCI => next_reg_H6_cry_25, S => \N6_data[26]\, 
        Y => OPEN, FCO => next_reg_H6_cry_26);
    
    \reg_H2[7]\ : SLE
      port map(D => \N2_data[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[7]\);
    
    next_reg_H5_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[23]\, B => 
        hash_control_st_reg_i(6), C => R5_data(23), D => 
        GND_net_1, FCI => next_reg_H5_cry_22, S => \N5_data[23]\, 
        Y => OPEN, FCO => next_reg_H5_cry_23);
    
    \reg_H3[16]\ : SLE
      port map(D => \N3_data[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[16]\);
    
    next_reg_H0_cry_3_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[3]\, B => 
        hash_control_st_reg_i(6), C => R0_data(3), D => GND_net_1, 
        FCI => next_reg_H0_cry_2, S => \N0_data[3]\, Y => OPEN, 
        FCO => next_reg_H0_cry_3);
    
    \reg_H6[28]\ : SLE
      port map(D => \N6_data[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[28]\);
    
    \reg_H3[25]\ : SLE
      port map(D => \N3_data[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[25]\);
    
    next_reg_H7_cry_19_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[19]\, B => 
        hash_control_st_reg_i(6), C => R7_data(19), D => 
        GND_net_1, FCI => next_reg_H7_cry_18, S => \N7_data[19]\, 
        Y => OPEN, FCO => next_reg_H7_cry_19);
    
    \reg_H7[2]\ : SLE
      port map(D => \N7_data[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[2]\);
    
    \reg_H2[1]\ : SLE
      port map(D => \N2_data[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[1]\);
    
    next_reg_H7_cry_9_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[9]\, B => 
        hash_control_st_reg_i(6), C => R7_data(9), D => GND_net_1, 
        FCI => next_reg_H7_cry_8, S => \N7_data[9]\, Y => OPEN, 
        FCO => next_reg_H7_cry_9);
    
    next_reg_H0_cry_0_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[0]\, B => 
        hash_control_st_reg_i(6), C => R0_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H0_cry_0_0_Y\, 
        FCO => next_reg_H0_cry_0);
    
    \reg_H2[8]\ : SLE
      port map(D => \N2_data[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[8]\);
    
    next_reg_H7_cry_0_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[0]\, B => 
        hash_control_st_reg_i(6), C => R7_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H7_cry_0_0_Y\, 
        FCO => next_reg_H7_cry_0);
    
    \reg_H5[7]\ : SLE
      port map(D => \N5_data[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[7]\);
    
    next_reg_H4_cry_15_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[15]\, B => 
        hash_control_st_reg_i(6), C => R4_data(15), D => 
        GND_net_1, FCI => next_reg_H4_cry_14, S => \N4_data[15]\, 
        Y => OPEN, FCO => next_reg_H4_cry_15);
    
    \reg_H3[1]\ : SLE
      port map(D => \N3_data[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[1]\);
    
    \reg_H0[28]\ : SLE
      port map(D => \N0_data[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[28]\);
    
    \reg_H2[13]\ : SLE
      port map(D => \N2_data[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[13]\);
    
    next_reg_H6_cry_9_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[9]\, B => 
        hash_control_st_reg_i(6), C => R6_data(9), D => GND_net_1, 
        FCI => next_reg_H6_cry_8, S => \N6_data[9]\, Y => OPEN, 
        FCO => next_reg_H6_cry_9);
    
    \reg_H6[25]\ : SLE
      port map(D => \N6_data[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[25]\);
    
    \reg_H6[13]\ : SLE
      port map(D => \N6_data[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[13]\);
    
    \reg_H2[14]\ : SLE
      port map(D => \N2_data[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[14]\);
    
    \reg_H6[14]\ : SLE
      port map(D => \N6_data[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[14]\);
    
    next_reg_H4_cry_8_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[8]\, B => 
        hash_control_st_reg_i(6), C => R4_data(8), D => GND_net_1, 
        FCI => next_reg_H4_cry_7, S => \N4_data[8]\, Y => OPEN, 
        FCO => next_reg_H4_cry_8);
    
    next_reg_H5_cry_19_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[19]\, B => 
        hash_control_st_reg_i(6), C => R5_data(19), D => 
        GND_net_1, FCI => next_reg_H5_cry_18, S => \N5_data[19]\, 
        Y => OPEN, FCO => next_reg_H5_cry_19);
    
    \reg_H7[3]\ : SLE
      port map(D => \N7_data[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[3]\);
    
    next_reg_H2_cry_13_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[13]\, B => 
        hash_control_st_reg_i(6), C => R2_data(13), D => 
        GND_net_1, FCI => next_reg_H2_cry_12, S => \N2_data[13]\, 
        Y => OPEN, FCO => next_reg_H2_cry_13);
    
    \reg_H4[23]\ : SLE
      port map(D => \N4_data[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[23]\);
    
    \reg_H7[20]\ : SLE
      port map(D => \N7_data[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[20]\);
    
    \reg_H4[24]\ : SLE
      port map(D => \N4_data[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[24]\);
    
    next_reg_H6_cry_12_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[12]\, B => 
        hash_control_st_reg_i(6), C => R6_data(12), D => 
        GND_net_1, FCI => next_reg_H6_cry_11, S => \N6_data[12]\, 
        Y => OPEN, FCO => next_reg_H6_cry_12);
    
    next_reg_H0_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[27]\, B => 
        hash_control_st_reg_i(6), C => R0_data(27), D => 
        GND_net_1, FCI => next_reg_H0_cry_26, S => \N0_data[27]\, 
        Y => OPEN, FCO => next_reg_H0_cry_27);
    
    next_reg_H6_cry_29_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[29]\, B => 
        hash_control_st_reg_i(6), C => R6_data(29), D => 
        GND_net_1, FCI => next_reg_H6_cry_28, S => \N6_data[29]\, 
        Y => OPEN, FCO => next_reg_H6_cry_29);
    
    next_reg_H6_cry_10_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[10]\, B => 
        hash_control_st_reg_i(6), C => R6_data(10), D => 
        GND_net_1, FCI => next_reg_H6_cry_9, S => \N6_data[10]\, 
        Y => OPEN, FCO => next_reg_H6_cry_10);
    
    next_reg_H1_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[23]\, B => 
        hash_control_st_reg_i(6), C => R1_data(23), D => 
        GND_net_1, FCI => next_reg_H1_cry_22, S => \N1_data[23]\, 
        Y => OPEN, FCO => next_reg_H1_cry_23);
    
    \reg_H5[8]\ : SLE
      port map(D => \N5_data[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[8]\);
    
    \reg_H0[3]\ : SLE
      port map(D => \N0_data[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[3]\);
    
    \reg_H0[25]\ : SLE
      port map(D => \N0_data[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[25]\);
    
    next_reg_H3_cry_28_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[28]\, B => 
        hash_control_st_reg_i(6), C => R3_data(28), D => 
        GND_net_1, FCI => next_reg_H3_cry_27, S => \N3_data[28]\, 
        Y => OPEN, FCO => next_reg_H3_cry_28);
    
    next_reg_H1_cry_9_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[9]\, B => 
        hash_control_st_reg_i(6), C => R1_data(9), D => GND_net_1, 
        FCI => next_reg_H1_cry_8, S => \N1_data[9]\, Y => OPEN, 
        FCO => next_reg_H1_cry_9);
    
    \reg_H3[21]\ : SLE
      port map(D => \N3_data[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[21]\);
    
    next_reg_H1_cry_7_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[7]\, B => 
        hash_control_st_reg_i(6), C => R1_data(7), D => GND_net_1, 
        FCI => next_reg_H1_cry_6, S => \N1_data[7]\, Y => OPEN, 
        FCO => next_reg_H1_cry_7);
    
    \reg_H5[2]\ : SLE
      port map(D => \N5_data[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[2]\);
    
    \reg_H0[0]\ : SLE
      port map(D => \next_reg_H0_cry_0_0_Y\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[0]\);
    
    next_reg_H7_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[27]\, B => 
        hash_control_st_reg_i(6), C => R7_data(27), D => 
        GND_net_1, FCI => next_reg_H7_cry_26, S => \N7_data[27]\, 
        Y => OPEN, FCO => next_reg_H7_cry_27);
    
    next_reg_H2_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[23]\, B => 
        hash_control_st_reg_i(6), C => R2_data(23), D => 
        GND_net_1, FCI => next_reg_H2_cry_22, S => \N2_data[23]\, 
        Y => OPEN, FCO => next_reg_H2_cry_23);
    
    \reg_H3[31]\ : SLE
      port map(D => \N3_data[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[31]\);
    
    next_reg_H5_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[27]\, B => 
        hash_control_st_reg_i(6), C => R5_data(27), D => 
        GND_net_1, FCI => next_reg_H5_cry_26, S => \N5_data[27]\, 
        Y => OPEN, FCO => next_reg_H5_cry_27);
    
    \reg_H3[12]\ : SLE
      port map(D => \N3_data[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[12]\);
    
    \reg_H0[9]\ : SLE
      port map(D => \N0_data[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[9]\);
    
    \reg_H6[0]\ : SLE
      port map(D => \next_reg_H6_cry_0_0_Y\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[0]\);
    
    \reg_H0[5]\ : SLE
      port map(D => \N0_data[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[5]\);
    
    next_reg_H4_cry_25_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[25]\, B => 
        hash_control_st_reg_i(6), C => R4_data(25), D => 
        GND_net_1, FCI => next_reg_H4_cry_24, S => \N4_data[25]\, 
        Y => OPEN, FCO => next_reg_H4_cry_25);
    
    \reg_H3[17]\ : SLE
      port map(D => \N3_data[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[17]\);
    
    next_reg_H7_cry_12_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[12]\, B => 
        hash_control_st_reg_i(6), C => R7_data(12), D => 
        GND_net_1, FCI => next_reg_H7_cry_11, S => \N7_data[12]\, 
        Y => OPEN, FCO => next_reg_H7_cry_12);
    
    \reg_H7[29]\ : SLE
      port map(D => \N7_data[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[29]\);
    
    next_reg_H0_cry_13_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[13]\, B => 
        hash_control_st_reg_i(6), C => R0_data(13), D => 
        GND_net_1, FCI => next_reg_H0_cry_12, S => \N0_data[13]\, 
        Y => OPEN, FCO => next_reg_H0_cry_13);
    
    \reg_H6[21]\ : SLE
      port map(D => \N6_data[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[21]\);
    
    next_reg_H7_cry_10_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[10]\, B => 
        hash_control_st_reg_i(6), C => R7_data(10), D => 
        GND_net_1, FCI => next_reg_H7_cry_9, S => \N7_data[10]\, 
        Y => OPEN, FCO => next_reg_H7_cry_10);
    
    \reg_H5[3]\ : SLE
      port map(D => \N5_data[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[3]\);
    
    next_reg_H6_cry_6_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[6]\, B => 
        hash_control_st_reg_i(6), C => R6_data(6), D => GND_net_1, 
        FCI => next_reg_H6_cry_5, S => \N6_data[6]\, Y => OPEN, 
        FCO => next_reg_H6_cry_6);
    
    next_reg_H0_cry_24_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[24]\, B => 
        hash_control_st_reg_i(6), C => R0_data(24), D => 
        GND_net_1, FCI => next_reg_H0_cry_23, S => \N0_data[24]\, 
        Y => OPEN, FCO => next_reg_H0_cry_24);
    
    \reg_H3[26]\ : SLE
      port map(D => \N3_data[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[26]\);
    
    next_reg_H4_cry_3_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[3]\, B => 
        hash_control_st_reg_i(6), C => R4_data(3), D => GND_net_1, 
        FCI => next_reg_H4_cry_2, S => \N4_data[3]\, Y => OPEN, 
        FCO => next_reg_H4_cry_3);
    
    next_reg_H1_cry_0_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[0]\, B => 
        hash_control_st_reg_i(6), C => R1_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H1_cry_0_0_Y\, 
        FCO => next_reg_H1_cry_0);
    
    next_reg_H3_s_31 : ARI1
      generic map(INIT => x"47D00")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R3_data(31), D => \SHA256_BLOCK_0_H3_o[31]\, FCI => 
        next_reg_H3_cry_30, S => \N3_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    \reg_H7[10]\ : SLE
      port map(D => \N7_data[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[10]\);
    
    \reg_H1[9]\ : SLE
      port map(D => \N1_data[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[9]\);
    
    next_reg_H3_cry_21_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[21]\, B => 
        hash_control_st_reg_i(6), C => R3_data(21), D => 
        GND_net_1, FCI => next_reg_H3_cry_20, S => \N3_data[21]\, 
        Y => OPEN, FCO => next_reg_H3_cry_21);
    
    next_reg_H2_cry_7_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[7]\, B => 
        hash_control_st_reg_i(6), C => R2_data(7), D => GND_net_1, 
        FCI => next_reg_H2_cry_6, S => \N2_data[7]\, Y => OPEN, 
        FCO => next_reg_H2_cry_7);
    
    next_reg_H0_cry_8_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[8]\, B => 
        hash_control_st_reg_i(6), C => R0_data(8), D => GND_net_1, 
        FCI => next_reg_H0_cry_7, S => \N0_data[8]\, Y => OPEN, 
        FCO => next_reg_H0_cry_8);
    
    next_reg_H3_cry_13_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[13]\, B => 
        hash_control_st_reg_i(6), C => R3_data(13), D => 
        GND_net_1, FCI => next_reg_H3_cry_12, S => \N3_data[13]\, 
        Y => OPEN, FCO => next_reg_H3_cry_13);
    
    \reg_H1[10]\ : SLE
      port map(D => \N1_data[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[10]\);
    
    \reg_H6[30]\ : SLE
      port map(D => \N6_data[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[30]\);
    
    next_reg_H2_cry_17_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[17]\, B => 
        hash_control_st_reg_i(6), C => R2_data(17), D => 
        GND_net_1, FCI => next_reg_H2_cry_16, S => \N2_data[17]\, 
        Y => OPEN, FCO => next_reg_H2_cry_17);
    
    \reg_H0[21]\ : SLE
      port map(D => \N0_data[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[21]\);
    
    next_reg_H1_cry_16_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[16]\, B => 
        hash_control_st_reg_i(6), C => R1_data(16), D => 
        GND_net_1, FCI => next_reg_H1_cry_15, S => \N1_data[16]\, 
        Y => OPEN, FCO => next_reg_H1_cry_16);
    
    \reg_H0[30]\ : SLE
      port map(D => \N0_data[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[30]\);
    
    \reg_H3[9]\ : SLE
      port map(D => \N3_data[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[9]\);
    
    next_reg_H5_cry_12_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[12]\, B => 
        hash_control_st_reg_i(6), C => R5_data(12), D => 
        GND_net_1, FCI => next_reg_H5_cry_11, S => \N5_data[12]\, 
        Y => OPEN, FCO => next_reg_H5_cry_12);
    
    next_reg_H0_s_31 : ARI1
      generic map(INIT => x"42800")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R0_data(31), D => \SHA256_BLOCK_0_H0_o[31]\, FCI => 
        next_reg_H0_cry_30, S => \N0_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_H5_cry_30_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[30]\, B => 
        hash_control_st_reg_i(6), C => R5_data(30), D => 
        GND_net_1, FCI => next_reg_H5_cry_29, S => \N5_data[30]\, 
        Y => OPEN, FCO => next_reg_H5_cry_30);
    
    next_reg_H5_cry_10_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[10]\, B => 
        hash_control_st_reg_i(6), C => R5_data(10), D => 
        GND_net_1, FCI => next_reg_H5_cry_9, S => \N5_data[10]\, 
        Y => OPEN, FCO => next_reg_H5_cry_10);
    
    next_reg_H7_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[24]\, B => 
        hash_control_st_reg_i(6), C => R7_data(24), D => 
        GND_net_1, FCI => next_reg_H7_cry_23, S => \N7_data[24]\, 
        Y => OPEN, FCO => next_reg_H7_cry_24);
    
    next_reg_H2_cry_1_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[1]\, B => 
        hash_control_st_reg_i(6), C => R2_data(1), D => GND_net_1, 
        FCI => next_reg_H2_cry_0, S => \N2_data[1]\, Y => OPEN, 
        FCO => next_reg_H2_cry_1);
    
    next_reg_H1_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[27]\, B => 
        hash_control_st_reg_i(6), C => R1_data(27), D => 
        GND_net_1, FCI => next_reg_H1_cry_26, S => \N1_data[27]\, 
        Y => OPEN, FCO => next_reg_H1_cry_27);
    
    \reg_H6[26]\ : SLE
      port map(D => \N6_data[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[26]\);
    
    \reg_H2[5]\ : SLE
      port map(D => \N2_data[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[5]\);
    
    next_reg_H5_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[24]\, B => 
        hash_control_st_reg_i(6), C => R5_data(24), D => 
        GND_net_1, FCI => next_reg_H5_cry_23, S => \N5_data[24]\, 
        Y => OPEN, FCO => next_reg_H5_cry_24);
    
    \reg_H7[8]\ : SLE
      port map(D => \N7_data[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[8]\);
    
    \reg_H4[18]\ : SLE
      port map(D => \N4_data[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[18]\);
    
    next_reg_H6_cry_22_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[22]\, B => 
        hash_control_st_reg_i(6), C => R6_data(22), D => 
        GND_net_1, FCI => next_reg_H6_cry_21, S => \N6_data[22]\, 
        Y => OPEN, FCO => next_reg_H6_cry_22);
    
    next_reg_H7_cry_1_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[1]\, B => 
        hash_control_st_reg_i(6), C => R7_data(1), D => GND_net_1, 
        FCI => next_reg_H7_cry_0, S => \N7_data[1]\, Y => OPEN, 
        FCO => next_reg_H7_cry_1);
    
    next_reg_H5_cry_6_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[6]\, B => 
        hash_control_st_reg_i(6), C => R5_data(6), D => GND_net_1, 
        FCI => next_reg_H5_cry_5, S => \N5_data[6]\, Y => OPEN, 
        FCO => next_reg_H5_cry_6);
    
    \reg_H5[5]\ : SLE
      port map(D => \N5_data[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[5]\);
    
    next_reg_H6_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[20]\, B => 
        hash_control_st_reg_i(6), C => R6_data(20), D => 
        GND_net_1, FCI => next_reg_H6_cry_19, S => \N6_data[20]\, 
        Y => OPEN, FCO => next_reg_H6_cry_20);
    
    \reg_H3[13]\ : SLE
      port map(D => \N3_data[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[13]\);
    
    next_reg_H3_cry_7_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[7]\, B => 
        hash_control_st_reg_i(6), C => R3_data(7), D => GND_net_1, 
        FCI => next_reg_H3_cry_6, S => \N3_data[7]\, Y => OPEN, 
        FCO => next_reg_H3_cry_7);
    
    \reg_H3[14]\ : SLE
      port map(D => \N3_data[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[14]\);
    
    next_reg_H4_cry_16_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[16]\, B => 
        hash_control_st_reg_i(6), C => R4_data(16), D => 
        GND_net_1, FCI => next_reg_H4_cry_15, S => \N4_data[16]\, 
        Y => OPEN, FCO => next_reg_H4_cry_16);
    
    \reg_H5[4]\ : SLE
      port map(D => \N5_data[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[4]\);
    
    next_reg_H4_cry_7_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[7]\, B => 
        hash_control_st_reg_i(6), C => R4_data(7), D => GND_net_1, 
        FCI => next_reg_H4_cry_6, S => \N4_data[7]\, Y => OPEN, 
        FCO => next_reg_H4_cry_7);
    
    \reg_H2[10]\ : SLE
      port map(D => \N2_data[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[10]\);
    
    next_reg_H7_cry_7_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[7]\, B => 
        hash_control_st_reg_i(6), C => R7_data(7), D => GND_net_1, 
        FCI => next_reg_H7_cry_6, S => \N7_data[7]\, Y => OPEN, 
        FCO => next_reg_H7_cry_7);
    
    \reg_H6[10]\ : SLE
      port map(D => \N6_data[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[10]\);
    
    \reg_H0[26]\ : SLE
      port map(D => \N0_data[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[26]\);
    
    next_reg_H6_cry_0_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[0]\, B => 
        hash_control_st_reg_i(6), C => R6_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H6_cry_0_0_Y\, 
        FCO => next_reg_H6_cry_0);
    
    next_reg_H2_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[27]\, B => 
        hash_control_st_reg_i(6), C => R2_data(27), D => 
        GND_net_1, FCI => next_reg_H2_cry_26, S => \N2_data[27]\, 
        Y => OPEN, FCO => next_reg_H2_cry_27);
    
    \reg_H7[19]\ : SLE
      port map(D => \N7_data[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[19]\);
    
    \reg_H1[19]\ : SLE
      port map(D => \N1_data[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[19]\);
    
    \reg_H6[7]\ : SLE
      port map(D => \N6_data[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[7]\);
    
    \reg_H5[18]\ : SLE
      port map(D => \N5_data[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[18]\);
    
    \reg_H4[20]\ : SLE
      port map(D => \N4_data[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[20]\);
    
    \reg_H4[15]\ : SLE
      port map(D => \N4_data[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[15]\);
    
    next_reg_H6_cry_13_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[13]\, B => 
        hash_control_st_reg_i(6), C => R6_data(13), D => 
        GND_net_1, FCI => next_reg_H6_cry_12, S => \N6_data[13]\, 
        Y => OPEN, FCO => next_reg_H6_cry_13);
    
    \reg_H1[30]\ : SLE
      port map(D => \N1_data[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[30]\);
    
    next_reg_H2_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[14]\, B => 
        hash_control_st_reg_i(6), C => R2_data(14), D => 
        GND_net_1, FCI => next_reg_H2_cry_13, S => \N2_data[14]\, 
        Y => OPEN, FCO => next_reg_H2_cry_14);
    
    next_reg_H1_cry_19_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[19]\, B => 
        hash_control_st_reg_i(6), C => R1_data(19), D => 
        GND_net_1, FCI => next_reg_H1_cry_18, S => \N1_data[19]\, 
        Y => OPEN, FCO => next_reg_H1_cry_19);
    
    next_reg_H0_cry_17_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[17]\, B => 
        hash_control_st_reg_i(6), C => R0_data(17), D => 
        GND_net_1, FCI => next_reg_H0_cry_16, S => \N0_data[17]\, 
        Y => OPEN, FCO => next_reg_H0_cry_17);
    
    \reg_H4[31]\ : SLE
      port map(D => \N4_data[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[31]\);
    
    \reg_H5[28]\ : SLE
      port map(D => \N5_data[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[28]\);
    
    \reg_H3[22]\ : SLE
      port map(D => \N3_data[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[22]\);
    
    next_reg_H5_cry_5_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[5]\, B => 
        hash_control_st_reg_i(6), C => R5_data(5), D => GND_net_1, 
        FCI => next_reg_H5_cry_4, S => \N5_data[5]\, Y => OPEN, 
        FCO => next_reg_H5_cry_5);
    
    next_reg_H4_cry_2_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[2]\, B => 
        hash_control_st_reg_i(6), C => R4_data(2), D => GND_net_1, 
        FCI => next_reg_H4_cry_1, S => \N4_data[2]\, Y => OPEN, 
        FCO => next_reg_H4_cry_2);
    
    next_reg_H3_cry_0_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[0]\, B => 
        hash_control_st_reg_i(6), C => R3_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H3_cry_0_0_Y\, 
        FCO => next_reg_H3_cry_0);
    
    next_reg_H1_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[24]\, B => 
        hash_control_st_reg_i(6), C => R1_data(24), D => 
        GND_net_1, FCI => next_reg_H1_cry_23, S => \N1_data[24]\, 
        Y => OPEN, FCO => next_reg_H1_cry_24);
    
    next_reg_H0_cry_28_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[28]\, B => 
        hash_control_st_reg_i(6), C => R0_data(28), D => 
        GND_net_1, FCI => next_reg_H0_cry_27, S => \N0_data[28]\, 
        Y => OPEN, FCO => next_reg_H0_cry_28);
    
    next_reg_H3_cry_3_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[3]\, B => 
        hash_control_st_reg_i(6), C => R3_data(3), D => GND_net_1, 
        FCI => next_reg_H3_cry_2, S => \N3_data[3]\, Y => OPEN, 
        FCO => next_reg_H3_cry_3);
    
    next_reg_H3_cry_17_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[17]\, B => 
        hash_control_st_reg_i(6), C => R3_data(17), D => 
        GND_net_1, FCI => next_reg_H3_cry_16, S => \N3_data[17]\, 
        Y => OPEN, FCO => next_reg_H3_cry_17);
    
    \reg_H3[27]\ : SLE
      port map(D => \N3_data[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[27]\);
    
    \reg_H5[15]\ : SLE
      port map(D => \N5_data[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[15]\);
    
    next_reg_H2_cry_30_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[30]\, B => 
        hash_control_st_reg_i(6), C => R2_data(30), D => 
        GND_net_1, FCI => next_reg_H2_cry_29, S => \N2_data[30]\, 
        Y => OPEN, FCO => next_reg_H2_cry_30);
    
    next_reg_H4_cry_19_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[19]\, B => 
        hash_control_st_reg_i(6), C => R4_data(19), D => 
        GND_net_1, FCI => next_reg_H4_cry_18, S => \N4_data[19]\, 
        Y => OPEN, FCO => next_reg_H4_cry_19);
    
    \reg_H7[6]\ : SLE
      port map(D => \N7_data[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[6]\);
    
    \reg_H2[19]\ : SLE
      port map(D => \N2_data[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[19]\);
    
    next_reg_H3_cry_25_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[25]\, B => 
        hash_control_st_reg_i(6), C => R3_data(25), D => 
        GND_net_1, FCI => next_reg_H3_cry_24, S => \N3_data[25]\, 
        Y => OPEN, FCO => next_reg_H3_cry_25);
    
    \reg_H6[19]\ : SLE
      port map(D => \N6_data[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[19]\);
    
    next_reg_H4_cry_30_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[30]\, B => 
        hash_control_st_reg_i(6), C => R4_data(30), D => 
        GND_net_1, FCI => next_reg_H4_cry_29, S => \N4_data[30]\, 
        Y => OPEN, FCO => next_reg_H4_cry_30);
    
    \reg_H5[25]\ : SLE
      port map(D => \N5_data[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[25]\);
    
    \reg_H2[28]\ : SLE
      port map(D => \N2_data[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[28]\);
    
    \reg_H6[22]\ : SLE
      port map(D => \N6_data[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[22]\);
    
    next_reg_H7_cry_13_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[13]\, B => 
        hash_control_st_reg_i(6), C => R7_data(13), D => 
        GND_net_1, FCI => next_reg_H7_cry_12, S => \N7_data[13]\, 
        Y => OPEN, FCO => next_reg_H7_cry_13);
    
    next_reg_H4_cry_26_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[26]\, B => 
        hash_control_st_reg_i(6), C => R4_data(26), D => 
        GND_net_1, FCI => next_reg_H4_cry_25, S => \N4_data[26]\, 
        Y => OPEN, FCO => next_reg_H4_cry_26);
    
    next_reg_H2_cry_24_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[24]\, B => 
        hash_control_st_reg_i(6), C => R2_data(24), D => 
        GND_net_1, FCI => next_reg_H2_cry_23, S => \N2_data[24]\, 
        Y => OPEN, FCO => next_reg_H2_cry_24);
    
    \reg_H4[29]\ : SLE
      port map(D => \N4_data[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[29]\);
    
    \reg_H3[5]\ : SLE
      port map(D => \N3_data[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[5]\);
    
    next_reg_H7_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[28]\, B => 
        hash_control_st_reg_i(6), C => R7_data(28), D => 
        GND_net_1, FCI => next_reg_H7_cry_27, S => \N7_data[28]\, 
        Y => OPEN, FCO => next_reg_H7_cry_28);
    
    \reg_H6[27]\ : SLE
      port map(D => \N6_data[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[27]\);
    
    next_reg_H5_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[28]\, B => 
        hash_control_st_reg_i(6), C => R5_data(28), D => 
        GND_net_1, FCI => next_reg_H5_cry_27, S => \N5_data[28]\, 
        Y => OPEN, FCO => next_reg_H5_cry_28);
    
    \reg_H7[9]\ : SLE
      port map(D => \N7_data[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[9]\);
    
    \reg_H1[7]\ : SLE
      port map(D => \N1_data[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[7]\);
    
    \reg_H4[11]\ : SLE
      port map(D => \N4_data[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[11]\);
    
    next_reg_H0_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[14]\, B => 
        hash_control_st_reg_i(6), C => R0_data(14), D => 
        GND_net_1, FCI => next_reg_H0_cry_13, S => \N0_data[14]\, 
        Y => OPEN, FCO => next_reg_H0_cry_14);
    
    next_reg_H4_cry_6_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[6]\, B => 
        hash_control_st_reg_i(6), C => R4_data(6), D => GND_net_1, 
        FCI => next_reg_H4_cry_5, S => \N4_data[6]\, Y => OPEN, 
        FCO => next_reg_H4_cry_6);
    
    next_reg_H0_cry_2_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[2]\, B => 
        hash_control_st_reg_i(6), C => R0_data(2), D => GND_net_1, 
        FCI => next_reg_H0_cry_1, S => \N0_data[2]\, Y => OPEN, 
        FCO => next_reg_H0_cry_2);
    
    next_reg_H0_cry_21_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[21]\, B => 
        hash_control_st_reg_i(6), C => R0_data(21), D => 
        GND_net_1, FCI => next_reg_H0_cry_20, S => \N0_data[21]\, 
        Y => OPEN, FCO => next_reg_H0_cry_21);
    
    \reg_H0[22]\ : SLE
      port map(D => \N0_data[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[22]\);
    
    \reg_H2[25]\ : SLE
      port map(D => \N2_data[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[25]\);
    
    next_reg_H2_s_31 : ARI1
      generic map(INIT => x"42800")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R2_data(31), D => \SHA256_BLOCK_0_H2_o[31]\, FCI => 
        next_reg_H2_cry_30, S => \N2_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_H1_cry_3_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[3]\, B => 
        hash_control_st_reg_i(6), C => R1_data(3), D => GND_net_1, 
        FCI => next_reg_H1_cry_2, S => \N1_data[3]\, Y => OPEN, 
        FCO => next_reg_H1_cry_3);
    
    \reg_H0[27]\ : SLE
      port map(D => \N0_data[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[27]\);
    
    \reg_H0[18]\ : SLE
      port map(D => \N0_data[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[18]\);
    
    next_reg_H5_cry_13_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[13]\, B => 
        hash_control_st_reg_i(6), C => R5_data(13), D => 
        GND_net_1, FCI => next_reg_H5_cry_12, S => \N5_data[13]\, 
        Y => OPEN, FCO => next_reg_H5_cry_13);
    
    next_reg_H3_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[14]\, B => 
        hash_control_st_reg_i(6), C => R3_data(14), D => 
        GND_net_1, FCI => next_reg_H3_cry_13, S => \N3_data[14]\, 
        Y => OPEN, FCO => next_reg_H3_cry_14);
    
    \reg_H5[1]\ : SLE
      port map(D => \N5_data[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[1]\);
    
    next_reg_H6_cry_17_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[17]\, B => 
        hash_control_st_reg_i(6), C => R6_data(17), D => 
        GND_net_1, FCI => next_reg_H6_cry_16, S => \N6_data[17]\, 
        Y => OPEN, FCO => next_reg_H6_cry_17);
    
    \reg_H3[23]\ : SLE
      port map(D => \N3_data[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[23]\);
    
    \reg_H3[24]\ : SLE
      port map(D => \N3_data[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[24]\);
    
    \reg_H5[11]\ : SLE
      port map(D => \N5_data[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[11]\);
    
    \reg_H2[3]\ : SLE
      port map(D => \N2_data[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[3]\);
    
    \reg_H2[31]\ : SLE
      port map(D => \N2_data[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[31]\);
    
    next_reg_H6_cry_23_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[23]\, B => 
        hash_control_st_reg_i(6), C => R6_data(23), D => 
        GND_net_1, FCI => next_reg_H6_cry_22, S => \N6_data[23]\, 
        Y => OPEN, FCO => next_reg_H6_cry_23);
    
    next_reg_H2_cry_18_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[18]\, B => 
        hash_control_st_reg_i(6), C => R2_data(18), D => 
        GND_net_1, FCI => next_reg_H2_cry_17, S => \N2_data[18]\, 
        Y => OPEN, FCO => next_reg_H2_cry_18);
    
    next_reg_H1_cry_12_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[12]\, B => 
        hash_control_st_reg_i(6), C => R1_data(12), D => 
        GND_net_1, FCI => next_reg_H1_cry_11, S => \N1_data[12]\, 
        Y => OPEN, FCO => next_reg_H1_cry_12);
    
    next_reg_H7_cry_21_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[21]\, B => 
        hash_control_st_reg_i(6), C => R7_data(21), D => 
        GND_net_1, FCI => next_reg_H7_cry_20, S => \N7_data[21]\, 
        Y => OPEN, FCO => next_reg_H7_cry_21);
    
    \reg_H2[4]\ : SLE
      port map(D => \N2_data[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[4]\);
    
    \reg_H4[16]\ : SLE
      port map(D => \N4_data[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[16]\);
    
    next_reg_H5_cry_21_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[21]\, B => 
        hash_control_st_reg_i(6), C => R5_data(21), D => 
        GND_net_1, FCI => next_reg_H5_cry_20, S => \N5_data[21]\, 
        Y => OPEN, FCO => next_reg_H5_cry_21);
    
    next_reg_H4_cry_29_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[29]\, B => 
        hash_control_st_reg_i(6), C => R4_data(29), D => 
        GND_net_1, FCI => next_reg_H4_cry_28, S => \N4_data[29]\, 
        Y => OPEN, FCO => next_reg_H4_cry_29);
    
    next_reg_H1_cry_10_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[10]\, B => 
        hash_control_st_reg_i(6), C => R1_data(10), D => 
        GND_net_1, FCI => next_reg_H1_cry_9, S => \N1_data[10]\, 
        Y => OPEN, FCO => next_reg_H1_cry_10);
    
    \reg_H3[10]\ : SLE
      port map(D => \N3_data[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[10]\);
    
    \reg_H5[21]\ : SLE
      port map(D => \N5_data[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[21]\);
    
    \reg_H4[9]\ : SLE
      port map(D => \N4_data[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[9]\);
    
    next_reg_H1_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[28]\, B => 
        hash_control_st_reg_i(6), C => R1_data(28), D => 
        GND_net_1, FCI => next_reg_H1_cry_27, S => \N1_data[28]\, 
        Y => OPEN, FCO => next_reg_H1_cry_28);
    
    \reg_H0[15]\ : SLE
      port map(D => \N0_data[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[15]\);
    
    \reg_H6[23]\ : SLE
      port map(D => \N6_data[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[23]\);
    
    next_reg_H1_cry_4_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[4]\, B => 
        hash_control_st_reg_i(6), C => R1_data(4), D => GND_net_1, 
        FCI => next_reg_H1_cry_3, S => \N1_data[4]\, Y => OPEN, 
        FCO => next_reg_H1_cry_4);
    
    \reg_H7[1]\ : SLE
      port map(D => \N7_data[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[1]\);
    
    \reg_H6[24]\ : SLE
      port map(D => \N6_data[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[24]\);
    
    next_reg_H4_cry_12_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[12]\, B => 
        hash_control_st_reg_i(6), C => R4_data(12), D => 
        GND_net_1, FCI => next_reg_H4_cry_11, S => \N4_data[12]\, 
        Y => OPEN, FCO => next_reg_H4_cry_12);
    
    next_reg_H7_cry_17_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[17]\, B => 
        hash_control_st_reg_i(6), C => R7_data(17), D => 
        GND_net_1, FCI => next_reg_H7_cry_16, S => \N7_data[17]\, 
        Y => OPEN, FCO => next_reg_H7_cry_17);
    
    next_reg_H4_s_31 : ARI1
      generic map(INIT => x"42800")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R4_data(31), D => \SHA256_BLOCK_0_H4_o[31]\, FCI => 
        next_reg_H4_cry_30, S => \N4_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_H3_cry_30_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[30]\, B => 
        hash_control_st_reg_i(6), C => R3_data(30), D => 
        GND_net_1, FCI => next_reg_H3_cry_29, S => \N3_data[30]\, 
        Y => OPEN, FCO => next_reg_H3_cry_30);
    
    \reg_H5[16]\ : SLE
      port map(D => \N5_data[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[16]\);
    
    \reg_H4[6]\ : SLE
      port map(D => \N4_data[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[6]\);
    
    next_reg_H4_cry_10_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[10]\, B => 
        hash_control_st_reg_i(6), C => R4_data(10), D => 
        GND_net_1, FCI => next_reg_H4_cry_9, S => \N4_data[10]\, 
        Y => OPEN, FCO => next_reg_H4_cry_10);
    
    next_reg_H2_cry_6_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[6]\, B => 
        hash_control_st_reg_i(6), C => R2_data(6), D => GND_net_1, 
        FCI => next_reg_H2_cry_5, S => \N2_data[6]\, Y => OPEN, 
        FCO => next_reg_H2_cry_6);
    
    next_reg_H2_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[28]\, B => 
        hash_control_st_reg_i(6), C => R2_data(28), D => 
        GND_net_1, FCI => next_reg_H2_cry_27, S => \N2_data[28]\, 
        Y => OPEN, FCO => next_reg_H2_cry_28);
    
    \reg_H2[6]\ : SLE
      port map(D => \N2_data[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[6]\);
    
    \reg_H1[28]\ : SLE
      port map(D => \N1_data[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[28]\);
    
    \reg_H2[2]\ : SLE
      port map(D => \N2_data[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[2]\);
    
    \reg_H0[23]\ : SLE
      port map(D => \N0_data[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[23]\);
    
    next_reg_H6_s_31 : ARI1
      generic map(INIT => x"42800")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R6_data(31), D => \SHA256_BLOCK_0_H6_o[31]\, FCI => 
        next_reg_H6_cry_30, S => \N6_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_H1_cry_5_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[5]\, B => 
        hash_control_st_reg_i(6), C => R1_data(5), D => GND_net_1, 
        FCI => next_reg_H1_cry_4, S => \N1_data[5]\, Y => OPEN, 
        FCO => next_reg_H1_cry_5);
    
    \reg_H2[21]\ : SLE
      port map(D => \N2_data[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[21]\);
    
    \reg_H0[24]\ : SLE
      port map(D => \N0_data[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[24]\);
    
    next_reg_H6_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[14]\, B => 
        hash_control_st_reg_i(6), C => R6_data(14), D => 
        GND_net_1, FCI => next_reg_H6_cry_13, S => \N6_data[14]\, 
        Y => OPEN, FCO => next_reg_H6_cry_14);
    
    next_reg_H6_cry_3_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[3]\, B => 
        hash_control_st_reg_i(6), C => R6_data(3), D => GND_net_1, 
        FCI => next_reg_H6_cry_2, S => \N6_data[3]\, Y => OPEN, 
        FCO => next_reg_H6_cry_3);
    
    next_reg_H2_cry_11_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[11]\, B => 
        hash_control_st_reg_i(6), C => R2_data(11), D => 
        GND_net_1, FCI => next_reg_H2_cry_10, S => \N2_data[11]\, 
        Y => OPEN, FCO => next_reg_H2_cry_11);
    
    next_reg_H4_cry_5_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[5]\, B => 
        hash_control_st_reg_i(6), C => R4_data(5), D => GND_net_1, 
        FCI => next_reg_H4_cry_4, S => \N4_data[5]\, Y => OPEN, 
        FCO => next_reg_H4_cry_5);
    
    \reg_H5[26]\ : SLE
      port map(D => \N5_data[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[26]\);
    
    next_reg_H7_cry_6_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[6]\, B => 
        hash_control_st_reg_i(6), C => R7_data(6), D => GND_net_1, 
        FCI => next_reg_H7_cry_5, S => \N7_data[6]\, Y => OPEN, 
        FCO => next_reg_H7_cry_6);
    
    next_reg_H0_cry_18_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[18]\, B => 
        hash_control_st_reg_i(6), C => R0_data(18), D => 
        GND_net_1, FCI => next_reg_H0_cry_17, S => \N0_data[18]\, 
        Y => OPEN, FCO => next_reg_H0_cry_18);
    
    next_reg_H1_cry_21_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[21]\, B => 
        hash_control_st_reg_i(6), C => R1_data(21), D => 
        GND_net_1, FCI => next_reg_H1_cry_20, S => \N1_data[21]\, 
        Y => OPEN, FCO => next_reg_H1_cry_21);
    
    \reg_H4[3]\ : SLE
      port map(D => \N4_data[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[3]\);
    
    \reg_H3[19]\ : SLE
      port map(D => \N3_data[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[19]\);
    
    next_reg_H0_cry_1_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[1]\, B => 
        hash_control_st_reg_i(6), C => R0_data(1), D => GND_net_1, 
        FCI => next_reg_H0_cry_0, S => \N0_data[1]\, Y => OPEN, 
        FCO => next_reg_H0_cry_1);
    
    next_reg_H5_cry_7_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[7]\, B => 
        hash_control_st_reg_i(6), C => R5_data(7), D => GND_net_1, 
        FCI => next_reg_H5_cry_6, S => \N5_data[7]\, Y => OPEN, 
        FCO => next_reg_H5_cry_7);
    
    next_reg_H6_cry_5_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[5]\, B => 
        hash_control_st_reg_i(6), C => R6_data(5), D => GND_net_1, 
        FCI => next_reg_H6_cry_4, S => \N6_data[5]\, Y => OPEN, 
        FCO => next_reg_H6_cry_5);
    
    next_reg_H5_cry_17_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[17]\, B => 
        hash_control_st_reg_i(6), C => R5_data(17), D => 
        GND_net_1, FCI => next_reg_H5_cry_16, S => \N5_data[17]\, 
        Y => OPEN, FCO => next_reg_H5_cry_17);
    
    \reg_H1[25]\ : SLE
      port map(D => \N1_data[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[25]\);
    
    next_reg_H3_cry_26_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[26]\, B => 
        hash_control_st_reg_i(6), C => R3_data(26), D => 
        GND_net_1, FCI => next_reg_H3_cry_25, S => \N3_data[26]\, 
        Y => OPEN, FCO => next_reg_H3_cry_26);
    
    next_reg_H3_cry_18_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[18]\, B => 
        hash_control_st_reg_i(6), C => R3_data(18), D => 
        GND_net_1, FCI => next_reg_H3_cry_17, S => \N3_data[18]\, 
        Y => OPEN, FCO => next_reg_H3_cry_18);
    
    next_reg_H0_cry_25_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[25]\, B => 
        hash_control_st_reg_i(6), C => R0_data(25), D => 
        GND_net_1, FCI => next_reg_H0_cry_24, S => \N0_data[25]\, 
        Y => OPEN, FCO => next_reg_H0_cry_25);
    
    next_reg_H6_cry_1_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[1]\, B => 
        hash_control_st_reg_i(6), C => R6_data(1), D => GND_net_1, 
        FCI => next_reg_H6_cry_0, S => \N6_data[1]\, Y => OPEN, 
        FCO => next_reg_H6_cry_1);
    
    next_reg_H3_cry_4_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[4]\, B => 
        hash_control_st_reg_i(6), C => R3_data(4), D => GND_net_1, 
        FCI => next_reg_H3_cry_3, S => \N3_data[4]\, Y => OPEN, 
        FCO => next_reg_H3_cry_4);
    
    next_reg_H2_cry_3_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[3]\, B => 
        hash_control_st_reg_i(6), C => R2_data(3), D => GND_net_1, 
        FCI => next_reg_H2_cry_2, S => \N2_data[3]\, Y => OPEN, 
        FCO => next_reg_H2_cry_3);
    
    \reg_H0[7]\ : SLE
      port map(D => \N0_data[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[7]\);
    
    \reg_H0[11]\ : SLE
      port map(D => \N0_data[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[11]\);
    
    next_reg_H6_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[27]\, B => 
        hash_control_st_reg_i(6), C => R6_data(27), D => 
        GND_net_1, FCI => next_reg_H6_cry_26, S => \N6_data[27]\, 
        Y => OPEN, FCO => next_reg_H6_cry_27);
    
    \reg_H2[26]\ : SLE
      port map(D => \N2_data[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_168_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[26]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_padding is

    port( raddr_pos                   : in    std_logic_vector(3 downto 2);
          Kt_addr                     : in    std_logic_vector(0 to 0);
          st_cnt_reg                  : in    std_logic_vector(6 to 6);
          hash_control_st_reg         : in    std_logic_vector(2 to 2);
          Kt_addr_fast                : in    std_logic_vector(5 downto 2);
          sha256_controller_0_bytes_o : in    std_logic_vector(1 to 1);
          W_out_2_0                   : out   std_logic_vector(5 to 5);
          W_out_i_0                   : out   std_logic_vector(2 downto 0);
          W_out_i_i_1_1               : out   std_logic_vector(31 to 31);
          W_out_2_0_1                 : out   std_logic_vector(7 to 7);
          W_out_i_i_1                 : out   std_logic_vector(31 to 31);
          W_out_2_0_a4_1_0_RNIFI1DA   : out   std_logic_vector(23 to 23);
          W_out_2_0_a4_1_0_RNI32U7B   : out   std_logic_vector(23 to 23);
          msg_bitlen                  : in    std_logic_vector(63 downto 3);
          state_2                     : in    std_logic;
          state_0                     : in    std_logic;
          state_3                     : in    std_logic;
          W_out_2_0_0_20              : out   std_logic;
          W_out_2_0_0_12              : out   std_logic;
          W_out_2_0_0_4               : out   std_logic;
          W_out_2_0_0_1               : out   std_logic;
          W_out_2_0_0_3               : out   std_logic;
          W_out_2_0_0_0               : out   std_logic;
          W_out_2_i_0_22              : out   std_logic;
          W_out_2_i_0_17              : out   std_logic;
          W_out_2_i_0_21              : out   std_logic;
          W_out_2_i_0_20              : out   std_logic;
          W_out_2_i_0_16              : out   std_logic;
          W_out_2_i_0_18              : out   std_logic;
          W_out_2_i_0_19              : out   std_logic;
          W_out_2_i_2_0               : out   std_logic;
          W_out_2_i_2_5               : out   std_logic;
          W_out_2_i_2_6               : out   std_logic;
          W_out_2_i_1_1               : out   std_logic;
          W_out_2_i_1_0               : out   std_logic;
          W_out_2_i_1_22              : out   std_logic;
          W_out_2_i_1_17              : out   std_logic;
          W_out_2_i_1_21              : out   std_logic;
          W_out_2_i_1_20              : out   std_logic;
          W_out_2_i_1_16              : out   std_logic;
          W_out_2_i_1_18              : out   std_logic;
          W_out_2_i_1_19              : out   std_logic;
          W_out_2_i_1_13              : out   std_logic;
          W_out_2_i_1_10              : out   std_logic;
          W_out_2_i_1_12              : out   std_logic;
          W_out_2_i_1_14              : out   std_logic;
          W_out_2_i_1_9               : out   std_logic;
          W_out_2_i_1_11              : out   std_logic;
          W_out_2_i_1_8               : out   std_logic;
          W_out_2_i_1_2               : out   std_logic;
          W_out_2_i_1_4               : out   std_logic;
          W_out_2_i_1_3               : out   std_logic;
          N_1696                      : in    std_logic;
          SHA256_Module_0_di_req_o    : in    std_logic;
          N_1400                      : in    std_logic;
          N_1624                      : in    std_logic;
          N_920                       : in    std_logic;
          N_1144                      : in    std_logic;
          N_1399                      : in    std_logic;
          N_1623                      : in    std_logic;
          N_919                       : in    std_logic;
          N_1143                      : in    std_logic;
          N_1401                      : in    std_logic;
          N_1625                      : in    std_logic;
          N_921                       : in    std_logic;
          N_1145                      : in    std_logic;
          one_insert                  : in    std_logic;
          N_388                       : out   std_logic;
          W_m4_e_2                    : out   std_logic;
          Kt_addr_1_rep1              : in    std_logic;
          N_102                       : in    std_logic;
          N_105                       : out   std_logic;
          ren_pos                     : in    std_logic;
          sha256_controller_0_end_o   : in    std_logic;
          Kt_addr_0_rep2              : in    std_logic;
          sha_last_blk_reg            : in    std_logic;
          sha_last_blk_next_0_o2_0    : in    std_logic;
          N_387                       : in    std_logic;
          N_98                        : out   std_logic;
          N_111                       : in    std_logic;
          N_1694                      : in    std_logic;
          N_1692                      : in    std_logic;
          N_349                       : out   std_logic;
          N_1693                      : in    std_logic;
          N_251                       : out   std_logic;
          N_1691                      : in    std_logic;
          N_248                       : out   std_logic;
          N_1690                      : in    std_logic;
          N_245                       : out   std_logic;
          N_89                        : in    std_logic;
          N_1695                      : in    std_logic;
          N_1708                      : in    std_logic;
          N_1709                      : in    std_logic;
          N_1707                      : in    std_logic;
          N_1706                      : in    std_logic;
          N_1705                      : in    std_logic;
          N_1704                      : in    std_logic;
          N_1703                      : in    std_logic;
          N_1700                      : in    std_logic;
          N_1701                      : in    std_logic;
          N_1697                      : in    std_logic;
          N_1699                      : in    std_logic;
          N_1698                      : in    std_logic;
          N_1717                      : in    std_logic;
          N_1712                      : in    std_logic;
          N_1716                      : in    std_logic;
          N_1715                      : in    std_logic;
          N_1711                      : in    std_logic;
          N_1713                      : in    std_logic;
          N_1714                      : in    std_logic;
          N_1718                      : in    std_logic;
          N_1702                      : in    std_logic;
          N_1710                      : in    std_logic;
          N_263                       : out   std_logic;
          N_301                       : out   std_logic;
          N_304                       : out   std_logic;
          N_298                       : out   std_logic;
          N_295                       : out   std_logic;
          N_292                       : out   std_logic;
          N_289                       : out   std_logic;
          N_286                       : out   std_logic;
          N_278                       : out   std_logic;
          N_275                       : out   std_logic;
          N_272                       : out   std_logic;
          N_268                       : out   std_logic;
          N_265                       : out   std_logic
        );

end sha256_padding;

architecture DEF_ARCH of sha256_padding is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal W_N_9_mux, d_m7_0, \W_out_2_i_0[9]_net_1\, d_m6_0_1_2, 
        \W_out_i_1_RNO[1]_net_1\, d_m6_1_6, 
        \W_out_i_1_RNO[0]_net_1\, d_m6_1_1_2, 
        \W_out_i_1_RNO[2]_net_1\, N_109, 
        \W_out_2_i_o2_1_0_1[16]_net_1\, N_259, 
        \W_out_2_i_o2_1_1_1[16]_net_1\, \N_388\, W_m4_e_2_net_1, 
        \W_m4_e_4\, \N_105\, \W_out_2_0_a4_2[7]\, W_N_5_mux, 
        \W_out_2_i_o2_0_d[16]_net_1\, 
        \W_out_2_i_o2_0_c[16]_net_1\, N_311, N_306_1, N_333_1, 
        \W_out_2_i_0[13]_net_1\, \W_out_2_i_0[14]_net_1\, 
        \W_out_i_i_0[31]_net_1\, N_255, \W_out_2_i_0[8]_net_1\, 
        N_3429_tz, N_300, N_93, N_303, N_297, N_294, N_291, N_288, 
        N_285, \W_out_2_i_1[13]_net_1\, \W_out_2_i_1[14]_net_1\, 
        \W_out_2_i_0[10]_net_1\, \W_out_2_i_0[12]_net_1\, 
        \W_out_2_i_0[11]_net_1\, GND_net_1, VCC_net_1
         : std_logic;

begin 

    N_388 <= \N_388\;
    W_m4_e_2 <= W_m4_e_2_net_1;
    N_105 <= \N_105\;

    \W_out_2_i_0[25]\ : CFG4
      generic map(INIT => x"0537")

      port map(A => msg_bitlen(57), B => msg_bitlen(25), C => 
        N_111, D => N_109, Y => W_out_2_i_0_17);
    
    \W_out_2_0_a2_0[15]\ : CFG2
      generic map(INIT => x"4")

      port map(A => Kt_addr(0), B => one_insert, Y => \N_388\);
    
    \W_out_2_i_a4_0[21]\ : CFG4
      generic map(INIT => x"1303")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(21), 
        C => N_109, D => N_111, Y => N_301);
    
    \W_out_2_i_1[28]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1715, B => N_311, C => d_m7_0, D => 
        W_N_9_mux, Y => W_out_2_i_1_20);
    
    \W_out_2_i_2[14]\ : CFG4
      generic map(INIT => x"F1F0")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(14), 
        C => \W_out_2_i_1[14]_net_1\, D => N_111, Y => 
        W_out_2_i_2_6);
    
    \W_out_2_i_1[8]\ : CFG4
      generic map(INIT => x"FFF1")

      port map(A => msg_bitlen(8), B => N_109, C => N_311, D => 
        \W_out_2_i_0[8]_net_1\, Y => W_out_2_i_1_0);
    
    \W_out_2_i_0[11]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1698, B => N_311, C => d_m7_0, D => 
        W_N_9_mux, Y => \W_out_2_i_0[11]_net_1\);
    
    \W_out_i_1_RNO[2]\ : CFG4
      generic map(INIT => x"4C7C")

      port map(A => N_1401, B => d_m6_1_1_2, C => raddr_pos(3), D
         => N_1625, Y => \W_out_i_1_RNO[2]_net_1\);
    
    \W_out_2_i_1[13]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1700, B => \W_out_2_i_0[13]_net_1\, C => 
        d_m7_0, D => W_N_9_mux, Y => \W_out_2_i_1[13]_net_1\);
    
    \W_out_2_0_0[6]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(38), B => msg_bitlen(6), C => 
        N_111, D => N_109, Y => W_out_2_0_0_3);
    
    \W_out_2_i_a4[19]\ : CFG3
      generic map(INIT => x"07")

      port map(A => N_1706, B => d_m7_0, C => W_N_9_mux, Y => 
        N_294);
    
    \W_out_2_i_0[10]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1697, B => N_311, C => d_m7_0, D => 
        W_N_9_mux, Y => \W_out_2_i_0[10]_net_1\);
    
    \W_out_2_i_1[22]\ : CFG4
      generic map(INIT => x"FDFC")

      port map(A => msg_bitlen(54), B => N_311, C => N_303, D => 
        N_93, Y => W_out_2_i_1_14);
    
    \W_out_2_i_0[24]\ : CFG4
      generic map(INIT => x"0537")

      port map(A => msg_bitlen(56), B => msg_bitlen(24), C => 
        N_111, D => N_109, Y => W_out_2_i_0_16);
    
    \W_m4_e_2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => st_cnt_reg(6), B => Kt_addr_fast(5), C => 
        Kt_addr_fast(2), D => hash_control_st_reg(2), Y => 
        W_m4_e_2_net_1);
    
    \W_out_2_i_a4[22]\ : CFG3
      generic map(INIT => x"07")

      port map(A => N_1709, B => d_m7_0, C => W_N_9_mux, Y => 
        N_303);
    
    \W_out_2_i_0[28]\ : CFG4
      generic map(INIT => x"0537")

      port map(A => msg_bitlen(60), B => msg_bitlen(28), C => 
        N_111, D => N_109, Y => W_out_2_i_0_20);
    
    \W_out_2_i_a4[21]\ : CFG3
      generic map(INIT => x"07")

      port map(A => N_1708, B => d_m7_0, C => W_N_9_mux, Y => 
        N_300);
    
    \W_out_i_i_0[31]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(63), B => msg_bitlen(31), C => 
        N_111, D => N_109, Y => \W_out_i_i_0[31]_net_1\);
    
    W_m4_e_4 : CFG4
      generic map(INIT => x"4000")

      port map(A => Kt_addr_fast(4), B => Kt_addr_fast(3), C => 
        W_m4_e_2_net_1, D => Kt_addr_1_rep1, Y => \W_m4_e_4\);
    
    \W_out_2_0_o2[7]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => sha_last_blk_reg, B => Kt_addr_0_rep2, C => 
        \N_105\, Y => N_109);
    
    \W_out_2_0_a4[6]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_387, B => d_m7_0, C => W_N_9_mux, D => 
        N_1693, Y => N_251);
    
    \W_out_2_0_a4_2_0[7]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => one_insert, B => SHA256_Module_0_di_req_o, C
         => sha256_controller_0_bytes_o(1), D => 
        sha256_controller_0_end_o, Y => \W_out_2_0_a4_2[7]\);
    
    \W_out_2_0_0[15]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(47), B => msg_bitlen(15), C => 
        N_111, D => N_109, Y => W_out_2_0_0_12);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \W_out_2_i_a4_0[10]\ : CFG4
      generic map(INIT => x"1033")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(42), 
        C => N_109, D => N_111, Y => N_265);
    
    \W_out_2_i_1[14]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1701, B => \W_out_2_i_0[14]_net_1\, C => 
        d_m7_0, D => W_N_9_mux, Y => \W_out_2_i_1[14]_net_1\);
    
    \W_out_i_1[2]\ : CFG4
      generic map(INIT => x"F535")

      port map(A => msg_bitlen(34), B => d_m7_0, C => N_111, D
         => \W_out_i_1_RNO[2]_net_1\, Y => W_out_i_0(2));
    
    \W_out_2_i_1[18]\ : CFG4
      generic map(INIT => x"FDFC")

      port map(A => msg_bitlen(50), B => N_311, C => N_291, D => 
        N_93, Y => W_out_2_i_1_10);
    
    \W_out_2_i_a4[20]\ : CFG3
      generic map(INIT => x"07")

      port map(A => N_1707, B => d_m7_0, C => W_N_9_mux, Y => 
        N_297);
    
    \W_out_2_i_0[8]\ : CFG4
      generic map(INIT => x"0D0F")

      port map(A => ren_pos, B => N_89, C => W_N_9_mux, D => 
        N_1695, Y => \W_out_2_i_0[8]_net_1\);
    
    \W_out_i_1[1]\ : CFG4
      generic map(INIT => x"F535")

      port map(A => msg_bitlen(33), B => d_m7_0, C => N_111, D
         => \W_out_i_1_RNO[1]_net_1\, Y => W_out_i_0(1));
    
    \W_out_2_i_0[13]\ : CFG4
      generic map(INIT => x"0357")

      port map(A => msg_bitlen(13), B => SHA256_Module_0_di_req_o, 
        C => W_N_9_mux, D => N_109, Y => \W_out_2_i_0[13]_net_1\);
    
    \W_out_2_a4[5]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_387, B => d_m7_0, C => W_N_9_mux, D => 
        N_1692, Y => N_349);
    
    \W_out_2_i_a4_0[17]\ : CFG4
      generic map(INIT => x"1303")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(17), 
        C => N_109, D => N_111, Y => N_289);
    
    \W_out_i_1_RNO_0[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => raddr_pos(3), B => raddr_pos(2), C => N_921, 
        D => N_1145, Y => d_m6_1_1_2);
    
    \W_out_2_i_1[12]\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => msg_bitlen(12), B => 
        \W_out_2_i_o2_0_d[16]_net_1\, C => 
        \W_out_2_i_o2_0_c[16]_net_1\, D => 
        \W_out_2_i_0[12]_net_1\, Y => W_out_2_i_1_4);
    
    \W_out_2_i_o2_1_0[16]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_109, B => \W_out_2_i_o2_1_0_1[16]_net_1\, Y
         => N_259);
    
    \W_out_2_0_a4_1_0_RNIFI1DA[23]\ : CFG3
      generic map(INIT => x"80")

      port map(A => d_m7_0, B => N_1702, C => N_3429_tz, Y => 
        W_out_2_0_a4_1_0_RNIFI1DA(23));
    
    \W_out_i_i_1_1[31]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => one_insert, B => N_333_1, C => 
        \W_out_i_i_0[31]_net_1\, Y => W_out_i_i_1_1(31));
    
    \W_out_2_i_1[26]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1713, B => N_311, C => d_m7_0, D => 
        W_N_9_mux, Y => W_out_2_i_1_18);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \W_out_2_i_a4_0[20]\ : CFG4
      generic map(INIT => x"1303")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(20), 
        C => N_109, D => N_111, Y => N_298);
    
    \W_out_2_0_0[4]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(36), B => msg_bitlen(4), C => 
        N_111, D => N_109, Y => W_out_2_0_0_1);
    
    \W_out_2_0_a4[4]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_387, B => d_m7_0, C => W_N_9_mux, D => 
        N_1691, Y => N_248);
    
    \W_out_2_0_0[3]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(35), B => msg_bitlen(3), C => 
        N_111, D => N_109, Y => W_out_2_0_0_0);
    
    \W_out_2_0_a4_1_0[23]\ : CFG4
      generic map(INIT => x"F200")

      port map(A => Kt_addr(0), B => sha_last_blk_reg, C => 
        \N_105\, D => SHA256_Module_0_di_req_o, Y => N_306_1);
    
    \W_out_2_i_o2_0_0[16]\ : CFG4
      generic map(INIT => x"1303")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(9), 
        C => N_109, D => N_111, Y => N_263);
    
    \W_out_2_i_1[21]\ : CFG4
      generic map(INIT => x"FDFC")

      port map(A => msg_bitlen(53), B => N_311, C => N_300, D => 
        N_93, Y => W_out_2_i_1_13);
    
    \W_out_2_i_0[14]\ : CFG4
      generic map(INIT => x"0357")

      port map(A => msg_bitlen(14), B => SHA256_Module_0_di_req_o, 
        C => W_N_9_mux, D => N_109, Y => \W_out_2_i_0[14]_net_1\);
    
    \W_out_i_1_RNO[1]\ : CFG4
      generic map(INIT => x"4C7C")

      port map(A => N_1400, B => d_m6_0_1_2, C => raddr_pos(3), D
         => N_1624, Y => \W_out_i_1_RNO[1]_net_1\);
    
    \W_out_2_i_1[27]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1714, B => N_311, C => d_m7_0, D => 
        W_N_9_mux, Y => W_out_2_i_1_19);
    
    W_out_2_0_237_0 : CFG4
      generic map(INIT => x"AAA8")

      port map(A => ren_pos, B => state_2, C => state_0, D => 
        state_3, Y => d_m7_0);
    
    \W_out_2_i_1[20]\ : CFG4
      generic map(INIT => x"FDFC")

      port map(A => msg_bitlen(52), B => N_311, C => N_297, D => 
        N_93, Y => W_out_2_i_1_12);
    
    \W_out_i_o2_0[0]\ : CFG3
      generic map(INIT => x"72")

      port map(A => W_N_5_mux, B => sha_last_blk_next_0_o2_0, C
         => N_387, Y => N_98);
    
    \W_out_2_i_0[26]\ : CFG4
      generic map(INIT => x"0537")

      port map(A => msg_bitlen(58), B => msg_bitlen(26), C => 
        N_111, D => N_109, Y => W_out_2_i_0_18);
    
    \W_out_i_i_a4_1_0[31]\ : CFG4
      generic map(INIT => x"00F7")

      port map(A => Kt_addr(0), B => sha_last_blk_reg, C => 
        \N_105\, D => SHA256_Module_0_di_req_o, Y => N_333_1);
    
    \W_out_2_i_1[9]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_109, B => \W_out_2_i_0[9]_net_1\, C => 
        \W_out_2_i_o2_1_1_1[16]_net_1\, Y => W_out_2_i_1_1);
    
    \W_out_2_i_o2_1[16]\ : CFG4
      generic map(INIT => x"0C5D")

      port map(A => \N_105\, B => N_109, C => 
        SHA256_Module_0_di_req_o, D => sha_last_blk_next_0_o2_0, 
        Y => N_93);
    
    \W_out_2_i_1[29]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1716, B => N_311, C => d_m7_0, D => 
        W_N_9_mux, Y => W_out_2_i_1_21);
    
    \W_out_2_0_a4_1_0_RNIUJM61[23]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => SHA256_Module_0_di_req_o, B => \N_388\, C => 
        N_306_1, Y => N_3429_tz);
    
    \W_out_2_i_a4_0[13]\ : CFG4
      generic map(INIT => x"1033")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(45), 
        C => N_109, D => N_111, Y => N_275);
    
    \W_out_2_i_0[12]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1699, B => N_311, C => d_m7_0, D => 
        W_N_9_mux, Y => \W_out_2_i_0[12]_net_1\);
    
    \W_out_2_i_a4_0[12]\ : CFG4
      generic map(INIT => x"1033")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(44), 
        C => N_109, D => N_111, Y => N_272);
    
    \W_out_2_0_a4_0[7]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_387, B => d_m7_0, C => W_N_9_mux, D => 
        N_1694, Y => N_255);
    
    \W_out_2_i_a4_0[19]\ : CFG4
      generic map(INIT => x"1303")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(19), 
        C => N_109, D => N_111, Y => N_295);
    
    \W_out_2_i_a4[18]\ : CFG3
      generic map(INIT => x"07")

      port map(A => N_1705, B => d_m7_0, C => W_N_9_mux, Y => 
        N_291);
    
    \W_out_2_i_0[27]\ : CFG4
      generic map(INIT => x"0537")

      port map(A => msg_bitlen(59), B => msg_bitlen(27), C => 
        N_111, D => N_109, Y => W_out_2_i_0_19);
    
    \W_out_i_1_RNO[0]\ : CFG4
      generic map(INIT => x"4C7C")

      port map(A => N_1399, B => d_m6_1_6, C => raddr_pos(3), D
         => N_1623, Y => \W_out_i_1_RNO[0]_net_1\);
    
    \W_out_2_i_a4[17]\ : CFG3
      generic map(INIT => x"07")

      port map(A => N_1704, B => d_m7_0, C => W_N_9_mux, Y => 
        N_288);
    
    \W_out_2_i_a4[16]\ : CFG3
      generic map(INIT => x"07")

      port map(A => N_1703, B => d_m7_0, C => W_N_9_mux, Y => 
        N_285);
    
    \W_out_2_i_1[16]\ : CFG4
      generic map(INIT => x"FDFC")

      port map(A => msg_bitlen(48), B => N_311, C => N_285, D => 
        N_93, Y => W_out_2_i_1_8);
    
    \W_out_i_1[0]\ : CFG4
      generic map(INIT => x"F535")

      port map(A => msg_bitlen(32), B => d_m7_0, C => N_111, D
         => \W_out_i_1_RNO[0]_net_1\, Y => W_out_i_0(0));
    
    \W_out_2_i_a4_0[14]\ : CFG4
      generic map(INIT => x"1033")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(46), 
        C => N_109, D => N_111, Y => N_278);
    
    \W_out_2_i_0[9]\ : CFG4
      generic map(INIT => x"1555")

      port map(A => W_N_9_mux, B => N_1696, C => 
        SHA256_Module_0_di_req_o, D => d_m7_0, Y => 
        \W_out_2_i_0[9]_net_1\);
    
    \W_out_2_i_o2_0_c[16]\ : CFG4
      generic map(INIT => x"08FF")

      port map(A => Kt_addr(0), B => sha_last_blk_reg, C => 
        \N_105\, D => SHA256_Module_0_di_req_o, Y => 
        \W_out_2_i_o2_0_c[16]_net_1\);
    
    \W_out_2_0[5]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(37), B => msg_bitlen(5), C => 
        N_111, D => N_109, Y => W_out_2_0(5));
    
    \W_out_2_i_2[8]\ : CFG4
      generic map(INIT => x"FF10")

      port map(A => msg_bitlen(8), B => SHA256_Module_0_di_req_o, 
        C => N_111, D => N_259, Y => W_out_2_i_2_0);
    
    \W_out_2_i_1[11]\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => msg_bitlen(11), B => 
        \W_out_2_i_o2_0_d[16]_net_1\, C => 
        \W_out_2_i_o2_0_c[16]_net_1\, D => 
        \W_out_2_i_0[11]_net_1\, Y => W_out_2_i_1_3);
    
    \W_out_2_0_a4[3]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_387, B => d_m7_0, C => W_N_9_mux, D => 
        N_1690, Y => N_245);
    
    \W_out_2_0_0[7]\ : CFG4
      generic map(INIT => x"DC50")

      port map(A => N_111, B => N_109, C => msg_bitlen(39), D => 
        \W_out_2_0_a4_2[7]\, Y => W_out_2_0_0_4);
    
    \W_out_2_i_0[29]\ : CFG4
      generic map(INIT => x"0537")

      port map(A => msg_bitlen(61), B => msg_bitlen(29), C => 
        N_111, D => N_109, Y => W_out_2_i_0_21);
    
    \W_out_2_i_1[17]\ : CFG4
      generic map(INIT => x"FDFC")

      port map(A => msg_bitlen(49), B => N_311, C => N_288, D => 
        N_93, Y => W_out_2_i_1_9);
    
    W_m4_e : CFG4
      generic map(INIT => x"80C4")

      port map(A => Kt_addr_0_rep2, B => \W_m4_e_4\, C => 
        sha_last_blk_reg, D => one_insert, Y => W_N_9_mux);
    
    \W_out_2_i_1[10]\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => msg_bitlen(10), B => 
        \W_out_2_i_o2_0_d[16]_net_1\, C => 
        \W_out_2_i_o2_0_c[16]_net_1\, D => 
        \W_out_2_i_0[10]_net_1\, Y => W_out_2_i_1_2);
    
    \W_out_2_0_o2_0[15]\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => hash_control_st_reg(2), B => Kt_addr_fast(5), 
        C => N_102, D => Kt_addr_fast(4), Y => \N_105\);
    
    \W_out_2_i_a4_0[11]\ : CFG4
      generic map(INIT => x"1033")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(43), 
        C => N_109, D => N_111, Y => N_268);
    
    \W_out_i_1_RNO_0[1]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => raddr_pos(3), B => raddr_pos(2), C => N_920, 
        D => N_1144, Y => d_m6_0_1_2);
    
    \W_out_2_0_1[7]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => N_255, B => msg_bitlen(7), C => N_109, Y => 
        W_out_2_0_1(7));
    
    \W_out_2_i_o2_1_0_1[16]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => msg_bitlen(40), B => SHA256_Module_0_di_req_o, 
        C => sha_last_blk_next_0_o2_0, D => \N_105\, Y => 
        \W_out_2_i_o2_1_0_1[16]_net_1\);
    
    \W_out_i_1_RNO_0[0]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => raddr_pos(3), B => raddr_pos(2), C => N_919, 
        D => N_1143, Y => d_m6_1_6);
    
    \W_out_2_i_a4_0[16]\ : CFG4
      generic map(INIT => x"1303")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(16), 
        C => N_109, D => N_111, Y => N_286);
    
    \W_out_2_i_1[25]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1712, B => N_311, C => d_m7_0, D => 
        W_N_9_mux, Y => W_out_2_i_1_17);
    
    \W_out_2_i_o2_0_d[16]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \N_105\, B => one_insert, C => Kt_addr(0), Y
         => \W_out_2_i_o2_0_d[16]_net_1\);
    
    \W_out_i_o2_0_RNO[0]\ : CFG4
      generic map(INIT => x"2031")

      port map(A => Kt_addr(0), B => \N_105\, C => 
        sha_last_blk_reg, D => one_insert, Y => W_N_5_mux);
    
    \W_out_2_i_a4_0[22]\ : CFG4
      generic map(INIT => x"1303")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(22), 
        C => N_109, D => N_111, Y => N_304);
    
    \W_out_2_i_2[13]\ : CFG4
      generic map(INIT => x"F1F0")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(13), 
        C => \W_out_2_i_1[13]_net_1\, D => N_111, Y => 
        W_out_2_i_2_5);
    
    \W_out_2_i_1[19]\ : CFG4
      generic map(INIT => x"FDFC")

      port map(A => msg_bitlen(51), B => N_311, C => N_294, D => 
        N_93, Y => W_out_2_i_1_11);
    
    \W_out_2_i_a4_0[18]\ : CFG4
      generic map(INIT => x"1303")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(18), 
        C => N_109, D => N_111, Y => N_292);
    
    \W_out_2_i_0[30]\ : CFG4
      generic map(INIT => x"0537")

      port map(A => msg_bitlen(62), B => msg_bitlen(30), C => 
        N_111, D => N_109, Y => W_out_2_i_0_22);
    
    \W_out_2_i_a4[24]\ : CFG2
      generic map(INIT => x"1")

      port map(A => W_N_9_mux, B => SHA256_Module_0_di_req_o, Y
         => N_311);
    
    \W_out_2_0_a4_1_0_RNI32U7B[23]\ : CFG3
      generic map(INIT => x"80")

      port map(A => d_m7_0, B => N_1710, C => N_3429_tz, Y => 
        W_out_2_0_a4_1_0_RNI32U7B(23));
    
    \W_out_i_i_1[31]\ : CFG4
      generic map(INIT => x"C800")

      port map(A => \N_388\, B => d_m7_0, C => N_306_1, D => 
        N_1718, Y => W_out_i_i_1(31));
    
    \W_out_2_i_1[30]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1717, B => N_311, C => d_m7_0, D => 
        W_N_9_mux, Y => W_out_2_i_1_22);
    
    \W_out_2_i_o2_1_1_1[16]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => msg_bitlen(41), B => SHA256_Module_0_di_req_o, 
        C => sha_last_blk_next_0_o2_0, D => \N_105\, Y => 
        \W_out_2_i_o2_1_1_1[16]_net_1\);
    
    \W_out_2_i_1[24]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_1711, B => N_311, C => d_m7_0, D => 
        W_N_9_mux, Y => W_out_2_i_1_16);
    
    \W_out_2_0_0[23]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(55), B => msg_bitlen(23), C => 
        N_111, D => N_109, Y => W_out_2_0_0_20);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_msg_sch is

    port( Wt_data                      : out   std_logic_vector(31 downto 0);
          W_out_2_0                    : in    std_logic_vector(5 to 5);
          W_out_i_0                    : in    std_logic_vector(2 downto 0);
          W_out_i_i_1_1                : in    std_logic_vector(31 to 31);
          W_out_i_i_1                  : in    std_logic_vector(31 to 31);
          W_out_2_i_0                  : in    std_logic_vector(30 downto 24);
          W_out_2_0_a4_1_0_RNI32U7B    : in    std_logic_vector(23 to 23);
          W_out_2_0_a4_1_0_RNIFI1DA    : in    std_logic_vector(23 to 23);
          W_out_2_0_1                  : in    std_logic_vector(7 to 7);
          W_out_2_0_0_3                : in    std_logic;
          W_out_2_0_0_1                : in    std_logic;
          W_out_2_0_0_0                : in    std_logic;
          W_out_2_0_0_20               : in    std_logic;
          W_out_2_0_0_12               : in    std_logic;
          W_out_2_0_0_4                : in    std_logic;
          W_out_2_i_2_0                : in    std_logic;
          W_out_2_i_2_6                : in    std_logic;
          W_out_2_i_2_5                : in    std_logic;
          W_out_2_i_1_22               : in    std_logic;
          W_out_2_i_1_21               : in    std_logic;
          W_out_2_i_1_20               : in    std_logic;
          W_out_2_i_1_19               : in    std_logic;
          W_out_2_i_1_18               : in    std_logic;
          W_out_2_i_1_17               : in    std_logic;
          W_out_2_i_1_16               : in    std_logic;
          W_out_2_i_1_0                : in    std_logic;
          W_out_2_i_1_14               : in    std_logic;
          W_out_2_i_1_13               : in    std_logic;
          W_out_2_i_1_12               : in    std_logic;
          W_out_2_i_1_11               : in    std_logic;
          W_out_2_i_1_10               : in    std_logic;
          W_out_2_i_1_9                : in    std_logic;
          W_out_2_i_1_8                : in    std_logic;
          W_out_2_i_1_4                : in    std_logic;
          W_out_2_i_1_3                : in    std_logic;
          W_out_2_i_1_2                : in    std_logic;
          W_out_2_i_1_1                : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK : in    std_logic;
          N_244_i_0                    : in    std_logic;
          next_r0_0_cry_0_Y            : out   std_logic;
          N_251                        : in    std_logic;
          ld_i_i_3                     : in    std_logic;
          N_349                        : in    std_logic;
          N_248                        : in    std_logic;
          N_245                        : in    std_logic;
          N_98                         : in    std_logic;
          N_304                        : in    std_logic;
          N_301                        : in    std_logic;
          N_298                        : in    std_logic;
          N_295                        : in    std_logic;
          N_292                        : in    std_logic;
          N_289                        : in    std_logic;
          N_286                        : in    std_logic;
          N_278                        : in    std_logic;
          N_275                        : in    std_logic;
          N_272                        : in    std_logic;
          N_268                        : in    std_logic;
          N_265                        : in    std_logic;
          N_263                        : in    std_logic
        );

end sha256_msg_sch;

architecture DEF_ARCH of sha256_msg_sch is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \r13[18]_net_1\, VCC_net_1, \r14[18]_net_1\, 
        GND_net_1, \r13[19]_net_1\, \r14[19]_net_1\, 
        \r13[20]_net_1\, \r14[20]_net_1\, \r13[21]_net_1\, 
        \r14[21]_net_1\, \r13[22]_net_1\, \r14[22]_net_1\, 
        \r13[23]_net_1\, \r14[23]_net_1\, \r13[24]_net_1\, 
        \r14[24]_net_1\, \r13[25]_net_1\, \r14[25]_net_1\, 
        \r13[26]_net_1\, \r14[26]_net_1\, \r13[27]_net_1\, 
        \r14[27]_net_1\, \r13[28]_net_1\, \r14[28]_net_1\, 
        \r13[29]_net_1\, \r14[29]_net_1\, \r13[30]_net_1\, 
        \r14[30]_net_1\, \r13[31]_net_1\, \r14[31]_net_1\, 
        \r13[3]_net_1\, \r14[3]_net_1\, \r13[4]_net_1\, 
        \r14[4]_net_1\, \r13[5]_net_1\, \r14[5]_net_1\, 
        \r13[6]_net_1\, \r14[6]_net_1\, \r13[7]_net_1\, 
        \r14[7]_net_1\, \r13[8]_net_1\, \r14[8]_net_1\, 
        \r13[9]_net_1\, \r14[9]_net_1\, \r13[10]_net_1\, 
        \r14[10]_net_1\, \r13[11]_net_1\, \r14[11]_net_1\, 
        \r13[12]_net_1\, \r14[12]_net_1\, \r13[13]_net_1\, 
        \r14[13]_net_1\, \r13[14]_net_1\, \r14[14]_net_1\, 
        \r13[15]_net_1\, \r14[15]_net_1\, \r13[16]_net_1\, 
        \r14[16]_net_1\, \r13[17]_net_1\, \r14[17]_net_1\, 
        \r15[20]_net_1\, \r15[21]_net_1\, \r15[22]_net_1\, 
        \r15[23]_net_1\, \r15[24]_net_1\, \r15[25]_net_1\, 
        \r15[26]_net_1\, \r15[27]_net_1\, \r15[28]_net_1\, 
        \r15[29]_net_1\, \r15[30]_net_1\, \r15[31]_net_1\, 
        \r13[0]_net_1\, \r14[0]_net_1\, \r13[1]_net_1\, 
        \r14[1]_net_1\, \r13[2]_net_1\, \r14[2]_net_1\, 
        \r15[5]_net_1\, \r15[6]_net_1\, \r15[7]_net_1\, 
        \r15[8]_net_1\, \r15[9]_net_1\, \r15[10]_net_1\, 
        \r15[11]_net_1\, \r15[12]_net_1\, \r15[13]_net_1\, 
        \r15[14]_net_1\, \r15[15]_net_1\, \r15[16]_net_1\, 
        \r15[17]_net_1\, \r15[18]_net_1\, \r15[19]_net_1\, 
        \r6[22]_net_1\, \r7[22]_net_1\, \r6[23]_net_1\, 
        \r7[23]_net_1\, \r6[24]_net_1\, \r7[24]_net_1\, 
        \r6[25]_net_1\, \r7[25]_net_1\, \r6[26]_net_1\, 
        \r7[26]_net_1\, \r6[27]_net_1\, \r7[27]_net_1\, 
        \r6[28]_net_1\, \r7[28]_net_1\, \r6[29]_net_1\, 
        \r7[29]_net_1\, \r6[30]_net_1\, \r7[30]_net_1\, 
        \r6[31]_net_1\, \r7[31]_net_1\, \r15[0]_net_1\, 
        \r15[1]_net_1\, \r15[2]_net_1\, \r15[3]_net_1\, 
        \r15[4]_net_1\, \r6[7]_net_1\, \r7[7]_net_1\, 
        \r6[8]_net_1\, \r7[8]_net_1\, \r6[9]_net_1\, 
        \r7[9]_net_1\, \r6[10]_net_1\, \r7[10]_net_1\, 
        \r6[11]_net_1\, \r7[11]_net_1\, \r6[12]_net_1\, 
        \r7[12]_net_1\, \r6[13]_net_1\, \r7[13]_net_1\, 
        \r6[14]_net_1\, \r7[14]_net_1\, \r6[15]_net_1\, 
        \r7[15]_net_1\, \r6[16]_net_1\, \r7[16]_net_1\, 
        \r6[17]_net_1\, \r7[17]_net_1\, \r6[18]_net_1\, 
        \r7[18]_net_1\, \r6[19]_net_1\, \r7[19]_net_1\, 
        \r6[20]_net_1\, \r7[20]_net_1\, \r6[21]_net_1\, 
        \r7[21]_net_1\, \r5[24]_net_1\, \r5[25]_net_1\, 
        \r5[26]_net_1\, \r5[27]_net_1\, \r5[28]_net_1\, 
        \r5[29]_net_1\, \r5[30]_net_1\, \r5[31]_net_1\, 
        \r6[0]_net_1\, \r7[0]_net_1\, \r6[1]_net_1\, 
        \r7[1]_net_1\, \r6[2]_net_1\, \r7[2]_net_1\, 
        \r6[3]_net_1\, \r7[3]_net_1\, \r6[4]_net_1\, 
        \r7[4]_net_1\, \r6[5]_net_1\, \r7[5]_net_1\, 
        \r6[6]_net_1\, \r7[6]_net_1\, \r5[9]_net_1\, 
        \r5[10]_net_1\, \r5[11]_net_1\, \r5[12]_net_1\, 
        \r5[13]_net_1\, \r5[14]_net_1\, \r5[15]_net_1\, 
        \r5[16]_net_1\, \r5[17]_net_1\, \r5[18]_net_1\, 
        \r5[19]_net_1\, \r5[20]_net_1\, \r5[21]_net_1\, 
        \r5[22]_net_1\, \r5[23]_net_1\, \r4[26]_net_1\, 
        \r4[27]_net_1\, \r4[28]_net_1\, \r4[29]_net_1\, 
        \r4[30]_net_1\, \r4[31]_net_1\, \r5[0]_net_1\, 
        \r5[1]_net_1\, \r5[2]_net_1\, \r5[3]_net_1\, 
        \r5[4]_net_1\, \r5[5]_net_1\, \r5[6]_net_1\, 
        \r5[7]_net_1\, \r5[8]_net_1\, \r4[11]_net_1\, 
        \r4[12]_net_1\, \r4[13]_net_1\, \r4[14]_net_1\, 
        \r4[15]_net_1\, \r4[16]_net_1\, \r4[17]_net_1\, 
        \r4[18]_net_1\, \r4[19]_net_1\, \r4[20]_net_1\, 
        \r4[21]_net_1\, \r4[22]_net_1\, \r4[23]_net_1\, 
        \r4[24]_net_1\, \r4[25]_net_1\, \r3[28]_net_1\, 
        \r3[29]_net_1\, \r3[30]_net_1\, \r3[31]_net_1\, 
        \r4[0]_net_1\, \r4[1]_net_1\, \r4[2]_net_1\, 
        \r4[3]_net_1\, \r4[4]_net_1\, \r4[5]_net_1\, 
        \r4[6]_net_1\, \r4[7]_net_1\, \r4[8]_net_1\, 
        \r4[9]_net_1\, \r4[10]_net_1\, \r3[13]_net_1\, 
        \r3[14]_net_1\, \r3[15]_net_1\, \r3[16]_net_1\, 
        \r3[17]_net_1\, \r3[18]_net_1\, \r3[19]_net_1\, 
        \r3[20]_net_1\, \r3[21]_net_1\, \r3[22]_net_1\, 
        \r3[23]_net_1\, \r3[24]_net_1\, \r3[25]_net_1\, 
        \r3[26]_net_1\, \r3[27]_net_1\, \r2[30]_net_1\, 
        \r2[31]_net_1\, \r3[0]_net_1\, \r3[1]_net_1\, 
        \r3[2]_net_1\, \r3[3]_net_1\, \r3[4]_net_1\, 
        \r3[5]_net_1\, \r3[6]_net_1\, \r3[7]_net_1\, 
        \r3[8]_net_1\, \r3[9]_net_1\, \r3[10]_net_1\, 
        \r3[11]_net_1\, \r3[12]_net_1\, \r2[15]_net_1\, 
        \r2[16]_net_1\, \r2[17]_net_1\, \r2[18]_net_1\, 
        \r2[19]_net_1\, \r2[20]_net_1\, \r2[21]_net_1\, 
        \r2[22]_net_1\, \r2[23]_net_1\, \r2[24]_net_1\, 
        \r2[25]_net_1\, \r2[26]_net_1\, \r2[27]_net_1\, 
        \r2[28]_net_1\, \r2[29]_net_1\, \r2[0]_net_1\, 
        \r2[1]_net_1\, \r2[2]_net_1\, \r2[3]_net_1\, 
        \r2[4]_net_1\, \r2[5]_net_1\, \r2[6]_net_1\, 
        \r2[7]_net_1\, \r2[8]_net_1\, \r2[9]_net_1\, 
        \r2[10]_net_1\, \r2[11]_net_1\, \r2[12]_net_1\, 
        \r2[13]_net_1\, \r2[14]_net_1\, \r1[17]_net_1\, 
        \r1[18]_net_1\, \r1[19]_net_1\, \r1[20]_net_1\, 
        \r1[21]_net_1\, \r1[22]_net_1\, \r1[23]_net_1\, 
        \r1[24]_net_1\, \r1[25]_net_1\, \r1[26]_net_1\, 
        \r1[27]_net_1\, \r1[28]_net_1\, \r1[29]_net_1\, 
        \r1[30]_net_1\, \r1[31]_net_1\, \r1[2]_net_1\, 
        \r1[3]_net_1\, \r1[4]_net_1\, \r1[5]_net_1\, 
        \r1[6]_net_1\, \r1[7]_net_1\, \r1[8]_net_1\, 
        \r1[9]_net_1\, \r1[10]_net_1\, \r1[11]_net_1\, 
        \r1[12]_net_1\, \r1[13]_net_1\, \r1[14]_net_1\, 
        \r1[15]_net_1\, \r1[16]_net_1\, \r0[19]_net_1\, 
        \Wt_data[19]\, \r0[20]_net_1\, \Wt_data[20]\, 
        \r0[21]_net_1\, \Wt_data[21]\, \r0[22]_net_1\, 
        \Wt_data[22]\, \r0[23]_net_1\, \Wt_data[23]\, 
        \r0[24]_net_1\, \Wt_data[24]\, \r0[25]_net_1\, 
        \Wt_data[25]\, \r0[26]_net_1\, \Wt_data[26]\, 
        \r0[27]_net_1\, \Wt_data[27]\, \r0[28]_net_1\, 
        \Wt_data[28]\, \r0[29]_net_1\, \Wt_data[29]\, 
        \r0[30]_net_1\, \Wt_data[30]\, \r0[31]_net_1\, 
        \Wt_data[31]\, \r1[0]_net_1\, \r1[1]_net_1\, 
        \r0[4]_net_1\, \Wt_data[4]\, \r0[5]_net_1\, \Wt_data[5]\, 
        \r0[6]_net_1\, \Wt_data[6]\, \r0[7]_net_1\, \Wt_data[7]\, 
        \r0[8]_net_1\, \Wt_data[8]\, \r0[9]_net_1\, \Wt_data[9]\, 
        \r0[10]_net_1\, \Wt_data[10]\, \r0[11]_net_1\, 
        \Wt_data[11]\, \r0[12]_net_1\, \Wt_data[12]\, 
        \r0[13]_net_1\, \Wt_data[13]\, \r0[14]_net_1\, 
        \Wt_data[14]\, \r0[15]_net_1\, \Wt_data[15]\, 
        \r0[16]_net_1\, \Wt_data[16]\, \r0[17]_net_1\, 
        \Wt_data[17]\, \r0[18]_net_1\, \Wt_data[18]\, 
        \r0[0]_net_1\, \Wt_data[0]\, \r0[1]_net_1\, \Wt_data[1]\, 
        \r0[2]_net_1\, \Wt_data[2]\, \r0[3]_net_1\, \Wt_data[3]\, 
        \r10[23]_net_1\, \r11[23]_net_1\, \r10[24]_net_1\, 
        \r11[24]_net_1\, \r10[25]_net_1\, \r11[25]_net_1\, 
        \r10[26]_net_1\, \r11[26]_net_1\, \r10[27]_net_1\, 
        \r11[27]_net_1\, \r10[28]_net_1\, \r11[28]_net_1\, 
        \r10[29]_net_1\, \r11[29]_net_1\, \r10[30]_net_1\, 
        \r11[30]_net_1\, \r10[31]_net_1\, \r11[31]_net_1\, 
        \r10[8]_net_1\, \r11[8]_net_1\, \r10[9]_net_1\, 
        \r11[9]_net_1\, \r10[10]_net_1\, \r11[10]_net_1\, 
        \r10[11]_net_1\, \r11[11]_net_1\, \r10[12]_net_1\, 
        \r11[12]_net_1\, \r10[13]_net_1\, \r11[13]_net_1\, 
        \r10[14]_net_1\, \r11[14]_net_1\, \r10[15]_net_1\, 
        \r11[15]_net_1\, \r10[16]_net_1\, \r11[16]_net_1\, 
        \r10[17]_net_1\, \r11[17]_net_1\, \r10[18]_net_1\, 
        \r11[18]_net_1\, \r10[19]_net_1\, \r11[19]_net_1\, 
        \r10[20]_net_1\, \r11[20]_net_1\, \r10[21]_net_1\, 
        \r11[21]_net_1\, \r10[22]_net_1\, \r11[22]_net_1\, 
        \r9[25]_net_1\, \r9[26]_net_1\, \r9[27]_net_1\, 
        \r9[28]_net_1\, \r9[29]_net_1\, \r9[30]_net_1\, 
        \r9[31]_net_1\, \r10[0]_net_1\, \r11[0]_net_1\, 
        \r10[1]_net_1\, \r11[1]_net_1\, \r10[2]_net_1\, 
        \r11[2]_net_1\, \r10[3]_net_1\, \r11[3]_net_1\, 
        \r10[4]_net_1\, \r11[4]_net_1\, \r10[5]_net_1\, 
        \r11[5]_net_1\, \r10[6]_net_1\, \r11[6]_net_1\, 
        \r10[7]_net_1\, \r11[7]_net_1\, \r9[10]_net_1\, 
        \r9[11]_net_1\, \r9[12]_net_1\, \r9[13]_net_1\, 
        \r9[14]_net_1\, \r9[15]_net_1\, \r9[16]_net_1\, 
        \r9[17]_net_1\, \r9[18]_net_1\, \r9[19]_net_1\, 
        \r9[20]_net_1\, \r9[21]_net_1\, \r9[22]_net_1\, 
        \r9[23]_net_1\, \r9[24]_net_1\, \r12[27]_net_1\, 
        \r12[28]_net_1\, \r12[29]_net_1\, \r12[30]_net_1\, 
        \r12[31]_net_1\, \r9[0]_net_1\, \r9[1]_net_1\, 
        \r9[2]_net_1\, \r9[3]_net_1\, \r9[4]_net_1\, 
        \r9[5]_net_1\, \r9[6]_net_1\, \r9[7]_net_1\, 
        \r9[8]_net_1\, \r9[9]_net_1\, \r12[12]_net_1\, 
        \r12[13]_net_1\, \r12[14]_net_1\, \r12[15]_net_1\, 
        \r12[16]_net_1\, \r12[17]_net_1\, \r12[18]_net_1\, 
        \r12[19]_net_1\, \r12[20]_net_1\, \r12[21]_net_1\, 
        \r12[22]_net_1\, \r12[23]_net_1\, \r12[24]_net_1\, 
        \r12[25]_net_1\, \r12[26]_net_1\, \r12[0]_net_1\, 
        \r12[1]_net_1\, \r12[2]_net_1\, \r12[3]_net_1\, 
        \r12[4]_net_1\, \r12[5]_net_1\, \r12[6]_net_1\, 
        \r12[7]_net_1\, \r12[8]_net_1\, \r12[9]_net_1\, 
        \r12[10]_net_1\, \r12[11]_net_1\, \r8[31]_net_1\, 
        \r8[16]_net_1\, \r8[17]_net_1\, \r8[18]_net_1\, 
        \r8[19]_net_1\, \r8[20]_net_1\, \r8[21]_net_1\, 
        \r8[22]_net_1\, \r8[23]_net_1\, \r8[24]_net_1\, 
        \r8[25]_net_1\, \r8[26]_net_1\, \r8[27]_net_1\, 
        \r8[28]_net_1\, \r8[29]_net_1\, \r8[30]_net_1\, 
        \r8[1]_net_1\, \r8[2]_net_1\, \r8[3]_net_1\, 
        \r8[4]_net_1\, \r8[5]_net_1\, \r8[6]_net_1\, 
        \r8[7]_net_1\, \r8[8]_net_1\, \r8[9]_net_1\, 
        \r8[10]_net_1\, \r8[11]_net_1\, \r8[12]_net_1\, 
        \r8[13]_net_1\, \r8[14]_net_1\, \r8[15]_net_1\, 
        \r8[0]_net_1\, \next_r0_0_cry_0\, \next_r0_0_cry_0_Y\, 
        sum0_5_cry_0_Y, sum0_4_cry_0_Y, \next_r0_0_cry_1\, 
        next_r0_0_cry_1_S, \sum0_4[1]\, \sum0_5[1]\, 
        \next_r0_0_cry_2\, next_r0_0_cry_2_S, \sum0_4[2]\, 
        \sum0_5[2]\, \next_r0_0_cry_3\, next_r0_0_cry_3_S, 
        \sum0_4[3]\, \sum0_5[3]\, \next_r0_0_cry_4\, 
        next_r0_0_cry_4_S, \sum0_4[4]\, \sum0_5[4]\, 
        \next_r0_0_cry_5\, next_r0_0_cry_5_S, \sum0_4[5]\, 
        \sum0_5[5]\, \next_r0_0_cry_6\, next_r0_0_cry_6_S, 
        \sum0_4[6]\, \sum0_5[6]\, \next_r0_0_cry_7\, 
        next_r0_0_cry_7_S, \sum0_4[7]\, \sum0_5[7]\, 
        \next_r0_0_cry_8\, next_r0_0_cry_8_S, \sum0_4[8]\, 
        \sum0_5[8]\, \next_r0_0_cry_9\, next_r0_0_cry_9_S, 
        \sum0_4[9]\, \sum0_5[9]\, \next_r0_0_cry_10\, 
        next_r0_0_cry_10_S, \sum0_4[10]\, \sum0_5[10]\, 
        \next_r0_0_cry_11\, next_r0_0_cry_11_S, \sum0_4[11]\, 
        \sum0_5[11]\, \next_r0_0_cry_12\, next_r0_0_cry_12_S, 
        \sum0_4[12]\, \sum0_5[12]\, \next_r0_0_cry_13\, 
        next_r0_0_cry_13_S, \sum0_4[13]\, \sum0_5[13]\, 
        \next_r0_0_cry_14\, next_r0_0_cry_14_S, \sum0_4[14]\, 
        \sum0_5[14]\, \next_r0_0_cry_15\, next_r0_0_cry_15_S, 
        \sum0_4[15]\, \sum0_5[15]\, \next_r0_0_cry_16\, 
        next_r0_0_cry_16_S, \sum0_4[16]\, \sum0_5[16]\, 
        \next_r0_0_cry_17\, next_r0_0_cry_17_S, \sum0_4[17]\, 
        \sum0_5[17]\, \next_r0_0_cry_18\, next_r0_0_cry_18_S, 
        \sum0_4[18]\, \sum0_5[18]\, \next_r0_0_cry_19\, 
        next_r0_0_cry_19_S, \sum0_4[19]\, \sum0_5[19]\, 
        \next_r0_0_cry_20\, next_r0_0_cry_20_S, \sum0_4[20]\, 
        \sum0_5[20]\, \next_r0_0_cry_21\, next_r0_0_cry_21_S, 
        \sum0_4[21]\, \sum0_5[21]\, \next_r0_0_cry_22\, 
        next_r0_0_cry_22_S, \sum0_4[22]\, \sum0_5[22]\, 
        \next_r0_0_cry_23\, next_r0_0_cry_23_S, \sum0_4[23]\, 
        \sum0_5[23]\, \next_r0_0_cry_24\, next_r0_0_cry_24_S, 
        \sum0_4[24]\, \sum0_5[24]\, \next_r0_0_cry_25\, 
        next_r0_0_cry_25_S, \sum0_4[25]\, \sum0_5[25]\, 
        \next_r0_0_cry_26\, next_r0_0_cry_26_S, \sum0_4[26]\, 
        \sum0_5[26]\, \next_r0_0_cry_27\, next_r0_0_cry_27_S, 
        \sum0_4[27]\, \sum0_5[27]\, \next_r0_0_cry_28\, 
        next_r0_0_cry_28_S, \sum0_4[28]\, \sum0_5[28]\, 
        \next_r0_0_cry_29\, next_r0_0_cry_29_S, \sum0_4[29]\, 
        \sum0_5[29]\, next_r0_0_s_31_S, \sum0_4[31]\, 
        \sum0_5[31]\, \next_r0_0_cry_30\, next_r0_0_cry_30_S, 
        \sum0_4[30]\, \sum0_5[30]\, \sum0_4_cry_0\, \s0_0[0]\, 
        \sum0_4[0]\, \sum0_4_cry_1\, \s0_0[1]\, \sum0_4_axb_1\, 
        \sum0_4_cry_2\, \s0_0[2]\, \sum0_4_axb_2\, \sum0_4_cry_3\, 
        \s0_0[3]\, \sum0_4_axb_3\, \sum0_4_cry_4\, \s0_0[4]\, 
        \sum0_4_axb_4\, \sum0_4_cry_5\, \s0_0[5]\, \sum0_4_axb_5\, 
        \sum0_4_cry_6\, \s0_0[6]\, \sum0_4_axb_6\, \sum0_4_cry_7\, 
        \s0_0[7]\, \sum0_4_axb_7\, \sum0_4_cry_8\, \s0_0[8]\, 
        \sum0_4_axb_8\, \sum0_4_cry_9\, \s0_0[9]\, \sum0_4_axb_9\, 
        \sum0_4_cry_10\, \s0_0[10]\, \sum0_4_axb_10\, 
        \sum0_4_cry_11\, \s0_0[11]\, \sum0_4_axb_11\, 
        \sum0_4_cry_12\, \s0_0[12]\, \sum0_4_axb_12\, 
        \sum0_4_cry_13\, \s0_0[13]\, \sum0_4_axb_13\, 
        \sum0_4_cry_14\, \s0_0[14]\, \sum0_4_axb_14\, 
        \sum0_4_cry_15\, \s0_0[15]\, \sum0_4_axb_15\, 
        \sum0_4_cry_16\, \s0_0[16]\, \sum0_4_axb_16\, 
        \sum0_4_cry_17\, \s0_0[17]\, \sum0_4_axb_17\, 
        \sum0_4_cry_18\, \s0_0[18]\, \sum0_4_axb_18\, 
        \sum0_4_cry_19\, \s0_0[19]\, \sum0_4_axb_19\, 
        \sum0_4_cry_20\, \s0_0[20]\, \sum0_4_axb_20\, 
        \sum0_4_cry_21\, \s0_0[21]\, \sum0_4_axb_21\, 
        \sum0_4_cry_22\, \s0_0[22]\, \sum0_4_axb_22\, 
        \sum0_4_cry_23\, \s0_0[23]\, \sum0_4_axb_23\, 
        \sum0_4_cry_24\, \s0_0[24]\, \sum0_4_axb_24\, 
        \sum0_4_cry_25\, \s0_0[25]\, \sum0_4_axb_25\, 
        \sum0_4_cry_26\, \s0_0[26]\, \sum0_4_axb_26\, 
        \sum0_4_cry_27\, \s0_0[27]\, \sum0_4_axb_27\, 
        \sum0_4_cry_28\, \s0_0[28]\, \sum0_4_axb_28\, 
        \sum0_4_cry_29\, \s0_0[29]\, \sum0_4_axb_29\, 
        \sum0_4_cry_30\, \s0_0[30]\, \sum0_4_axb_30\, 
        \sum0_5_cry_0\, \sum0_5_cry_1\, \sum0_5_cry_2\, 
        \sum0_5_cry_3\, \sum0_5_cry_4\, \sum0_5_cry_5\, 
        \sum0_5_cry_6\, \sum0_5_cry_7\, \sum0_5_cry_8\, 
        \sum0_5_cry_9\, \sum0_5_cry_10\, \sum0_5_cry_11\, 
        \sum0_5_cry_12\, \sum0_5_cry_13\, \sum0_5_cry_14\, 
        \sum0_5_cry_15\, \sum0_5_cry_16\, \sum0_5_cry_17\, 
        \sum0_5_cry_18\, \sum0_5_cry_19\, \sum0_5_cry_20\, 
        \sum0_5_cry_21\, \sum0_5_cry_22\, \sum0_5_cry_23\, 
        \sum0_5_cry_24\, \sum0_5_cry_25\, \sum0_5_cry_26\, 
        \sum0_5_cry_27\, \sum0_5_cry_28\, \sum0_5_cry_29\, 
        \sum0_5_cry_30\, \s0[29]_net_1\, \s0[30]_net_1\, 
        \s0[21]_net_1\, \s0[22]_net_1\, \s0[23]_net_1\, 
        \s0[24]_net_1\, \s0[25]_net_1\, \s0[26]_net_1\, 
        \s0[27]_net_1\, \s0[28]_net_1\, \s0[6]_net_1\, 
        \s0[7]_net_1\, \s0[8]_net_1\, \s0[9]_net_1\, 
        \s0[10]_net_1\, \s0[11]_net_1\, \s0[12]_net_1\, 
        \s0[13]_net_1\, \s0[14]_net_1\, \s0[15]_net_1\, 
        \s0[16]_net_1\, \s0[17]_net_1\, \s0[18]_net_1\, 
        \s0[19]_net_1\, \s0[20]_net_1\, \s0[0]_net_1\, 
        \s0[1]_net_1\, \s0[2]_net_1\, \s0[3]_net_1\, 
        \s0[4]_net_1\, \s0[5]_net_1\ : std_logic;

begin 

    Wt_data(31) <= \Wt_data[31]\;
    Wt_data(30) <= \Wt_data[30]\;
    Wt_data(29) <= \Wt_data[29]\;
    Wt_data(28) <= \Wt_data[28]\;
    Wt_data(27) <= \Wt_data[27]\;
    Wt_data(26) <= \Wt_data[26]\;
    Wt_data(25) <= \Wt_data[25]\;
    Wt_data(24) <= \Wt_data[24]\;
    Wt_data(23) <= \Wt_data[23]\;
    Wt_data(22) <= \Wt_data[22]\;
    Wt_data(21) <= \Wt_data[21]\;
    Wt_data(20) <= \Wt_data[20]\;
    Wt_data(19) <= \Wt_data[19]\;
    Wt_data(18) <= \Wt_data[18]\;
    Wt_data(17) <= \Wt_data[17]\;
    Wt_data(16) <= \Wt_data[16]\;
    Wt_data(15) <= \Wt_data[15]\;
    Wt_data(14) <= \Wt_data[14]\;
    Wt_data(13) <= \Wt_data[13]\;
    Wt_data(12) <= \Wt_data[12]\;
    Wt_data(11) <= \Wt_data[11]\;
    Wt_data(10) <= \Wt_data[10]\;
    Wt_data(9) <= \Wt_data[9]\;
    Wt_data(8) <= \Wt_data[8]\;
    Wt_data(7) <= \Wt_data[7]\;
    Wt_data(6) <= \Wt_data[6]\;
    Wt_data(5) <= \Wt_data[5]\;
    Wt_data(4) <= \Wt_data[4]\;
    Wt_data(3) <= \Wt_data[3]\;
    Wt_data(2) <= \Wt_data[2]\;
    Wt_data(1) <= \Wt_data[1]\;
    Wt_data(0) <= \Wt_data[0]\;
    next_r0_0_cry_0_Y <= \next_r0_0_cry_0_Y\;

    \r4[9]\ : SLE
      port map(D => \r5[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[9]_net_1\);
    
    \r5[22]\ : SLE
      port map(D => \r6[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[22]_net_1\);
    
    \r12[21]\ : SLE
      port map(D => \r13[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[21]_net_1\);
    
    \r12[0]\ : SLE
      port map(D => \r13[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[0]_net_1\);
    
    \r10[21]\ : SLE
      port map(D => \r11[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[21]_net_1\);
    
    sum0_4_cry_0_1030 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[12]_net_1\, B => \r2[1]_net_1\, C => 
        \r2[29]_net_1\, Y => \s0_0[26]\);
    
    \r1[13]\ : SLE
      port map(D => \r2[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[13]_net_1\);
    
    sum0_4_cry_0 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[0]\, C => \sum0_4[0]\, 
        D => GND_net_1, FCI => GND_net_1, S => OPEN, Y => 
        sum0_4_cry_0_Y, FCO => \sum0_4_cry_0\);
    
    \r9[18]\ : SLE
      port map(D => \r10[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[18]_net_1\);
    
    \r6[0]\ : SLE
      port map(D => \r7[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[0]_net_1\);
    
    \r9[29]\ : SLE
      port map(D => \r10[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[29]_net_1\);
    
    \r6[9]\ : SLE
      port map(D => \r7[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[9]_net_1\);
    
    \r13[28]\ : SLE
      port map(D => \r14[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[28]_net_1\);
    
    \r3[24]\ : SLE
      port map(D => \r4[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[24]_net_1\);
    
    \r15[14]\ : SLE
      port map(D => \r0[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[14]_net_1\);
    
    \r3[18]\ : SLE
      port map(D => \r4[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[18]_net_1\);
    
    \r3[3]\ : SLE
      port map(D => \r4[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[3]_net_1\);
    
    sum0_4_cry_0_1041 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[18]_net_1\, B => \r2[1]_net_1\, C => 
        \r2[22]_net_1\, Y => \s0_0[15]\);
    
    \next_r0[14]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_278, C => next_r0_0_cry_14_S, 
        D => W_out_2_i_2_6, Y => \Wt_data[14]\);
    
    \next_r0[17]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_289, C => next_r0_0_cry_17_S, 
        D => W_out_2_i_1_9, Y => \Wt_data[17]\);
    
    \r15[12]\ : SLE
      port map(D => \r0[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[12]_net_1\);
    
    \r15[24]\ : SLE
      port map(D => \r0[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[24]_net_1\);
    
    \r5[31]\ : SLE
      port map(D => \r6[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[31]_net_1\);
    
    sum0_4_cry_20 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[20]\, C => 
        \sum0_4_axb_20\, D => GND_net_1, FCI => \sum0_4_cry_19\, 
        S => \sum0_4[20]\, Y => OPEN, FCO => \sum0_4_cry_20\);
    
    \r15[22]\ : SLE
      port map(D => \r0[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[22]_net_1\);
    
    \r15[31]\ : SLE
      port map(D => \r0[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[31]_net_1\);
    
    \r13[3]\ : SLE
      port map(D => \r14[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[3]_net_1\);
    
    \r4[17]\ : SLE
      port map(D => \r5[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[17]_net_1\);
    
    \r0[3]\ : SLE
      port map(D => \Wt_data[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[3]_net_1\);
    
    sum0_5_cry_11 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[11]_net_1\, B => \r10[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_10\, S => 
        \sum0_5[11]\, Y => OPEN, FCO => \sum0_5_cry_11\);
    
    sum0_5_cry_4 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[4]_net_1\, B => \r10[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_3\, S => 
        \sum0_5[4]\, Y => OPEN, FCO => \sum0_5_cry_4\);
    
    \r14[13]\ : SLE
      port map(D => \r15[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[13]_net_1\);
    
    \next_r0[18]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_292, C => next_r0_0_cry_18_S, 
        D => W_out_2_i_1_10, Y => \Wt_data[18]\);
    
    \r0[7]\ : SLE
      port map(D => \Wt_data[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[7]_net_1\);
    
    \r10[11]\ : SLE
      port map(D => \r11[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[11]_net_1\);
    
    \r11[0]\ : SLE
      port map(D => \r12[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[0]_net_1\);
    
    \r2[5]\ : SLE
      port map(D => \r3[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[5]_net_1\);
    
    \r5[5]\ : SLE
      port map(D => \r6[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[5]_net_1\);
    
    \r14[25]\ : SLE
      port map(D => \r15[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[25]_net_1\);
    
    next_r0_0_cry_0 : ARI1
      generic map(INIT => x"555AA")

      port map(A => sum0_5_cry_0_Y, B => sum0_4_cry_0_Y, C => 
        GND_net_1, D => GND_net_1, FCI => GND_net_1, S => OPEN, Y
         => \next_r0_0_cry_0_Y\, FCO => \next_r0_0_cry_0\);
    
    sum0_4_cry_23 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[23]\, C => 
        \sum0_4_axb_23\, D => GND_net_1, FCI => \sum0_4_cry_22\, 
        S => \sum0_4[23]\, Y => OPEN, FCO => \sum0_4_cry_23\);
    
    \r14[19]\ : SLE
      port map(D => \r15[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[19]_net_1\);
    
    \next_r0[23]\ : CFG4
      generic map(INIT => x"FE54")

      port map(A => ld_i_i_3, B => W_out_2_0_0_20, C => 
        W_out_2_0_a4_1_0_RNI32U7B(23), D => next_r0_0_cry_23_S, Y
         => \Wt_data[23]\);
    
    sum0_4_cry_0_1031 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[11]_net_1\, B => \r2[0]_net_1\, C => 
        \r2[28]_net_1\, Y => \s0_0[25]\);
    
    next_r0_0_cry_11 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[11]\, B => \sum0_5[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_10\, S
         => next_r0_0_cry_11_S, Y => OPEN, FCO => 
        \next_r0_0_cry_11\);
    
    \r12[9]\ : SLE
      port map(D => \r13[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[9]_net_1\);
    
    sum0_4_cry_17 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[17]\, C => 
        \sum0_4_axb_17\, D => GND_net_1, FCI => \sum0_4_cry_16\, 
        S => \sum0_4[17]\, Y => OPEN, FCO => \sum0_4_cry_17\);
    
    next_r0_0_cry_21 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[21]\, B => \sum0_5[21]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_20\, S
         => next_r0_0_cry_21_S, Y => OPEN, FCO => 
        \next_r0_0_cry_21\);
    
    \r7[17]\ : SLE
      port map(D => \r8[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[17]_net_1\);
    
    \r8[9]\ : SLE
      port map(D => \r9[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[9]_net_1\);
    
    \r0[29]\ : SLE
      port map(D => \Wt_data[29]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[29]_net_1\);
    
    \r13[21]\ : SLE
      port map(D => \r14[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[21]_net_1\);
    
    \r0[19]\ : SLE
      port map(D => \Wt_data[19]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[19]_net_1\);
    
    sum0_4_cry_28 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[28]\, C => 
        \sum0_4_axb_28\, D => GND_net_1, FCI => \sum0_4_cry_27\, 
        S => \sum0_4[28]\, Y => OPEN, FCO => \sum0_4_cry_28\);
    
    \s0[4]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[22]_net_1\, B => \r2[11]_net_1\, C => 
        \r2[7]_net_1\, Y => \s0[4]_net_1\);
    
    \r6[2]\ : SLE
      port map(D => \r7[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[2]_net_1\);
    
    \r4[18]\ : SLE
      port map(D => \r5[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[18]_net_1\);
    
    \r1[24]\ : SLE
      port map(D => \r2[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[24]_net_1\);
    
    \r5[14]\ : SLE
      port map(D => \r6[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[14]_net_1\);
    
    \s0[5]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[23]_net_1\, B => \r2[12]_net_1\, C => 
        \r2[8]_net_1\, Y => \s0[5]_net_1\);
    
    \r5[8]\ : SLE
      port map(D => \r6[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[8]_net_1\);
    
    \r7[26]\ : SLE
      port map(D => \r8[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[26]_net_1\);
    
    \r4[24]\ : SLE
      port map(D => \r5[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[24]_net_1\);
    
    sum0_4_cry_0_1055 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[19]_net_1\, B => \r2[8]_net_1\, C => 
        \r2[4]_net_1\, Y => \s0_0[1]\);
    
    \r15[16]\ : SLE
      port map(D => \r0[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[16]_net_1\);
    
    \r14[14]\ : SLE
      port map(D => \r15[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[14]_net_1\);
    
    \s0[6]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[24]_net_1\, B => \r2[13]_net_1\, C => 
        \r2[9]_net_1\, Y => \s0[6]_net_1\);
    
    \r15[3]\ : SLE
      port map(D => \r0[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[3]_net_1\);
    
    \r15[26]\ : SLE
      port map(D => \r0[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[26]_net_1\);
    
    \r14[12]\ : SLE
      port map(D => \r15[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[12]_net_1\);
    
    \s0[25]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[11]_net_1\, B => \r2[0]_net_1\, C => 
        \r2[28]_net_1\, Y => \s0[25]_net_1\);
    
    \r9[15]\ : SLE
      port map(D => \r10[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[15]_net_1\);
    
    \s0[15]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[18]_net_1\, B => \r2[1]_net_1\, C => 
        \r2[22]_net_1\, Y => \s0[15]_net_1\);
    
    \r8[29]\ : SLE
      port map(D => \r9[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[29]_net_1\);
    
    \r1[17]\ : SLE
      port map(D => \r2[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[17]_net_1\);
    
    \r2[14]\ : SLE
      port map(D => \r3[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[14]_net_1\);
    
    \r11[8]\ : SLE
      port map(D => \r12[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[8]_net_1\);
    
    \r11[2]\ : SLE
      port map(D => \r12[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[2]_net_1\);
    
    \r7[21]\ : SLE
      port map(D => \r8[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[21]_net_1\);
    
    \r6[26]\ : SLE
      port map(D => \r7[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[26]_net_1\);
    
    \r3[15]\ : SLE
      port map(D => \r4[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[15]_net_1\);
    
    sum0_5_cry_30 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[30]_net_1\, B => \r10[30]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_29\, S => 
        \sum0_5[30]\, Y => OPEN, FCO => \sum0_5_cry_30\);
    
    \r11[30]\ : SLE
      port map(D => \r12[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[30]_net_1\);
    
    \r7[18]\ : SLE
      port map(D => \r8[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[18]_net_1\);
    
    \r13[30]\ : SLE
      port map(D => \r14[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[30]_net_1\);
    
    \r4[5]\ : SLE
      port map(D => \r5[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[5]_net_1\);
    
    next_r0_0_cry_18 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[18]\, B => \sum0_5[18]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_17\, S
         => next_r0_0_cry_18_S, Y => OPEN, FCO => 
        \next_r0_0_cry_18\);
    
    \r7[3]\ : SLE
      port map(D => \r8[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[3]_net_1\);
    
    next_r0_0_cry_28 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[28]\, B => \sum0_5[28]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_27\, S
         => next_r0_0_cry_28_S, Y => OPEN, FCO => 
        \next_r0_0_cry_28\);
    
    \r6[21]\ : SLE
      port map(D => \r7[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[21]_net_1\);
    
    \r14[27]\ : SLE
      port map(D => \r15[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[27]_net_1\);
    
    \r8[31]\ : SLE
      port map(D => \r9[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[31]_net_1\);
    
    \r2[1]\ : SLE
      port map(D => \r3[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[1]_net_1\);
    
    sum0_4_axb_28 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[13]_net_1\, B => \s0[28]_net_1\, C => 
        \r15[15]_net_1\, Y => \sum0_4_axb_28\);
    
    \r12[6]\ : SLE
      port map(D => \r13[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[6]_net_1\);
    
    sum0_5_cry_6 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[6]_net_1\, B => \r10[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_5\, S => 
        \sum0_5[6]\, Y => OPEN, FCO => \sum0_5_cry_6\);
    
    sum0_4_cry_14 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[14]\, C => 
        \sum0_4_axb_14\, D => GND_net_1, FCI => \sum0_4_cry_13\, 
        S => \sum0_4[14]\, Y => OPEN, FCO => \sum0_4_cry_14\);
    
    \r9[24]\ : SLE
      port map(D => \r10[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[24]_net_1\);
    
    \r8[10]\ : SLE
      port map(D => \r9[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[10]_net_1\);
    
    \r6[3]\ : SLE
      port map(D => \r7[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[3]_net_1\);
    
    \r8[3]\ : SLE
      port map(D => \r9[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[3]_net_1\);
    
    \s0[8]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[26]_net_1\, B => \r2[15]_net_1\, C => 
        \r2[11]_net_1\, Y => \s0[8]_net_1\);
    
    \r7[23]\ : SLE
      port map(D => \r8[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[23]_net_1\);
    
    \r15[5]\ : SLE
      port map(D => \r0[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[5]_net_1\);
    
    \r9[12]\ : SLE
      port map(D => \r10[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[12]_net_1\);
    
    \r1[18]\ : SLE
      port map(D => \r2[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[18]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    sum0_4_cry_29 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[29]\, C => 
        \sum0_4_axb_29\, D => GND_net_1, FCI => \sum0_4_cry_28\, 
        S => \sum0_4[29]\, Y => OPEN, FCO => \sum0_4_cry_29\);
    
    sum0_5_cry_21 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[21]_net_1\, B => \r10[21]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_20\, S => 
        \sum0_5[21]\, Y => OPEN, FCO => \sum0_5_cry_21\);
    
    \next_r0[13]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_275, C => next_r0_0_cry_13_S, 
        D => W_out_2_i_2_5, Y => \Wt_data[13]\);
    
    \r3[12]\ : SLE
      port map(D => \r4[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[12]_net_1\);
    
    \r6[16]\ : SLE
      port map(D => \r7[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[16]_net_1\);
    
    \r2[2]\ : SLE
      port map(D => \r3[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[2]_net_1\);
    
    \r14[16]\ : SLE
      port map(D => \r15[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[16]_net_1\);
    
    \r2[26]\ : SLE
      port map(D => \r3[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[26]_net_1\);
    
    \r9[0]\ : SLE
      port map(D => \r10[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[0]_net_1\);
    
    \r6[23]\ : SLE
      port map(D => \r7[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[23]_net_1\);
    
    sum0_4_cry_26 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[26]\, C => 
        \sum0_4_axb_26\, D => GND_net_1, FCI => \sum0_4_cry_25\, 
        S => \sum0_4[26]\, Y => OPEN, FCO => \sum0_4_cry_26\);
    
    sum0_5_cry_10 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[10]_net_1\, B => \r10[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_9\, S => 
        \sum0_5[10]\, Y => OPEN, FCO => \sum0_5_cry_10\);
    
    \s0[26]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[12]_net_1\, B => \r2[1]_net_1\, C => 
        \r2[29]_net_1\, Y => \s0[26]_net_1\);
    
    \r4[15]\ : SLE
      port map(D => \r5[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[15]_net_1\);
    
    \r9[30]\ : SLE
      port map(D => \r10[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[30]_net_1\);
    
    \s0[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[18]_net_1\, B => \r2[7]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0[0]_net_1\);
    
    \s0[16]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[19]_net_1\, B => \r2[2]_net_1\, C => 
        \r2[23]_net_1\, Y => \s0[16]_net_1\);
    
    \s0[20]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[23]_net_1\, B => \r2[6]_net_1\, C => 
        \r2[27]_net_1\, Y => \s0[20]_net_1\);
    
    \r7[0]\ : SLE
      port map(D => \r8[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[0]_net_1\);
    
    \r2[6]\ : SLE
      port map(D => \r3[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[6]_net_1\);
    
    \s0[10]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[28]_net_1\, B => \r2[13]_net_1\, C => 
        \r2[17]_net_1\, Y => \s0[10]_net_1\);
    
    \r6[11]\ : SLE
      port map(D => \r7[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[11]_net_1\);
    
    sum0_4_axb_6 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[16]_net_1\, B => \s0[6]_net_1\, C => 
        \r15[25]_net_1\, D => \r15[23]_net_1\, Y => 
        \sum0_4_axb_6\);
    
    \r3[26]\ : SLE
      port map(D => \r4[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[26]_net_1\);
    
    \r13[10]\ : SLE
      port map(D => \r14[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[10]_net_1\);
    
    \r12[10]\ : SLE
      port map(D => \r13[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[10]_net_1\);
    
    \r11[28]\ : SLE
      port map(D => \r12[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[28]_net_1\);
    
    \next_r0[8]\ : CFG4
      generic map(INIT => x"888D")

      port map(A => ld_i_i_3, B => next_r0_0_cry_8_S, C => 
        W_out_2_i_2_0, D => W_out_2_i_1_0, Y => \Wt_data[8]\);
    
    \r2[21]\ : SLE
      port map(D => \r3[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[21]_net_1\);
    
    \r3[9]\ : SLE
      port map(D => \r4[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[9]_net_1\);
    
    \r5[20]\ : SLE
      port map(D => \r6[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[20]_net_1\);
    
    \r11[18]\ : SLE
      port map(D => \r12[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[18]_net_1\);
    
    \r0[24]\ : SLE
      port map(D => \Wt_data[24]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[24]_net_1\);
    
    \r13[5]\ : SLE
      port map(D => \r14[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[5]_net_1\);
    
    \r0[14]\ : SLE
      port map(D => \Wt_data[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[14]_net_1\);
    
    sum0_5_cry_13 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[13]_net_1\, B => \r10[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_12\, S => 
        \sum0_5[13]\, Y => OPEN, FCO => \sum0_5_cry_13\);
    
    sum0_4_cry_0_1056 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[18]_net_1\, B => \r2[7]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0_0[0]\);
    
    \r1[2]\ : SLE
      port map(D => \r2[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[2]_net_1\);
    
    \r3[21]\ : SLE
      port map(D => \r4[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[21]_net_1\);
    
    \r11[5]\ : SLE
      port map(D => \r12[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[5]_net_1\);
    
    \r7[15]\ : SLE
      port map(D => \r8[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[15]_net_1\);
    
    sum0_4_cry_22 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[22]\, C => 
        \sum0_4_axb_22\, D => GND_net_1, FCI => \sum0_4_cry_21\, 
        S => \sum0_4[22]\, Y => OPEN, FCO => \sum0_4_cry_22\);
    
    \r1[0]\ : SLE
      port map(D => \r2[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[0]_net_1\);
    
    \r0[1]\ : SLE
      port map(D => \Wt_data[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[1]_net_1\);
    
    \next_r0[5]\ : CFG4
      generic map(INIT => x"CFCA")

      port map(A => N_349, B => next_r0_0_cry_5_S, C => ld_i_i_3, 
        D => W_out_2_0(5), Y => \Wt_data[5]\);
    
    \r14[23]\ : SLE
      port map(D => \r15[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[23]_net_1\);
    
    sum0_5_cry_18 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[18]_net_1\, B => \r10[18]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_17\, S => 
        \sum0_5[18]\, Y => OPEN, FCO => \sum0_5_cry_18\);
    
    \r6[13]\ : SLE
      port map(D => \r7[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[13]_net_1\);
    
    \r1[5]\ : SLE
      port map(D => \r2[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[5]_net_1\);
    
    \r4[12]\ : SLE
      port map(D => \r5[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[12]_net_1\);
    
    \r2[23]\ : SLE
      port map(D => \r3[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[23]_net_1\);
    
    \next_r0[29]\ : CFG4
      generic map(INIT => x"C0C5")

      port map(A => W_out_2_i_1_21, B => next_r0_0_cry_29_S, C
         => ld_i_i_3, D => W_out_2_i_0(29), Y => \Wt_data[29]\);
    
    \r8[24]\ : SLE
      port map(D => \r9[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[24]_net_1\);
    
    \r5[0]\ : SLE
      port map(D => \r6[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[0]_net_1\);
    
    \r6[7]\ : SLE
      port map(D => \r7[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[7]_net_1\);
    
    next_r0_0_cry_13 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[13]\, B => \sum0_5[13]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_12\, S
         => next_r0_0_cry_13_S, Y => OPEN, FCO => 
        \next_r0_0_cry_13\);
    
    \r9[7]\ : SLE
      port map(D => \r10[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[7]_net_1\);
    
    next_r0_0_cry_23 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[23]\, B => \sum0_5[23]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_22\, S
         => next_r0_0_cry_23_S, Y => OPEN, FCO => 
        \next_r0_0_cry_23\);
    
    \r14[29]\ : SLE
      port map(D => \r15[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[29]_net_1\);
    
    \next_r0[1]\ : CFG4
      generic map(INIT => x"C0E2")

      port map(A => N_98, B => ld_i_i_3, C => next_r0_0_cry_1_S, 
        D => W_out_i_0(1), Y => \Wt_data[1]\);
    
    sum0_5_s_31 : ARI1
      generic map(INIT => x"46600")

      port map(A => VCC_net_1, B => \r1[31]_net_1\, C => 
        \r10[31]_net_1\, D => GND_net_1, FCI => \sum0_5_cry_30\, 
        S => \sum0_5[31]\, Y => OPEN, FCO => OPEN);
    
    \r3[1]\ : SLE
      port map(D => \r4[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[1]_net_1\);
    
    \next_r0[6]\ : CFG4
      generic map(INIT => x"CFCA")

      port map(A => N_251, B => next_r0_0_cry_6_S, C => ld_i_i_3, 
        D => W_out_2_0_0_3, Y => \Wt_data[6]\);
    
    \r3[23]\ : SLE
      port map(D => \r4[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[23]_net_1\);
    
    \r11[21]\ : SLE
      port map(D => \r12[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[21]_net_1\);
    
    \r7[27]\ : SLE
      port map(D => \r8[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[27]_net_1\);
    
    \next_r0[22]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_304, C => next_r0_0_cry_22_S, 
        D => W_out_2_i_1_14, Y => \Wt_data[22]\);
    
    \r1[15]\ : SLE
      port map(D => \r2[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[15]_net_1\);
    
    \r11[11]\ : SLE
      port map(D => \r12[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[11]_net_1\);
    
    \r9[4]\ : SLE
      port map(D => \r10[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[4]_net_1\);
    
    \r1[26]\ : SLE
      port map(D => \r2[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[26]_net_1\);
    
    \r5[16]\ : SLE
      port map(D => \r6[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[16]_net_1\);
    
    \r3[31]\ : SLE
      port map(D => \r4[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[31]_net_1\);
    
    \r4[26]\ : SLE
      port map(D => \r5[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[26]_net_1\);
    
    \r7[12]\ : SLE
      port map(D => \r8[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[12]_net_1\);
    
    \next_r0[30]\ : CFG4
      generic map(INIT => x"C0C5")

      port map(A => W_out_2_i_1_22, B => next_r0_0_cry_30_S, C
         => ld_i_i_3, D => W_out_2_i_0(30), Y => \Wt_data[30]\);
    
    \r10[6]\ : SLE
      port map(D => \r11[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[6]_net_1\);
    
    next_r0_0_cry_4 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[4]\, B => \sum0_5[4]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_3\, S => 
        next_r0_0_cry_4_S, Y => OPEN, FCO => \next_r0_0_cry_4\);
    
    \r13[15]\ : SLE
      port map(D => \r14[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[15]_net_1\);
    
    \r12[15]\ : SLE
      port map(D => \r13[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[15]_net_1\);
    
    \r9[5]\ : SLE
      port map(D => \r10[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[5]_net_1\);
    
    \r8[19]\ : SLE
      port map(D => \r9[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[19]_net_1\);
    
    \r6[27]\ : SLE
      port map(D => \r7[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[27]_net_1\);
    
    \r14[24]\ : SLE
      port map(D => \r15[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[24]_net_1\);
    
    \r2[30]\ : SLE
      port map(D => \r3[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[30]_net_1\);
    
    \r14[22]\ : SLE
      port map(D => \r15[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[22]_net_1\);
    
    \r2[4]\ : SLE
      port map(D => \r3[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[4]_net_1\);
    
    \r2[16]\ : SLE
      port map(D => \r3[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[16]_net_1\);
    
    \r1[21]\ : SLE
      port map(D => \r2[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[21]_net_1\);
    
    sum0_4_cry_0_1045 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[29]_net_1\, B => \r2[18]_net_1\, C => 
        \r2[14]_net_1\, Y => \s0_0[11]\);
    
    \r5[11]\ : SLE
      port map(D => \r6[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[11]_net_1\);
    
    \r12[5]\ : SLE
      port map(D => \r13[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[5]_net_1\);
    
    \r15[18]\ : SLE
      port map(D => \r0[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[18]_net_1\);
    
    \r4[21]\ : SLE
      port map(D => \r5[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[21]_net_1\);
    
    \r11[9]\ : SLE
      port map(D => \r12[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[9]_net_1\);
    
    \r15[28]\ : SLE
      port map(D => \r0[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[28]_net_1\);
    
    \r7[5]\ : SLE
      port map(D => \r8[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[5]_net_1\);
    
    \r9[2]\ : SLE
      port map(D => \r10[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[2]_net_1\);
    
    \r4[7]\ : SLE
      port map(D => \r5[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[7]_net_1\);
    
    sum0_4_cry_1 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[1]\, C => 
        \sum0_4_axb_1\, D => GND_net_1, FCI => \sum0_4_cry_0\, S
         => \sum0_4[1]\, Y => OPEN, FCO => \sum0_4_cry_1\);
    
    sum0_4_cry_15 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[15]\, C => 
        \sum0_4_axb_15\, D => GND_net_1, FCI => \sum0_4_cry_14\, 
        S => \sum0_4[15]\, Y => OPEN, FCO => \sum0_4_cry_15\);
    
    \r7[28]\ : SLE
      port map(D => \r8[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[28]_net_1\);
    
    sum0_5_cry_20 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[20]_net_1\, B => \r10[20]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_19\, S => 
        \sum0_5[20]\, Y => OPEN, FCO => \sum0_5_cry_20\);
    
    \r1[12]\ : SLE
      port map(D => \r2[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[12]_net_1\);
    
    \next_r0[3]\ : CFG4
      generic map(INIT => x"CFCA")

      port map(A => N_245, B => next_r0_0_cry_3_S, C => ld_i_i_3, 
        D => W_out_2_0_0_0, Y => \Wt_data[3]\);
    
    \r8[4]\ : SLE
      port map(D => \r9[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[4]_net_1\);
    
    \r2[11]\ : SLE
      port map(D => \r3[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[11]_net_1\);
    
    sum0_5_cry_19 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[19]_net_1\, B => \r10[19]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_18\, S => 
        \sum0_5[19]\, Y => OPEN, FCO => \sum0_5_cry_19\);
    
    \r7[4]\ : SLE
      port map(D => \r8[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[4]_net_1\);
    
    \r6[6]\ : SLE
      port map(D => \r7[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[6]_net_1\);
    
    \r9[26]\ : SLE
      port map(D => \r10[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[26]_net_1\);
    
    \r10[9]\ : SLE
      port map(D => \r11[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[9]_net_1\);
    
    sum0_4_cry_7 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[7]\, C => 
        \sum0_4_axb_7\, D => GND_net_1, FCI => \sum0_4_cry_6\, S
         => \sum0_4[7]\, Y => OPEN, FCO => \sum0_4_cry_7\);
    
    \r4[3]\ : SLE
      port map(D => \r5[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[3]_net_1\);
    
    \r1[23]\ : SLE
      port map(D => \r2[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[23]_net_1\);
    
    sum0_5_cry_16 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[16]_net_1\, B => \r10[16]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_15\, S => 
        \sum0_5[16]\, Y => OPEN, FCO => \sum0_5_cry_16\);
    
    \r5[13]\ : SLE
      port map(D => \r6[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[13]_net_1\);
    
    \s0[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[27]_net_1\, B => \r2[16]_net_1\, C => 
        \r2[12]_net_1\, Y => \s0[9]_net_1\);
    
    \r4[23]\ : SLE
      port map(D => \r5[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[23]_net_1\);
    
    \r14[3]\ : SLE
      port map(D => \r15[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[3]_net_1\);
    
    next_r0_0_cry_5 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[5]\, B => \sum0_5[5]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_4\, S => 
        next_r0_0_cry_5_S, Y => OPEN, FCO => \next_r0_0_cry_5\);
    
    \s0[21]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[28]_net_1\, B => \r2[24]_net_1\, C => 
        \r2[7]_net_1\, Y => \s0[21]_net_1\);
    
    \r6[28]\ : SLE
      port map(D => \r7[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[28]_net_1\);
    
    \r6[17]\ : SLE
      port map(D => \r7[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[17]_net_1\);
    
    \r5[29]\ : SLE
      port map(D => \r6[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[29]_net_1\);
    
    \next_r0[19]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_295, C => next_r0_0_cry_19_S, 
        D => W_out_2_i_1_11, Y => \Wt_data[19]\);
    
    sum0_4_cry_0_1035 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[28]_net_1\, B => \r2[24]_net_1\, C => 
        \r2[7]_net_1\, Y => \s0_0[21]\);
    
    \s0[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[29]_net_1\, B => \r2[18]_net_1\, C => 
        \r2[14]_net_1\, Y => \s0[11]_net_1\);
    
    sum0_4_axb_18 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[3]_net_1\, B => \r15[5]_net_1\, C => 
        \s0[18]_net_1\, D => \r15[28]_net_1\, Y => 
        \sum0_4_axb_18\);
    
    \r5[7]\ : SLE
      port map(D => \r6[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[7]_net_1\);
    
    sum0_4_cry_0_1053 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[10]_net_1\, B => \r2[6]_net_1\, C => 
        \r2[21]_net_1\, Y => \s0_0[3]\);
    
    \r2[27]\ : SLE
      port map(D => \r3[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[27]_net_1\);
    
    sum0_5_cry_23 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[23]_net_1\, B => \r10[23]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_22\, S => 
        \sum0_5[23]\, Y => OPEN, FCO => \sum0_5_cry_23\);
    
    \r4[31]\ : SLE
      port map(D => \r5[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[31]_net_1\);
    
    \r2[8]\ : SLE
      port map(D => \r3[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[8]_net_1\);
    
    \r2[3]\ : SLE
      port map(D => \r3[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[3]_net_1\);
    
    \r9[21]\ : SLE
      port map(D => \r10[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[21]_net_1\);
    
    \r2[13]\ : SLE
      port map(D => \r3[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[13]_net_1\);
    
    \r13[17]\ : SLE
      port map(D => \r14[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[17]_net_1\);
    
    \r12[17]\ : SLE
      port map(D => \r13[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[17]_net_1\);
    
    \r15[11]\ : SLE
      port map(D => \r0[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[11]_net_1\);
    
    \r9[10]\ : SLE
      port map(D => \r10[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[10]_net_1\);
    
    \r14[26]\ : SLE
      port map(D => \r15[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[26]_net_1\);
    
    \s0[23]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[30]_net_1\, B => \r2[26]_net_1\, C => 
        \r2[9]_net_1\, Y => \s0[23]_net_1\);
    
    sum0_4_s_31 : ARI1
      generic map(INIT => x"46996")

      port map(A => \r15[18]_net_1\, B => \r2[6]_net_1\, C => 
        \r2[17]_net_1\, D => \r15[16]_net_1\, FCI => 
        \sum0_4_cry_30\, S => \sum0_4[31]\, Y => OPEN, FCO => 
        OPEN);
    
    \r13[2]\ : SLE
      port map(D => \r14[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[2]_net_1\);
    
    sum0_5_cry_28 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[28]_net_1\, B => \r10[28]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_27\, S => 
        \sum0_5[28]\, Y => OPEN, FCO => \sum0_5_cry_28\);
    
    \r14[9]\ : SLE
      port map(D => \r15[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[9]_net_1\);
    
    \s0[13]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[20]_net_1\, C => 
        \r2[16]_net_1\, Y => \s0[13]_net_1\);
    
    \r3[27]\ : SLE
      port map(D => \r4[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[27]_net_1\);
    
    \next_r0[12]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_272, C => next_r0_0_cry_12_S, 
        D => W_out_2_i_1_4, Y => \Wt_data[12]\);
    
    \r15[21]\ : SLE
      port map(D => \r0[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[21]_net_1\);
    
    sum0_4_cry_6 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[6]\, C => 
        \sum0_4_axb_6\, D => GND_net_1, FCI => \sum0_4_cry_5\, S
         => \sum0_4[6]\, Y => OPEN, FCO => \sum0_4_cry_6\);
    
    \r13[6]\ : SLE
      port map(D => \r14[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[6]_net_1\);
    
    \r6[5]\ : SLE
      port map(D => \r7[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[5]_net_1\);
    
    \r3[10]\ : SLE
      port map(D => \r4[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[10]_net_1\);
    
    \r3[7]\ : SLE
      port map(D => \r4[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[7]_net_1\);
    
    \r11[3]\ : SLE
      port map(D => \r12[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[3]_net_1\);
    
    sum0_5_cry_12 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[12]_net_1\, B => \r10[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_11\, S => 
        \sum0_5[12]\, Y => OPEN, FCO => \sum0_5_cry_12\);
    
    \r14[18]\ : SLE
      port map(D => \r15[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[18]_net_1\);
    
    \r9[3]\ : SLE
      port map(D => \r10[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[3]_net_1\);
    
    \r14[5]\ : SLE
      port map(D => \r15[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[5]_net_1\);
    
    \r12[20]\ : SLE
      port map(D => \r13[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[20]_net_1\);
    
    \r10[20]\ : SLE
      port map(D => \r11[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[20]_net_1\);
    
    \r9[23]\ : SLE
      port map(D => \r10[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[23]_net_1\);
    
    \r0[26]\ : SLE
      port map(D => \Wt_data[26]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[26]_net_1\);
    
    sum0_4_cry_0_1052 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[22]_net_1\, B => \r2[11]_net_1\, C => 
        \r2[7]_net_1\, Y => \s0_0[4]\);
    
    \r15[2]\ : SLE
      port map(D => \r0[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[2]_net_1\);
    
    \r6[18]\ : SLE
      port map(D => \r7[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[18]_net_1\);
    
    \r0[16]\ : SLE
      port map(D => \Wt_data[16]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[16]_net_1\);
    
    \r2[28]\ : SLE
      port map(D => \r3[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[28]_net_1\);
    
    \r6[30]\ : SLE
      port map(D => \r7[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[30]_net_1\);
    
    \r12[8]\ : SLE
      port map(D => \r13[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[8]_net_1\);
    
    sum0_4_cry_27 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[27]\, C => 
        \sum0_4_axb_27\, D => GND_net_1, FCI => \sum0_4_cry_26\, 
        S => \sum0_4[27]\, Y => OPEN, FCO => \sum0_4_cry_27\);
    
    sum0_4_axb_26 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[11]_net_1\, B => \s0[26]_net_1\, C => 
        \r15[13]_net_1\, Y => \sum0_4_axb_26\);
    
    \r1[1]\ : SLE
      port map(D => \r2[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[1]_net_1\);
    
    sum0_4_cry_4 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[4]\, C => 
        \sum0_4_axb_4\, D => GND_net_1, FCI => \sum0_4_cry_3\, S
         => \sum0_4[4]\, Y => OPEN, FCO => \sum0_4_cry_4\);
    
    \r7[25]\ : SLE
      port map(D => \r8[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[25]_net_1\);
    
    \r0[21]\ : SLE
      port map(D => \Wt_data[21]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[21]_net_1\);
    
    \r1[4]\ : SLE
      port map(D => \r2[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[4]_net_1\);
    
    \r15[30]\ : SLE
      port map(D => \r0[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[30]_net_1\);
    
    sum0_4_axb_29 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[14]_net_1\, B => \s0[29]_net_1\, C => 
        \r15[16]_net_1\, Y => \sum0_4_axb_29\);
    
    \r13[4]\ : SLE
      port map(D => \r14[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[4]_net_1\);
    
    sum0_4_cry_0_1046 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[28]_net_1\, B => \r2[13]_net_1\, C => 
        \r2[17]_net_1\, Y => \s0_0[10]\);
    
    \r8[14]\ : SLE
      port map(D => \r9[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[14]_net_1\);
    
    \r0[11]\ : SLE
      port map(D => \Wt_data[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[11]_net_1\);
    
    \r3[28]\ : SLE
      port map(D => \r4[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[28]_net_1\);
    
    \r8[26]\ : SLE
      port map(D => \r9[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[26]_net_1\);
    
    sum0_4_cry_8 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[8]\, C => 
        \sum0_4_axb_8\, D => GND_net_1, FCI => \sum0_4_cry_7\, S
         => \sum0_4[8]\, Y => OPEN, FCO => \sum0_4_cry_8\);
    
    \r12[2]\ : SLE
      port map(D => \r13[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[2]_net_1\);
    
    \r10[2]\ : SLE
      port map(D => \r11[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[2]_net_1\);
    
    sum0_4_cry_3 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[3]\, C => 
        \sum0_4_axb_3\, D => GND_net_1, FCI => \sum0_4_cry_2\, S
         => \sum0_4[3]\, Y => OPEN, FCO => \sum0_4_cry_3\);
    
    \r7[9]\ : SLE
      port map(D => \r8[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[9]_net_1\);
    
    \r10[10]\ : SLE
      port map(D => \r11[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[10]_net_1\);
    
    \r10[8]\ : SLE
      port map(D => \r11[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[8]_net_1\);
    
    \r6[25]\ : SLE
      port map(D => \r7[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[25]_net_1\);
    
    \r4[10]\ : SLE
      port map(D => \r5[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[10]_net_1\);
    
    \r1[27]\ : SLE
      port map(D => \r2[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[27]_net_1\);
    
    \r14[31]\ : SLE
      port map(D => \r15[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[31]_net_1\);
    
    \r14[11]\ : SLE
      port map(D => \r15[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[11]_net_1\);
    
    \r5[17]\ : SLE
      port map(D => \r6[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[17]_net_1\);
    
    \r4[27]\ : SLE
      port map(D => \r5[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[27]_net_1\);
    
    \r13[13]\ : SLE
      port map(D => \r14[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[13]_net_1\);
    
    \r12[13]\ : SLE
      port map(D => \r13[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[13]_net_1\);
    
    next_r0_0_cry_14 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[14]\, B => \sum0_5[14]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_13\, S
         => next_r0_0_cry_14_S, Y => OPEN, FCO => 
        \next_r0_0_cry_14\);
    
    sum0_4_axb_21 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[6]_net_1\, B => \r15[8]_net_1\, C => 
        \s0[21]_net_1\, D => \r15[31]_net_1\, Y => 
        \sum0_4_axb_21\);
    
    \r8[21]\ : SLE
      port map(D => \r9[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[21]_net_1\);
    
    \r0[23]\ : SLE
      port map(D => \Wt_data[23]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[23]_net_1\);
    
    next_r0_0_cry_24 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[24]\, B => \sum0_5[24]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_23\, S
         => next_r0_0_cry_24_S, Y => OPEN, FCO => 
        \next_r0_0_cry_24\);
    
    \r14[4]\ : SLE
      port map(D => \r15[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[4]_net_1\);
    
    sum0_5_cry_29 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[29]_net_1\, B => \r10[29]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_28\, S => 
        \sum0_5[29]\, Y => OPEN, FCO => \sum0_5_cry_29\);
    
    \r0[13]\ : SLE
      port map(D => \Wt_data[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[13]_net_1\);
    
    \r13[20]\ : SLE
      port map(D => \r14[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[20]_net_1\);
    
    sum0_4_cry_0_1036 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[23]_net_1\, B => \r2[6]_net_1\, C => 
        \r2[27]_net_1\, Y => \s0_0[20]\);
    
    \r13[1]\ : SLE
      port map(D => \r14[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[1]_net_1\);
    
    \r12[25]\ : SLE
      port map(D => \r13[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[25]_net_1\);
    
    \r10[25]\ : SLE
      port map(D => \r11[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[25]_net_1\);
    
    \r2[17]\ : SLE
      port map(D => \r3[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[17]_net_1\);
    
    sum0_5_cry_26 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[26]_net_1\, B => \r10[26]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_25\, S => 
        \sum0_5[26]\, Y => OPEN, FCO => \sum0_5_cry_26\);
    
    \r7[22]\ : SLE
      port map(D => \r8[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[22]_net_1\);
    
    \r14[1]\ : SLE
      port map(D => \r15[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[1]_net_1\);
    
    \r8[6]\ : SLE
      port map(D => \r9[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[6]_net_1\);
    
    \r1[30]\ : SLE
      port map(D => \r2[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[30]_net_1\);
    
    \r15[9]\ : SLE
      port map(D => \r0[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[9]_net_1\);
    
    \r13[19]\ : SLE
      port map(D => \r14[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[19]_net_1\);
    
    \r12[19]\ : SLE
      port map(D => \r13[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[19]_net_1\);
    
    sum0_4_axb_30 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[15]_net_1\, B => \s0[30]_net_1\, C => 
        \r15[17]_net_1\, Y => \sum0_4_axb_30\);
    
    \r2[0]\ : SLE
      port map(D => \r3[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[0]_net_1\);
    
    \r5[24]\ : SLE
      port map(D => \r6[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[24]_net_1\);
    
    sum0_4_cry_0_1054 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[20]_net_1\, B => \r2[9]_net_1\, C => 
        \r2[5]_net_1\, Y => \s0_0[2]\);
    
    \r7[31]\ : SLE
      port map(D => \r8[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[31]_net_1\);
    
    sum0_5_cry_7 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[7]_net_1\, B => \r10[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_6\, S => 
        \sum0_5[7]\, Y => OPEN, FCO => \sum0_5_cry_7\);
    
    \r7[10]\ : SLE
      port map(D => \r8[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[10]_net_1\);
    
    \s0[3]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[10]_net_1\, B => \r2[6]_net_1\, C => 
        \r2[21]_net_1\, Y => \s0[3]_net_1\);
    
    \next_r0[31]\ : CFG4
      generic map(INIT => x"AFAC")

      port map(A => next_r0_0_s_31_S, B => W_out_i_i_1_1(31), C
         => ld_i_i_3, D => W_out_i_i_1(31), Y => \Wt_data[31]\);
    
    sum0_4_cry_24 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[24]\, C => 
        \sum0_4_axb_24\, D => GND_net_1, FCI => \sum0_4_cry_23\, 
        S => \sum0_4[24]\, Y => OPEN, FCO => \sum0_4_cry_24\);
    
    \r4[0]\ : SLE
      port map(D => \r5[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[0]_net_1\);
    
    \r15[8]\ : SLE
      port map(D => \r0[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[8]_net_1\);
    
    \r8[23]\ : SLE
      port map(D => \r9[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[23]_net_1\);
    
    sum0_4_axb_22 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[7]_net_1\, B => \s0[22]_net_1\, C => 
        \r15[9]_net_1\, Y => \sum0_4_axb_22\);
    
    \r10[31]\ : SLE
      port map(D => \r11[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[31]_net_1\);
    
    \r6[22]\ : SLE
      port map(D => \r7[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[22]_net_1\);
    
    \r10[5]\ : SLE
      port map(D => \r11[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[5]_net_1\);
    
    \r1[28]\ : SLE
      port map(D => \r2[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[28]_net_1\);
    
    \r6[15]\ : SLE
      port map(D => \r7[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[15]_net_1\);
    
    \r5[18]\ : SLE
      port map(D => \r6[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[18]_net_1\);
    
    \s0[7]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[25]_net_1\, B => \r2[14]_net_1\, C => 
        \r2[10]_net_1\, Y => \s0[7]_net_1\);
    
    \r0[2]\ : SLE
      port map(D => \Wt_data[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[2]_net_1\);
    
    \r4[28]\ : SLE
      port map(D => \r5[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[28]_net_1\);
    
    \r2[25]\ : SLE
      port map(D => \r3[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[25]_net_1\);
    
    \r11[6]\ : SLE
      port map(D => \r12[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[6]_net_1\);
    
    \r9[27]\ : SLE
      port map(D => \r10[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[27]_net_1\);
    
    sum0_4_axb_25 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[10]_net_1\, B => \s0[25]_net_1\, C => 
        \r15[12]_net_1\, Y => \sum0_4_axb_25\);
    
    \r9[19]\ : SLE
      port map(D => \r10[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[19]_net_1\);
    
    \r12[31]\ : SLE
      port map(D => \r13[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[31]_net_1\);
    
    \r13[14]\ : SLE
      port map(D => \r14[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[14]_net_1\);
    
    \r12[14]\ : SLE
      port map(D => \r13[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[14]_net_1\);
    
    next_r0_0_cry_1 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[1]\, B => \sum0_5[1]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_0\, S => 
        next_r0_0_cry_1_S, Y => OPEN, FCO => \next_r0_0_cry_1\);
    
    next_r0_0_cry_19 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[19]\, B => \sum0_5[19]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_18\, S
         => next_r0_0_cry_19_S, Y => OPEN, FCO => 
        \next_r0_0_cry_19\);
    
    \r13[12]\ : SLE
      port map(D => \r14[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[12]_net_1\);
    
    \r12[12]\ : SLE
      port map(D => \r13[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[12]_net_1\);
    
    next_r0_0_cry_2 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[2]\, B => \sum0_5[2]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_1\, S => 
        next_r0_0_cry_2_S, Y => OPEN, FCO => \next_r0_0_cry_2\);
    
    sum0_5_cry_22 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[22]_net_1\, B => \r10[22]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_21\, S => 
        \sum0_5[22]\, Y => OPEN, FCO => \sum0_5_cry_22\);
    
    \r3[19]\ : SLE
      port map(D => \r4[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[19]_net_1\);
    
    next_r0_0_cry_29 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[29]\, B => \sum0_5[29]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_28\, S
         => next_r0_0_cry_29_S, Y => OPEN, FCO => 
        \next_r0_0_cry_29\);
    
    \r10[15]\ : SLE
      port map(D => \r11[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[15]_net_1\);
    
    \r2[18]\ : SLE
      port map(D => \r3[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[18]_net_1\);
    
    \r3[25]\ : SLE
      port map(D => \r4[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[25]_net_1\);
    
    \r1[10]\ : SLE
      port map(D => \r2[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[10]_net_1\);
    
    sum0_5_cry_0 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[0]_net_1\, B => \r10[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => GND_net_1, S => OPEN, Y
         => sum0_5_cry_0_Y, FCO => \sum0_5_cry_0\);
    
    \s0[27]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[13]_net_1\, B => \r2[2]_net_1\, C => 
        \r2[30]_net_1\, Y => \s0[27]_net_1\);
    
    \r14[0]\ : SLE
      port map(D => \r15[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[0]_net_1\);
    
    \next_r0[20]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_298, C => next_r0_0_cry_20_S, 
        D => W_out_2_i_1_12, Y => \Wt_data[20]\);
    
    sum0_4_cry_0_1026 : CFG2
      generic map(INIT => x"6")

      port map(A => \r2[5]_net_1\, B => \r2[16]_net_1\, Y => 
        \s0_0[30]\);
    
    \s0[17]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[24]_net_1\, B => \r2[20]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0[17]_net_1\);
    
    \r13[25]\ : SLE
      port map(D => \r14[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[25]_net_1\);
    
    \r8[0]\ : SLE
      port map(D => \r9[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[0]_net_1\);
    
    \r12[27]\ : SLE
      port map(D => \r13[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[27]_net_1\);
    
    \r10[27]\ : SLE
      port map(D => \r11[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[27]_net_1\);
    
    \r6[12]\ : SLE
      port map(D => \r7[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[12]_net_1\);
    
    \r3[5]\ : SLE
      port map(D => \r4[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[5]_net_1\);
    
    \r0[30]\ : SLE
      port map(D => \Wt_data[30]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[30]_net_1\);
    
    sum0_4_cry_0_1043 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[20]_net_1\, C => 
        \r2[16]_net_1\, Y => \s0_0[13]\);
    
    \r2[22]\ : SLE
      port map(D => \r3[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[22]_net_1\);
    
    \r9[28]\ : SLE
      port map(D => \r10[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[28]_net_1\);
    
    \r11[1]\ : SLE
      port map(D => \r12[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[1]_net_1\);
    
    sum0_5_cry_17 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[17]_net_1\, B => \r10[17]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_16\, S => 
        \sum0_5[17]\, Y => OPEN, FCO => \sum0_5_cry_17\);
    
    next_r0_0_cry_8 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[8]\, B => \sum0_5[8]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_7\, S => 
        next_r0_0_cry_8_S, Y => OPEN, FCO => \next_r0_0_cry_8\);
    
    \r0[27]\ : SLE
      port map(D => \Wt_data[27]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[27]_net_1\);
    
    next_r0_0_cry_6 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[6]\, B => \sum0_5[6]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_5\, S => 
        next_r0_0_cry_6_S, Y => OPEN, FCO => \next_r0_0_cry_6\);
    
    \r0[17]\ : SLE
      port map(D => \Wt_data[17]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[17]_net_1\);
    
    \r15[4]\ : SLE
      port map(D => \r0[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[4]_net_1\);
    
    \r14[8]\ : SLE
      port map(D => \r15[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[8]_net_1\);
    
    \r14[28]\ : SLE
      port map(D => \r15[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[28]_net_1\);
    
    \r12[7]\ : SLE
      port map(D => \r13[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[7]_net_1\);
    
    sum0_4_cry_0_1048 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[26]_net_1\, B => \r2[15]_net_1\, C => 
        \r2[11]_net_1\, Y => \s0_0[8]\);
    
    next_r0_0_cry_3 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[3]\, B => \sum0_5[3]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_2\, S => 
        next_r0_0_cry_3_S, Y => OPEN, FCO => \next_r0_0_cry_3\);
    
    \r3[22]\ : SLE
      port map(D => \r4[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[22]_net_1\);
    
    \r8[2]\ : SLE
      port map(D => \r9[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[2]_net_1\);
    
    \s0[28]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[14]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0[28]_net_1\);
    
    \s0[18]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[25]_net_1\, B => \r2[21]_net_1\, C => 
        \r2[4]_net_1\, Y => \s0[18]_net_1\);
    
    \r4[19]\ : SLE
      port map(D => \r5[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[19]_net_1\);
    
    sum0_4_cry_11 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[11]\, C => 
        \sum0_4_axb_11\, D => GND_net_1, FCI => \sum0_4_cry_10\, 
        S => \sum0_4[11]\, Y => OPEN, FCO => \sum0_4_cry_11\);
    
    \r13[16]\ : SLE
      port map(D => \r14[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[16]_net_1\);
    
    \r12[16]\ : SLE
      port map(D => \r13[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[16]_net_1\);
    
    \r5[30]\ : SLE
      port map(D => \r6[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[30]_net_1\);
    
    \r7[7]\ : SLE
      port map(D => \r8[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[7]_net_1\);
    
    sum0_4_axb_3 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[13]_net_1\, B => \s0[3]_net_1\, C => 
        \r15[22]_net_1\, D => \r15[20]_net_1\, Y => 
        \sum0_4_axb_3\);
    
    \r1[25]\ : SLE
      port map(D => \r2[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[25]_net_1\);
    
    \r5[15]\ : SLE
      port map(D => \r6[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[15]_net_1\);
    
    sum0_4_cry_0_1042 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[0]_net_1\, B => \r2[17]_net_1\, C => 
        \r2[21]_net_1\, Y => \s0_0[14]\);
    
    sum0_4_cry_0_1033 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[30]_net_1\, B => \r2[26]_net_1\, C => 
        \r2[9]_net_1\, Y => \s0_0[23]\);
    
    \r8[27]\ : SLE
      port map(D => \r9[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[27]_net_1\);
    
    \r10[17]\ : SLE
      port map(D => \r11[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[17]_net_1\);
    
    next_r0_0_cry_9 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[9]\, B => \sum0_5[9]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_8\, S => 
        next_r0_0_cry_9_S, Y => OPEN, FCO => \next_r0_0_cry_9\);
    
    \r4[25]\ : SLE
      port map(D => \r5[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[25]_net_1\);
    
    \r1[9]\ : SLE
      port map(D => \r2[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[9]_net_1\);
    
    \r8[16]\ : SLE
      port map(D => \r9[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[16]_net_1\);
    
    sum0_4_axb_16 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[1]_net_1\, B => \r15[3]_net_1\, C => 
        \s0[16]_net_1\, D => \r15[26]_net_1\, Y => 
        \sum0_4_axb_16\);
    
    \r10[1]\ : SLE
      port map(D => \r11[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[1]_net_1\);
    
    \s0[29]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \r2[4]_net_1\, B => \r2[15]_net_1\, Y => 
        \s0[29]_net_1\);
    
    \r0[28]\ : SLE
      port map(D => \Wt_data[28]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[28]_net_1\);
    
    \r9[6]\ : SLE
      port map(D => \r10[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[6]_net_1\);
    
    \s0[19]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[26]_net_1\, B => \r2[22]_net_1\, C => 
        \r2[5]_net_1\, Y => \s0[19]_net_1\);
    
    sum0_4_axb_19 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[4]_net_1\, B => \r15[6]_net_1\, C => 
        \s0[19]_net_1\, D => \r15[29]_net_1\, Y => 
        \sum0_4_axb_19\);
    
    sum0_4_cry_0_1038 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[25]_net_1\, B => \r2[21]_net_1\, C => 
        \r2[4]_net_1\, Y => \s0_0[18]\);
    
    \r0[18]\ : SLE
      port map(D => \Wt_data[18]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[18]_net_1\);
    
    \r2[15]\ : SLE
      port map(D => \r3[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[15]_net_1\);
    
    \r7[19]\ : SLE
      port map(D => \r8[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[19]_net_1\);
    
    \r13[27]\ : SLE
      port map(D => \r14[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[27]_net_1\);
    
    \r9[8]\ : SLE
      port map(D => \r10[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[8]_net_1\);
    
    \r8[11]\ : SLE
      port map(D => \r9[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[11]_net_1\);
    
    \r14[21]\ : SLE
      port map(D => \r15[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[21]_net_1\);
    
    \r12[23]\ : SLE
      port map(D => \r13[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[23]_net_1\);
    
    \r10[23]\ : SLE
      port map(D => \r11[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[23]_net_1\);
    
    \r9[14]\ : SLE
      port map(D => \r10[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[14]_net_1\);
    
    sum0_5_cry_14 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[14]_net_1\, B => \r10[14]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_13\, S => 
        \sum0_5[14]\, Y => OPEN, FCO => \sum0_5_cry_14\);
    
    \next_r0[10]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_265, C => next_r0_0_cry_10_S, 
        D => W_out_2_i_1_2, Y => \Wt_data[10]\);
    
    sum0_4_cry_0_1032 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[27]_net_1\, C => 
        \r2[10]_net_1\, Y => \s0_0[24]\);
    
    sum0_4_axb_8 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[18]_net_1\, B => \s0[8]_net_1\, C => 
        \r15[27]_net_1\, D => \r15[25]_net_1\, Y => 
        \sum0_4_axb_8\);
    
    \r1[22]\ : SLE
      port map(D => \r2[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[22]_net_1\);
    
    \r11[20]\ : SLE
      port map(D => \r12[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[20]_net_1\);
    
    \r5[12]\ : SLE
      port map(D => \r6[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[12]_net_1\);
    
    \r3[14]\ : SLE
      port map(D => \r4[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[14]_net_1\);
    
    \r8[28]\ : SLE
      port map(D => \r9[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[28]_net_1\);
    
    \r5[6]\ : SLE
      port map(D => \r6[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[6]_net_1\);
    
    sum0_4_axb_11 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[21]_net_1\, B => \s0[11]_net_1\, C => 
        \r15[30]_net_1\, D => \r15[28]_net_1\, Y => 
        \sum0_4_axb_11\);
    
    sum0_4_cry_2 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[2]\, C => 
        \sum0_4_axb_2\, D => GND_net_1, FCI => \sum0_4_cry_1\, S
         => \sum0_4[2]\, Y => OPEN, FCO => \sum0_4_cry_2\);
    
    \r11[10]\ : SLE
      port map(D => \r12[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[10]_net_1\);
    
    sum0_4_cry_25 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[25]\, C => 
        \sum0_4_axb_25\, D => GND_net_1, FCI => \sum0_4_cry_24\, 
        S => \sum0_4[25]\, Y => OPEN, FCO => \sum0_4_cry_25\);
    
    \r4[22]\ : SLE
      port map(D => \r5[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[22]_net_1\);
    
    \r9[25]\ : SLE
      port map(D => \r10[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[25]_net_1\);
    
    \next_r0[26]\ : CFG4
      generic map(INIT => x"C0C5")

      port map(A => W_out_2_i_1_18, B => next_r0_0_cry_26_S, C
         => ld_i_i_3, D => W_out_2_i_0(26), Y => \Wt_data[26]\);
    
    \r12[29]\ : SLE
      port map(D => \r13[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[29]_net_1\);
    
    \r10[29]\ : SLE
      port map(D => \r11[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[29]_net_1\);
    
    \r5[26]\ : SLE
      port map(D => \r6[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[26]_net_1\);
    
    \r1[19]\ : SLE
      port map(D => \r2[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[19]_net_1\);
    
    sum0_4_axb_23 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[8]_net_1\, B => \r15[10]_net_1\, C => 
        \s0[23]_net_1\, Y => \sum0_4_axb_23\);
    
    \r8[5]\ : SLE
      port map(D => \r9[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[5]_net_1\);
    
    sum0_4_axb_5 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[15]_net_1\, B => \s0[5]_net_1\, C => 
        \r15[24]_net_1\, D => \r15[22]_net_1\, Y => 
        \sum0_4_axb_5\);
    
    \r8[13]\ : SLE
      port map(D => \r9[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[13]_net_1\);
    
    \r9[31]\ : SLE
      port map(D => \r10[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[31]_net_1\);
    
    \r0[4]\ : SLE
      port map(D => \Wt_data[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[4]_net_1\);
    
    sum0_4_axb_20 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[5]_net_1\, B => \r15[7]_net_1\, C => 
        \s0[20]_net_1\, D => \r15[30]_net_1\, Y => 
        \sum0_4_axb_20\);
    
    \r7[20]\ : SLE
      port map(D => \r8[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[20]_net_1\);
    
    \r2[12]\ : SLE
      port map(D => \r3[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[12]_net_1\);
    
    \r15[0]\ : SLE
      port map(D => \r0[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[0]_net_1\);
    
    \r1[6]\ : SLE
      port map(D => \r2[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[6]_net_1\);
    
    \s0[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[19]_net_1\, B => \r2[8]_net_1\, C => 
        \r2[4]_net_1\, Y => \s0[1]_net_1\);
    
    \r0[5]\ : SLE
      port map(D => \Wt_data[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[5]_net_1\);
    
    sum0_4_cry_0_1044 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[30]_net_1\, B => \r2[19]_net_1\, C => 
        \r2[15]_net_1\, Y => \s0_0[12]\);
    
    \r15[6]\ : SLE
      port map(D => \r0[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[6]_net_1\);
    
    \r6[4]\ : SLE
      port map(D => \r7[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[4]_net_1\);
    
    \r5[21]\ : SLE
      port map(D => \r6[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[21]_net_1\);
    
    \r10[13]\ : SLE
      port map(D => \r11[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[13]_net_1\);
    
    \r0[6]\ : SLE
      port map(D => \Wt_data[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[6]_net_1\);
    
    sum0_4_cry_0_1028 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[14]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0_0[28]\);
    
    sum0_4_axb_12 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[22]_net_1\, B => \s0[12]_net_1\, C => 
        \r15[31]_net_1\, D => \r15[29]_net_1\, Y => 
        \sum0_4_axb_12\);
    
    \r4[2]\ : SLE
      port map(D => \r5[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[2]_net_1\);
    
    \r12[24]\ : SLE
      port map(D => \r13[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[24]_net_1\);
    
    \r10[24]\ : SLE
      port map(D => \r11[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[24]_net_1\);
    
    sum0_5_cry_27 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[27]_net_1\, B => \r10[27]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_26\, S => 
        \sum0_5[27]\, Y => OPEN, FCO => \sum0_5_cry_27\);
    
    \r6[20]\ : SLE
      port map(D => \r7[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[20]_net_1\);
    
    \r12[22]\ : SLE
      port map(D => \r13[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[22]_net_1\);
    
    \r10[22]\ : SLE
      port map(D => \r11[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[22]_net_1\);
    
    \r8[30]\ : SLE
      port map(D => \r9[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[30]_net_1\);
    
    \r3[6]\ : SLE
      port map(D => \r4[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[6]_net_1\);
    
    sum0_4_axb_15 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[0]_net_1\, B => \r15[2]_net_1\, C => 
        \s0[15]_net_1\, D => \r15[25]_net_1\, Y => 
        \sum0_4_axb_15\);
    
    sum0_4_axb_9 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[19]_net_1\, B => \s0[9]_net_1\, C => 
        \r15[28]_net_1\, D => \r15[26]_net_1\, Y => 
        \sum0_4_axb_9\);
    
    \r9[22]\ : SLE
      port map(D => \r10[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[22]_net_1\);
    
    \r13[23]\ : SLE
      port map(D => \r14[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[23]_net_1\);
    
    \r10[19]\ : SLE
      port map(D => \r11[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[19]_net_1\);
    
    \r0[25]\ : SLE
      port map(D => \Wt_data[25]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[25]_net_1\);
    
    sum0_4_cry_5 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[5]\, C => 
        \sum0_4_axb_5\, D => GND_net_1, FCI => \sum0_4_cry_4\, S
         => \sum0_4[5]\, Y => OPEN, FCO => \sum0_4_cry_5\);
    
    \r4[14]\ : SLE
      port map(D => \r5[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[14]_net_1\);
    
    \r0[15]\ : SLE
      port map(D => \Wt_data[15]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[15]_net_1\);
    
    \r5[23]\ : SLE
      port map(D => \r6[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[23]_net_1\);
    
    \r13[9]\ : SLE
      port map(D => \r14[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[9]_net_1\);
    
    \r11[25]\ : SLE
      port map(D => \r12[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[25]_net_1\);
    
    sum0_4_cry_10 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[10]\, C => 
        \sum0_4_axb_10\, D => GND_net_1, FCI => \sum0_4_cry_9\, S
         => \sum0_4[10]\, Y => OPEN, FCO => \sum0_4_cry_10\);
    
    sum0_4_cry_0_1034 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[29]_net_1\, B => \r2[25]_net_1\, C => 
        \r2[8]_net_1\, Y => \s0_0[22]\);
    
    next_r0_0_cry_7 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[7]\, B => \sum0_5[7]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_6\, S => 
        next_r0_0_cry_7_S, Y => OPEN, FCO => \next_r0_0_cry_7\);
    
    \r11[15]\ : SLE
      port map(D => \r12[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[15]_net_1\);
    
    sum0_4_cry_0_1049 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[25]_net_1\, B => \r2[14]_net_1\, C => 
        \r2[10]_net_1\, Y => \s0_0[7]\);
    
    \r13[29]\ : SLE
      port map(D => \r14[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[29]_net_1\);
    
    sum0_5_cry_3 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[3]_net_1\, B => \r10[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_2\, S => 
        \sum0_5[3]\, Y => OPEN, FCO => \sum0_5_cry_3\);
    
    \r0[8]\ : SLE
      port map(D => \Wt_data[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[8]_net_1\);
    
    next_r0_0_cry_10 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[10]\, B => \sum0_5[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_9\, S
         => next_r0_0_cry_10_S, Y => OPEN, FCO => 
        \next_r0_0_cry_10\);
    
    \r13[7]\ : SLE
      port map(D => \r14[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[7]_net_1\);
    
    \r14[2]\ : SLE
      port map(D => \r15[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[2]_net_1\);
    
    \next_r0[21]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_301, C => next_r0_0_cry_21_S, 
        D => W_out_2_i_1_13, Y => \Wt_data[21]\);
    
    \r10[14]\ : SLE
      port map(D => \r11[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[14]_net_1\);
    
    next_r0_0_cry_20 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[20]\, B => \sum0_5[20]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_19\, S
         => next_r0_0_cry_20_S, Y => OPEN, FCO => 
        \next_r0_0_cry_20\);
    
    \r15[10]\ : SLE
      port map(D => \r0[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[10]_net_1\);
    
    \r10[12]\ : SLE
      port map(D => \r11[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[12]_net_1\);
    
    \r8[25]\ : SLE
      port map(D => \r9[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[25]_net_1\);
    
    \r6[10]\ : SLE
      port map(D => \r7[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[10]_net_1\);
    
    \r7[14]\ : SLE
      port map(D => \r8[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[14]_net_1\);
    
    sum0_4_axb_0 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[10]_net_1\, B => \s0[0]_net_1\, C => 
        \r15[19]_net_1\, D => \r15[17]_net_1\, Y => \sum0_4[0]\);
    
    \r15[20]\ : SLE
      port map(D => \r0[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[20]_net_1\);
    
    \r2[20]\ : SLE
      port map(D => \r3[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[20]_net_1\);
    
    \next_r0[16]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_286, C => next_r0_0_cry_16_S, 
        D => W_out_2_i_1_8, Y => \Wt_data[16]\);
    
    sum0_4_cry_13 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[13]\, C => 
        \sum0_4_axb_13\, D => GND_net_1, FCI => \sum0_4_cry_12\, 
        S => \sum0_4[13]\, Y => OPEN, FCO => \sum0_4_cry_13\);
    
    sum0_4_axb_4 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[14]_net_1\, B => \s0[4]_net_1\, C => 
        \r15[23]_net_1\, D => \r15[21]_net_1\, Y => 
        \sum0_4_axb_4\);
    
    \r0[22]\ : SLE
      port map(D => \Wt_data[22]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[22]_net_1\);
    
    \r13[24]\ : SLE
      port map(D => \r14[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[24]_net_1\);
    
    \r12[26]\ : SLE
      port map(D => \r13[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[26]_net_1\);
    
    \r10[26]\ : SLE
      port map(D => \r11[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[26]_net_1\);
    
    \r2[31]\ : SLE
      port map(D => \r3[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[31]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \r0[12]\ : SLE
      port map(D => \Wt_data[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[12]_net_1\);
    
    sum0_5_cry_24 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[24]_net_1\, B => \r10[24]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_23\, S => 
        \sum0_5[24]\, Y => OPEN, FCO => \sum0_5_cry_24\);
    
    \r13[22]\ : SLE
      port map(D => \r14[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[22]_net_1\);
    
    \r8[17]\ : SLE
      port map(D => \r9[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[17]_net_1\);
    
    \r11[31]\ : SLE
      port map(D => \r12[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[31]_net_1\);
    
    \r0[0]\ : SLE
      port map(D => \Wt_data[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[0]_net_1\);
    
    \r5[2]\ : SLE
      port map(D => \r6[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[2]_net_1\);
    
    \r13[31]\ : SLE
      port map(D => \r14[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[31]_net_1\);
    
    sum0_4_cry_18 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[18]\, C => 
        \sum0_4_axb_18\, D => GND_net_1, FCI => \sum0_4_cry_17\, 
        S => \sum0_4[18]\, Y => OPEN, FCO => \sum0_4_cry_18\);
    
    \r3[20]\ : SLE
      port map(D => \r4[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[20]_net_1\);
    
    sum0_4_cry_0_1039 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[24]_net_1\, B => \r2[20]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0_0[17]\);
    
    \r12[3]\ : SLE
      port map(D => \r13[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[3]_net_1\);
    
    sum0_4_axb_2 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[12]_net_1\, B => \s0[2]_net_1\, C => 
        \r15[21]_net_1\, D => \r15[19]_net_1\, Y => 
        \sum0_4_axb_2\);
    
    sum0_4_cry_0_1050 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[24]_net_1\, B => \r2[13]_net_1\, C => 
        \r2[9]_net_1\, Y => \s0_0[6]\);
    
    sum0_4_axb_7 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[17]_net_1\, B => \s0[7]_net_1\, C => 
        \r15[26]_net_1\, D => \r15[24]_net_1\, Y => 
        \sum0_4_axb_7\);
    
    \r13[18]\ : SLE
      port map(D => \r14[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[18]_net_1\);
    
    \r12[18]\ : SLE
      port map(D => \r13[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[18]_net_1\);
    
    \r1[14]\ : SLE
      port map(D => \r2[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[14]_net_1\);
    
    \r8[22]\ : SLE
      port map(D => \r9[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[22]_net_1\);
    
    \r5[4]\ : SLE
      port map(D => \r6[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[4]_net_1\);
    
    \r3[2]\ : SLE
      port map(D => \r4[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[2]_net_1\);
    
    sum0_5_cry_1 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[1]_net_1\, B => \r10[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_0\, S => 
        \sum0_5[1]\, Y => OPEN, FCO => \sum0_5_cry_1\);
    
    sum0_5_cry_15 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[15]_net_1\, B => \r10[15]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_14\, S => 
        \sum0_5[15]\, Y => OPEN, FCO => \sum0_5_cry_15\);
    
    \s0[30]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \r2[5]_net_1\, B => \r2[16]_net_1\, Y => 
        \s0[30]_net_1\);
    
    next_r0_0_cry_30 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[30]\, B => \sum0_5[30]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_29\, S
         => next_r0_0_cry_30_S, Y => OPEN, FCO => 
        \next_r0_0_cry_30\);
    
    \r9[1]\ : SLE
      port map(D => \r10[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[1]_net_1\);
    
    \r7[6]\ : SLE
      port map(D => \r8[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[6]_net_1\);
    
    sum0_4_axb_24 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[9]_net_1\, B => \r15[11]_net_1\, C => 
        \s0[24]_net_1\, Y => \sum0_4_axb_24\);
    
    \r11[27]\ : SLE
      port map(D => \r12[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[27]_net_1\);
    
    \r7[29]\ : SLE
      port map(D => \r8[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[29]_net_1\);
    
    \r1[7]\ : SLE
      port map(D => \r2[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[7]_net_1\);
    
    \r11[17]\ : SLE
      port map(D => \r12[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[17]_net_1\);
    
    \r7[8]\ : SLE
      port map(D => \r8[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[8]_net_1\);
    
    \next_r0[4]\ : CFG4
      generic map(INIT => x"CFCA")

      port map(A => N_248, B => next_r0_0_cry_4_S, C => ld_i_i_3, 
        D => W_out_2_0_0_1, Y => \Wt_data[4]\);
    
    \r6[8]\ : SLE
      port map(D => \r7[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[8]_net_1\);
    
    \r13[0]\ : SLE
      port map(D => \r14[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[0]_net_1\);
    
    \r12[4]\ : SLE
      port map(D => \r13[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[4]_net_1\);
    
    \r10[0]\ : SLE
      port map(D => \r11[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[0]_net_1\);
    
    \r9[16]\ : SLE
      port map(D => \r10[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[16]_net_1\);
    
    \r10[16]\ : SLE
      port map(D => \r11[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[16]_net_1\);
    
    sum0_4_cry_0_1047 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[27]_net_1\, B => \r2[16]_net_1\, C => 
        \r2[12]_net_1\, Y => \s0_0[9]\);
    
    \r8[8]\ : SLE
      port map(D => \r9[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[8]_net_1\);
    
    \r8[18]\ : SLE
      port map(D => \r9[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[18]_net_1\);
    
    \r15[15]\ : SLE
      port map(D => \r0[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[15]_net_1\);
    
    \r14[30]\ : SLE
      port map(D => \r15[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[30]_net_1\);
    
    \r14[10]\ : SLE
      port map(D => \r15[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[10]_net_1\);
    
    \r3[30]\ : SLE
      port map(D => \r4[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[30]_net_1\);
    
    sum0_4_axb_27 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[12]_net_1\, B => \s0[27]_net_1\, C => 
        \r15[14]_net_1\, Y => \sum0_4_axb_27\);
    
    \r5[27]\ : SLE
      port map(D => \r6[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[27]_net_1\);
    
    \r3[16]\ : SLE
      port map(D => \r4[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[16]_net_1\);
    
    \r6[29]\ : SLE
      port map(D => \r7[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[29]_net_1\);
    
    \r15[25]\ : SLE
      port map(D => \r0[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[25]_net_1\);
    
    \next_r0[2]\ : CFG4
      generic map(INIT => x"C0E2")

      port map(A => N_98, B => ld_i_i_3, C => next_r0_0_cry_2_S, 
        D => W_out_i_0(2), Y => \Wt_data[2]\);
    
    \r3[8]\ : SLE
      port map(D => \r4[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[8]_net_1\);
    
    \r13[26]\ : SLE
      port map(D => \r14[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[26]_net_1\);
    
    \r9[11]\ : SLE
      port map(D => \r10[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[11]_net_1\);
    
    \next_r0[11]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_268, C => next_r0_0_cry_11_S, 
        D => W_out_2_i_1_3, Y => \Wt_data[11]\);
    
    sum0_4_cry_0_1029 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[13]_net_1\, B => \r2[2]_net_1\, C => 
        \r2[30]_net_1\, Y => \s0_0[27]\);
    
    sum0_4_cry_30 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[30]\, C => 
        \sum0_4_axb_30\, D => GND_net_1, FCI => \sum0_4_cry_29\, 
        S => \sum0_4[30]\, Y => OPEN, FCO => \sum0_4_cry_30\);
    
    \r1[20]\ : SLE
      port map(D => \r2[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[20]_net_1\);
    
    \r13[11]\ : SLE
      port map(D => \r14[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[11]_net_1\);
    
    \r12[11]\ : SLE
      port map(D => \r13[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[11]_net_1\);
    
    \r10[7]\ : SLE
      port map(D => \r11[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[7]_net_1\);
    
    \r5[10]\ : SLE
      port map(D => \r6[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[10]_net_1\);
    
    sum0_4_cry_0_1051 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[23]_net_1\, B => \r2[12]_net_1\, C => 
        \r2[8]_net_1\, Y => \s0_0[5]\);
    
    \r9[9]\ : SLE
      port map(D => \r10[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[9]_net_1\);
    
    \r4[20]\ : SLE
      port map(D => \r5[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[20]_net_1\);
    
    \r3[11]\ : SLE
      port map(D => \r4[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[11]_net_1\);
    
    sum0_4_axb_13 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[0]_net_1\, B => \r15[30]_net_1\, C => 
        \r15[23]_net_1\, D => \s0[13]_net_1\, Y => 
        \sum0_4_axb_13\);
    
    sum0_4_cry_19 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[19]\, C => 
        \sum0_4_axb_19\, D => GND_net_1, FCI => \sum0_4_cry_18\, 
        S => \sum0_4[19]\, Y => OPEN, FCO => \sum0_4_cry_19\);
    
    \r10[4]\ : SLE
      port map(D => \r11[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[4]_net_1\);
    
    sum0_4_cry_0_1037 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[26]_net_1\, B => \r2[22]_net_1\, C => 
        \r2[5]_net_1\, Y => \s0_0[19]\);
    
    sum0_4_axb_10 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[20]_net_1\, B => \s0[10]_net_1\, C => 
        \r15[29]_net_1\, D => \r15[27]_net_1\, Y => 
        \sum0_4_axb_10\);
    
    \r5[9]\ : SLE
      port map(D => \r6[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[9]_net_1\);
    
    \r2[7]\ : SLE
      port map(D => \r3[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[7]_net_1\);
    
    \r2[10]\ : SLE
      port map(D => \r3[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[10]_net_1\);
    
    \r10[30]\ : SLE
      port map(D => \r11[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[30]_net_1\);
    
    sum0_5_cry_5 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[5]_net_1\, B => \r10[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_4\, S => 
        \sum0_5[5]\, Y => OPEN, FCO => \sum0_5_cry_5\);
    
    sum0_4_cry_16 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[16]\, C => 
        \sum0_4_axb_16\, D => GND_net_1, FCI => \sum0_4_cry_15\, 
        S => \sum0_4[16]\, Y => OPEN, FCO => \sum0_4_cry_16\);
    
    \r9[13]\ : SLE
      port map(D => \r10[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[13]_net_1\);
    
    \r3[4]\ : SLE
      port map(D => \r4[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[4]_net_1\);
    
    \r5[28]\ : SLE
      port map(D => \r6[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[28]_net_1\);
    
    \r6[31]\ : SLE
      port map(D => \r7[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[31]_net_1\);
    
    \r6[19]\ : SLE
      port map(D => \r7[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[19]_net_1\);
    
    \r12[30]\ : SLE
      port map(D => \r13[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[30]_net_1\);
    
    \r3[13]\ : SLE
      port map(D => \r4[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[13]_net_1\);
    
    \next_r0[9]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_263, C => next_r0_0_cry_9_S, 
        D => W_out_2_i_1_1, Y => \Wt_data[9]\);
    
    \r2[29]\ : SLE
      port map(D => \r3[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[29]_net_1\);
    
    \r11[23]\ : SLE
      port map(D => \r12[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[23]_net_1\);
    
    \r10[3]\ : SLE
      port map(D => \r11[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[3]_net_1\);
    
    \r4[16]\ : SLE
      port map(D => \r5[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[16]_net_1\);
    
    \r4[8]\ : SLE
      port map(D => \r5[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[8]_net_1\);
    
    \r11[13]\ : SLE
      port map(D => \r12[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[13]_net_1\);
    
    next_r0_0_cry_16 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[16]\, B => \sum0_5[16]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_15\, S
         => next_r0_0_cry_16_S, Y => OPEN, FCO => 
        \next_r0_0_cry_16\);
    
    \r4[30]\ : SLE
      port map(D => \r5[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[30]_net_1\);
    
    \r14[6]\ : SLE
      port map(D => \r15[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[6]_net_1\);
    
    \r14[15]\ : SLE
      port map(D => \r15[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[15]_net_1\);
    
    next_r0_0_cry_26 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[26]\, B => \sum0_5[26]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_25\, S
         => next_r0_0_cry_26_S, Y => OPEN, FCO => 
        \next_r0_0_cry_26\);
    
    \r15[17]\ : SLE
      port map(D => \r0[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[17]_net_1\);
    
    \r9[20]\ : SLE
      port map(D => \r10[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[20]_net_1\);
    
    \r15[27]\ : SLE
      port map(D => \r0[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[27]_net_1\);
    
    \r3[29]\ : SLE
      port map(D => \r4[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[29]_net_1\);
    
    \r7[2]\ : SLE
      port map(D => \r8[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[2]_net_1\);
    
    \r3[0]\ : SLE
      port map(D => \r4[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[0]_net_1\);
    
    \r11[29]\ : SLE
      port map(D => \r12[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[29]_net_1\);
    
    sum0_4_cry_21 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[21]\, C => 
        \sum0_4_axb_21\, D => GND_net_1, FCI => \sum0_4_cry_20\, 
        S => \sum0_4[21]\, Y => OPEN, FCO => \sum0_4_cry_21\);
    
    sum0_4_cry_12 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[12]\, C => 
        \sum0_4_axb_12\, D => GND_net_1, FCI => \sum0_4_cry_11\, 
        S => \sum0_4[12]\, Y => OPEN, FCO => \sum0_4_cry_12\);
    
    \r4[11]\ : SLE
      port map(D => \r5[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[11]_net_1\);
    
    \r1[8]\ : SLE
      port map(D => \r2[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[8]_net_1\);
    
    \r11[19]\ : SLE
      port map(D => \r12[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[19]_net_1\);
    
    \r0[9]\ : SLE
      port map(D => \Wt_data[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[9]_net_1\);
    
    \next_r0[25]\ : CFG4
      generic map(INIT => x"C0C5")

      port map(A => W_out_2_i_1_17, B => next_r0_0_cry_25_S, C
         => ld_i_i_3, D => W_out_2_i_0(25), Y => \Wt_data[25]\);
    
    \r5[1]\ : SLE
      port map(D => \r6[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[1]_net_1\);
    
    next_r0_0_cry_12 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[12]\, B => \sum0_5[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_11\, S
         => next_r0_0_cry_12_S, Y => OPEN, FCO => 
        \next_r0_0_cry_12\);
    
    sum0_4_cry_9 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[9]\, C => 
        \sum0_4_axb_9\, D => GND_net_1, FCI => \sum0_4_cry_8\, S
         => \sum0_4[9]\, Y => OPEN, FCO => \sum0_4_cry_9\);
    
    \r8[15]\ : SLE
      port map(D => \r9[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[15]_net_1\);
    
    next_r0_0_cry_22 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[22]\, B => \sum0_5[22]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_21\, S
         => next_r0_0_cry_22_S, Y => OPEN, FCO => 
        \next_r0_0_cry_22\);
    
    sum0_5_cry_2 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[2]_net_1\, B => \r10[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_1\, S => 
        \sum0_5[2]\, Y => OPEN, FCO => \sum0_5_cry_2\);
    
    sum0_5_cry_25 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[25]_net_1\, B => \r10[25]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_24\, S => 
        \sum0_5[25]\, Y => OPEN, FCO => \sum0_5_cry_25\);
    
    \r7[16]\ : SLE
      port map(D => \r8[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[16]_net_1\);
    
    \r8[7]\ : SLE
      port map(D => \r9[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[7]_net_1\);
    
    sum0_4_cry_0_1027 : CFG2
      generic map(INIT => x"6")

      port map(A => \r2[4]_net_1\, B => \r2[15]_net_1\, Y => 
        \s0_0[29]\);
    
    sum0_5_cry_9 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[9]_net_1\, B => \r10[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_8\, S => 
        \sum0_5[9]\, Y => OPEN, FCO => \sum0_5_cry_9\);
    
    sum0_5_cry_8 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[8]_net_1\, B => \r10[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_7\, S => 
        \sum0_5[8]\, Y => OPEN, FCO => \sum0_5_cry_8\);
    
    \r7[24]\ : SLE
      port map(D => \r8[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[24]_net_1\);
    
    \r1[3]\ : SLE
      port map(D => \r2[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[3]_net_1\);
    
    \s0[2]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[20]_net_1\, B => \r2[9]_net_1\, C => 
        \r2[5]_net_1\, Y => \s0[2]_net_1\);
    
    \s0[24]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[27]_net_1\, C => 
        \r2[10]_net_1\, Y => \s0[24]_net_1\);
    
    next_r0_0_cry_17 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[17]\, B => \sum0_5[17]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_16\, S
         => next_r0_0_cry_17_S, Y => OPEN, FCO => 
        \next_r0_0_cry_17\);
    
    \s0[14]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[0]_net_1\, B => \r2[17]_net_1\, C => 
        \r2[21]_net_1\, Y => \s0[14]_net_1\);
    
    \r7[1]\ : SLE
      port map(D => \r8[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[1]_net_1\);
    
    next_r0_0_cry_27 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[27]\, B => \sum0_5[27]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_26\, S
         => next_r0_0_cry_27_S, Y => OPEN, FCO => 
        \next_r0_0_cry_27\);
    
    \next_r0[24]\ : CFG4
      generic map(INIT => x"C0C5")

      port map(A => W_out_2_i_1_16, B => next_r0_0_cry_24_S, C
         => ld_i_i_3, D => W_out_2_i_0(24), Y => \Wt_data[24]\);
    
    \r1[31]\ : SLE
      port map(D => \r2[31]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[31]_net_1\);
    
    \r11[24]\ : SLE
      port map(D => \r12[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[24]_net_1\);
    
    \next_r0[27]\ : CFG4
      generic map(INIT => x"C0C5")

      port map(A => W_out_2_i_1_19, B => next_r0_0_cry_27_S, C
         => ld_i_i_3, D => W_out_2_i_0(27), Y => \Wt_data[27]\);
    
    next_r0_0_cry_15 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[15]\, B => \sum0_5[15]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_14\, S
         => next_r0_0_cry_15_S, Y => OPEN, FCO => 
        \next_r0_0_cry_15\);
    
    \r13[8]\ : SLE
      port map(D => \r14[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r13[8]_net_1\);
    
    \r11[22]\ : SLE
      port map(D => \r12[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[22]_net_1\);
    
    \r11[14]\ : SLE
      port map(D => \r12[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[14]_net_1\);
    
    \r4[13]\ : SLE
      port map(D => \r5[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[13]_net_1\);
    
    next_r0_0_cry_25 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[25]\, B => \sum0_5[25]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_24\, S
         => next_r0_0_cry_25_S, Y => OPEN, FCO => 
        \next_r0_0_cry_25\);
    
    \r7[11]\ : SLE
      port map(D => \r8[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[11]_net_1\);
    
    \r11[12]\ : SLE
      port map(D => \r12[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[12]_net_1\);
    
    \r5[3]\ : SLE
      port map(D => \r6[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[3]_net_1\);
    
    \r6[24]\ : SLE
      port map(D => \r7[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[24]_net_1\);
    
    \s0[22]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[29]_net_1\, B => \r2[25]_net_1\, C => 
        \r2[8]_net_1\, Y => \s0[22]_net_1\);
    
    \next_r0[0]\ : CFG4
      generic map(INIT => x"A3A0")

      port map(A => \next_r0_0_cry_0_Y\, B => W_out_i_0(0), C => 
        ld_i_i_3, D => N_98, Y => \Wt_data[0]\);
    
    \r0[20]\ : SLE
      port map(D => \Wt_data[20]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[20]_net_1\);
    
    \r4[4]\ : SLE
      port map(D => \r5[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[4]_net_1\);
    
    \s0[12]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[30]_net_1\, B => \r2[19]_net_1\, C => 
        \r2[15]_net_1\, Y => \s0[12]_net_1\);
    
    \r15[1]\ : SLE
      port map(D => \r0[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[1]_net_1\);
    
    \r8[1]\ : SLE
      port map(D => \r9[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[1]_net_1\);
    
    \r12[28]\ : SLE
      port map(D => \r13[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[28]_net_1\);
    
    \r10[28]\ : SLE
      port map(D => \r11[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[28]_net_1\);
    
    \r0[10]\ : SLE
      port map(D => \Wt_data[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[10]_net_1\);
    
    \r1[16]\ : SLE
      port map(D => \r2[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[16]_net_1\);
    
    \next_r0[28]\ : CFG4
      generic map(INIT => x"C0C5")

      port map(A => W_out_2_i_1_20, B => next_r0_0_cry_28_S, C
         => ld_i_i_3, D => W_out_2_i_0(28), Y => \Wt_data[28]\);
    
    \r8[12]\ : SLE
      port map(D => \r9[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[12]_net_1\);
    
    \r12[1]\ : SLE
      port map(D => \r13[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r12[1]_net_1\);
    
    \r5[25]\ : SLE
      port map(D => \r6[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[25]_net_1\);
    
    sum0_4_axb_1 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[11]_net_1\, B => \s0[1]_net_1\, C => 
        \r15[20]_net_1\, D => \r15[18]_net_1\, Y => 
        \sum0_4_axb_1\);
    
    \r14[17]\ : SLE
      port map(D => \r15[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[17]_net_1\);
    
    \r1[29]\ : SLE
      port map(D => \r2[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[29]_net_1\);
    
    \r9[17]\ : SLE
      port map(D => \r10[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r9[17]_net_1\);
    
    sum0_4_cry_0_1040 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[19]_net_1\, B => \r2[2]_net_1\, C => 
        \r2[23]_net_1\, Y => \s0_0[16]\);
    
    \r5[19]\ : SLE
      port map(D => \r6[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r5[19]_net_1\);
    
    \r11[7]\ : SLE
      port map(D => \r12[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[7]_net_1\);
    
    \r4[29]\ : SLE
      port map(D => \r5[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[29]_net_1\);
    
    \r4[6]\ : SLE
      port map(D => \r5[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[6]_net_1\);
    
    \r15[13]\ : SLE
      port map(D => \r0[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[13]_net_1\);
    
    \r11[4]\ : SLE
      port map(D => \r12[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[4]_net_1\);
    
    \r7[13]\ : SLE
      port map(D => \r8[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[13]_net_1\);
    
    \r3[17]\ : SLE
      port map(D => \r4[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r3[17]_net_1\);
    
    \r1[11]\ : SLE
      port map(D => \r2[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r1[11]_net_1\);
    
    \r15[23]\ : SLE
      port map(D => \r0[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[23]_net_1\);
    
    sum0_4_axb_14 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[1]_net_1\, B => \r15[31]_net_1\, C => 
        \r15[24]_net_1\, D => \s0[14]_net_1\, Y => 
        \sum0_4_axb_14\);
    
    \r4[1]\ : SLE
      port map(D => \r5[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r4[1]_net_1\);
    
    \r8[20]\ : SLE
      port map(D => \r9[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r8[20]_net_1\);
    
    \r15[7]\ : SLE
      port map(D => \r0[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[7]_net_1\);
    
    \r2[9]\ : SLE
      port map(D => \r3[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[9]_net_1\);
    
    next_r0_0_s_31 : ARI1
      generic map(INIT => x"46600")

      port map(A => VCC_net_1, B => \sum0_4[31]\, C => 
        \sum0_5[31]\, D => GND_net_1, FCI => \next_r0_0_cry_30\, 
        S => next_r0_0_s_31_S, Y => OPEN, FCO => OPEN);
    
    \r2[19]\ : SLE
      port map(D => \r3[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[19]_net_1\);
    
    \r14[20]\ : SLE
      port map(D => \r15[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[20]_net_1\);
    
    \r15[19]\ : SLE
      port map(D => \r0[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[19]_net_1\);
    
    \r14[7]\ : SLE
      port map(D => \r15[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r14[7]_net_1\);
    
    \r6[14]\ : SLE
      port map(D => \r7[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[14]_net_1\);
    
    \r6[1]\ : SLE
      port map(D => \r7[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r6[1]_net_1\);
    
    \r10[18]\ : SLE
      port map(D => \r11[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r10[18]_net_1\);
    
    \r15[29]\ : SLE
      port map(D => \r0[29]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r15[29]_net_1\);
    
    sum0_4_axb_17 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[2]_net_1\, B => \r15[4]_net_1\, C => 
        \s0[17]_net_1\, D => \r15[27]_net_1\, Y => 
        \sum0_4_axb_17\);
    
    \next_r0[15]\ : CFG4
      generic map(INIT => x"FE54")

      port map(A => ld_i_i_3, B => W_out_2_0_0_12, C => 
        W_out_2_0_a4_1_0_RNIFI1DA(23), D => next_r0_0_cry_15_S, Y
         => \Wt_data[15]\);
    
    \r2[24]\ : SLE
      port map(D => \r3[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r2[24]_net_1\);
    
    \r11[26]\ : SLE
      port map(D => \r12[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[26]_net_1\);
    
    \r0[31]\ : SLE
      port map(D => \Wt_data[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r0[31]_net_1\);
    
    \r7[30]\ : SLE
      port map(D => \r8[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r7[30]_net_1\);
    
    \next_r0[7]\ : CFG4
      generic map(INIT => x"AFAC")

      port map(A => next_r0_0_cry_7_S, B => W_out_2_0_1(7), C => 
        ld_i_i_3, D => W_out_2_0_0_4, Y => \Wt_data[7]\);
    
    \r11[16]\ : SLE
      port map(D => \r12[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_244_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \r11[16]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_kt_rom is

    port( hash_control_st_reg_ns_i_0_a2_0 : in    std_logic_vector(4 to 4);
          hash_control_st_reg_ns_i_0_a2_2 : out   std_logic_vector(4 to 4);
          Kt_addr                         : in    std_logic_vector(5 downto 0);
          Kt_addr_fast                    : in    std_logic_vector(4 downto 0);
          Kt_data_0                       : out   std_logic;
          Kt_data_24                      : out   std_logic;
          Kt_data_15                      : out   std_logic;
          m10_bm                          : out   std_logic;
          m20_1                           : out   std_logic;
          m10_am                          : out   std_logic;
          Kt_addr_5_rep1                  : in    std_logic;
          Kt_addr_3_rep2                  : in    std_logic;
          Kt_addr_3_rep1                  : in    std_logic;
          m62_am                          : out   std_logic;
          Kt_addr_0_rep1                  : in    std_logic;
          m104_bm                         : out   std_logic;
          Kt_addr_2_rep1                  : in    std_logic;
          Kt_addr_0_rep2                  : in    std_logic;
          m49_am                          : out   std_logic;
          Kt_addr_1_rep1                  : in    std_logic;
          m49_bm                          : out   std_logic;
          m137_am                         : out   std_logic;
          m137_bm                         : out   std_logic;
          Kt_addr_2_rep2                  : in    std_logic;
          Kt_addr_1_rep2                  : in    std_logic;
          Kt_addr_4_rep2                  : in    std_logic;
          m215_am                         : out   std_logic;
          Kt_addr_4_rep1                  : in    std_logic;
          m215_bm                         : out   std_logic;
          m250_am                         : out   std_logic;
          m250_bm                         : out   std_logic;
          m207_1_1                        : out   std_logic;
          m207_1_0                        : out   std_logic;
          m95_1_1                         : out   std_logic;
          m95_1_0                         : out   std_logic;
          m197_1_1                        : out   std_logic;
          m197_1_0                        : out   std_logic;
          m316                            : out   std_logic;
          m34                             : out   std_logic;
          m157                            : out   std_logic;
          m325                            : out   std_logic;
          m168_1_1                        : out   std_logic;
          m168_1_0                        : out   std_logic;
          m230                            : out   std_logic;
          m296                            : out   std_logic;
          m254                            : out   std_logic;
          m114                            : out   std_logic;
          m304                            : out   std_logic;
          m73_0                           : out   std_logic;
          pad_one_reg_0_0_a2_0            : in    std_logic;
          m239                            : out   std_logic;
          m219                            : out   std_logic;
          m285                            : out   std_logic;
          m177                            : out   std_logic;
          m124                            : out   std_logic;
          m289                            : out   std_logic;
          m78                             : out   std_logic;
          m141                            : out   std_logic;
          i3_mux_1                        : out   std_logic;
          m67_ns                          : out   std_logic;
          m83_ns                          : out   std_logic;
          m110_ns                         : out   std_logic;
          m119_ns                         : out   std_logic;
          m144_ns                         : out   std_logic;
          m172_ns                         : out   std_logic;
          m222_ns                         : out   std_logic;
          m226_ns                         : out   std_logic;
          m235_ns                         : out   std_logic;
          m258_ns                         : out   std_logic;
          m276_ns                         : out   std_logic;
          m281_ns                         : out   std_logic;
          m292_ns                         : out   std_logic;
          m300_ns                         : out   std_logic;
          m273                            : out   std_logic;
          m104_am                         : out   std_logic;
          m62_bm                          : out   std_logic
        );

end sha256_kt_rom;

architecture DEF_ARCH of sha256_kt_rom is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \m10_bm\, \m20_1\, \m10_am\, m19_1_1, m19_1_0, 
        m62_am_1_0, m62_am_1, m54, m53, m51, m304_2, m104_bm_1, 
        m103_1, m79, m78_1, m49_am_1_0, m35, m48_2, m49_bm_1, 
        m48_1, m43, m137_am_1_0, m129, m126, m127, m137_bm_1_0, 
        m137_bm_1, m17, m133, m132, m215_am_1_0, m211_0, m209, 
        m92, m215_bm_1_0, m215_bm_1, m90, m22, m164, m273_2, 
        m250_am_1, m194, m85, m250_bm_1_0_1, m250_bm_1_0, m205, 
        m202, m207_1_0_1, m270_2, m270_1_1, m266, m263, m261, m93, 
        m91, m46, m87, m195, m193, m185, m191, m316_2, m316_1_1, 
        m313, m311, m310, m32, m34_1_2, m30, i2_mux, m23, m155, 
        m157_1_2, m153, m151, m148, 
        \hash_control_st_reg_ns_i_0_a2_2[4]\, m325_1_1, m325_1_0, 
        m323, m318, m325_1_0_1, m186, m188_1_2, m184, m181, m180, 
        m166, m163, m168_1_0_1, m230_0, m230_1_1, m227, m296_2, 
        m296_1_1, m16, m237, m254_1_1, m254_1_0, m252, m232, m105, 
        m1, m114_1_0, m63, m304_1_0, m304_1, m216, m73_1, m73_1_0, 
        m73, m71, m13, m239_1_2, m81, m219_1_2, m68, m285_1_1_1, 
        m285_1_1, m28, m177_2, m177_1_0, m177_1, m174, m124_1_2, 
        m120, m122, m289_1_1, m289_1_0, m37, m78_2, m78_1_0, 
        m141_1, m138, m117, m308_ns_1, m67_bm, m67_am, m83_bm, 
        m83_am, m110_bm, m110_am, m119_bm, m119_am, m144_bm, 
        m144_am, m172_bm, m172_am, m222_bm, m222_am, m226_bm, 
        m226_am, m235_bm, m235_am, m258_bm, m258_am, m276_bm, 
        m276_am, m281_bm, m281_am, m292_bm, m292_am, m300_bm, 
        m300_am, m2, m42, m15, m267, m242, m146, m111, m76, m70, 
        m45, m29, m273_0, m273_1, m98, m60, GND_net_1, VCC_net_1
         : std_logic;

begin 

    hash_control_st_reg_ns_i_0_a2_2(4) <= 
        \hash_control_st_reg_ns_i_0_a2_2[4]\;
    m10_bm <= \m10_bm\;
    m20_1 <= \m20_1\;
    m10_am <= \m10_am\;

    \next_rout_31_0_.m313\ : CFG4
      generic map(INIT => x"5A2F")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m313);
    
    \next_rout_31_0_.m71\ : CFG3
      generic map(INIT => x"71")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m71);
    
    \next_rout_31_0_.m227\ : CFG3
      generic map(INIT => x"4E")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep1, Y => m227);
    
    \next_rout_31_0_.m13\ : CFG3
      generic map(INIT => x"1B")

      port map(A => Kt_addr_fast(0), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, Y => m13);
    
    \next_rout_31_0_.m285_1_1\ : CFG4
      generic map(INIT => x"A2BD")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(2), C => 
        Kt_addr(1), D => m285_1_1_1, Y => m285_1_1);
    
    \next_rout_31_0_.m216\ : CFG3
      generic map(INIT => x"4A")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep1, Y => m216);
    
    \next_rout_31_0_.m2\ : CFG3
      generic map(INIT => x"21")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_0_rep1, C => 
        Kt_addr_1_rep1, Y => m2);
    
    \next_rout_31_0_.m137_am\ : CFG4
      generic map(INIT => x"EBAB")

      port map(A => m304_2, B => m137_am_1_0, C => Kt_addr_3_rep2, 
        D => m129, Y => m137_am);
    
    \next_rout_31_0_.m10_am\ : CFG4
      generic map(INIT => x"BA89")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => \m10_am\);
    
    \next_rout_31_0_.m289\ : CFG3
      generic map(INIT => x"47")

      port map(A => m289_1_1, B => Kt_addr(3), C => m289_1_0, Y
         => m289);
    
    \next_rout_31_0_.m177_1_0\ : CFG4
      generic map(INIT => x"0A1B")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => m174, D
         => pad_one_reg_0_0_a2_0, Y => m177_1_0);
    
    \next_rout_31_0_.m98\ : CFG4
      generic map(INIT => x"3479")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m98);
    
    \next_rout_31_0_.m119_am\ : CFG4
      generic map(INIT => x"D585")

      port map(A => Kt_addr_4_rep2, B => pad_one_reg_0_0_a2_0, C
         => Kt_addr_0_rep2, D => Kt_addr(1), Y => m119_am);
    
    \next_rout_31_0_.m250_am\ : CFG4
      generic map(INIT => x"0051")

      port map(A => m273_2, B => m250_am_1, C => Kt_addr_3_rep2, 
        D => m48_1, Y => m250_am);
    
    \next_rout_31_0_.m157_1_2\ : CFG4
      generic map(INIT => x"2637")

      port map(A => Kt_addr_5_rep1, B => Kt_addr_3_rep2, C => 
        m151, D => m148, Y => m157_1_2);
    
    \next_rout_31_0_.m141\ : CFG3
      generic map(INIT => x"FD")

      port map(A => m141_1, B => m211_0, C => m177_1, Y => m141);
    
    \next_rout_31_0_.m235_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m235_bm, C => m235_am, Y => 
        m235_ns);
    
    \next_rout_31_0_.m104_bm_1\ : CFG4
      generic map(INIT => x"41EB")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_0_rep1, D => m79, Y => m104_bm_1);
    
    \next_rout_31_0_.m144_am\ : CFG4
      generic map(INIT => x"011C")

      port map(A => Kt_addr(1), B => Kt_addr_4_rep2, C => 
        Kt_addr(2), D => Kt_addr_0_rep2, Y => m144_am);
    
    \next_rout_31_0_.m270_1_1\ : CFG4
      generic map(INIT => x"2637")

      port map(A => Kt_addr_5_rep1, B => Kt_addr_3_rep2, C => 
        m263, D => m261, Y => m270_1_1);
    
    \next_rout_31_0_.m289_1_0\ : CFG3
      generic map(INIT => x"74")

      port map(A => m237, B => Kt_addr(4), C => m46, Y => 
        m289_1_0);
    
    \next_rout_31_0_.m51\ : CFG3
      generic map(INIT => x"15")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m51);
    
    \next_rout_31_0_.m67_am\ : CFG4
      generic map(INIT => x"80D5")

      port map(A => Kt_addr_4_rep1, B => Kt_addr(2), C => 
        Kt_addr(1), D => m63, Y => m67_am);
    
    \next_rout_31_0_.m207_1_1\ : CFG3
      generic map(INIT => x"74")

      port map(A => m205, B => Kt_addr_3_rep2, C => m202, Y => 
        m207_1_1);
    
    \next_rout_31_0_.m168_1_0\ : CFG4
      generic map(INIT => x"2C5A")

      port map(A => Kt_addr_4_rep2, B => Kt_addr_3_rep2, C => 
        m168_1_0_1, D => Kt_addr(0), Y => m168_1_0);
    
    \next_rout_31_0_.m92\ : CFG3
      generic map(INIT => x"79")

      port map(A => Kt_addr_fast(1), B => Kt_addr_fast(0), C => 
        Kt_addr_2_rep1, Y => m92);
    
    \next_rout_31_0_.m62_am_1\ : CFG4
      generic map(INIT => x"0A1B")

      port map(A => Kt_addr_fast(4), B => Kt_addr_0_rep1, C => 
        m51, D => hash_control_st_reg_ns_i_0_a2_0(4), Y => 
        m62_am_1);
    
    \next_rout_31_0_.m43\ : CFG3
      generic map(INIT => x"4D")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m43);
    
    \next_rout_31_0_.m62_am\ : CFG3
      generic map(INIT => x"72")

      port map(A => Kt_addr_3_rep1, B => m62_am_1_0, C => 
        m62_am_1, Y => m62_am);
    
    \next_rout_31_0_.m316_3\ : CFG4
      generic map(INIT => x"8008")

      port map(A => Kt_addr_5_rep1, B => Kt_addr(3), C => 
        Kt_addr(4), D => m126, Y => m316_2);
    
    \next_rout_31_0_.m40_2\ : CFG3
      generic map(INIT => x"40")

      port map(A => Kt_addr_fast(4), B => m37, C => 
        Kt_addr_fast(3), Y => m78_1);
    
    \next_rout_31_0_.m292_am\ : CFG4
      generic map(INIT => x"E4EE")

      port map(A => Kt_addr(4), B => m54, C => Kt_addr(2), D => 
        Kt_addr(1), Y => m292_am);
    
    \next_rout_31_0_.m114_1_0\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr_3_rep2, B => m63, C => m35, Y => 
        m114_1_0);
    
    \next_rout_31_0_.m34\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => m32, B => Kt_addr_5_rep1, C => m34_1_2, D => 
        m30, Y => m34);
    
    \next_rout_31_0_.m23\ : CFG4
      generic map(INIT => x"75C3")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m23);
    
    \next_rout_31_0_.m166\ : CFG4
      generic map(INIT => x"5214")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_4_rep1, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m166);
    
    \next_rout_31_0_.m202\ : CFG4
      generic map(INIT => x"38BA")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m202);
    
    \next_rout_31_0_.m67_bm\ : CFG4
      generic map(INIT => x"494F")

      port map(A => Kt_addr_4_rep1, B => Kt_addr(2), C => 
        Kt_addr_0_rep2, D => Kt_addr(1), Y => m67_bm);
    
    \next_rout_31_0_.m226_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m226_bm, B => Kt_addr(3), C => m226_am, Y => 
        m226_ns);
    
    \next_rout_31_0_.m137_bm_1_0\ : CFG4
      generic map(INIT => x"5D08")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => m17, Y => m137_bm_1_0);
    
    \next_rout_31_0_.m83_am\ : CFG4
      generic map(INIT => x"52A7")

      port map(A => Kt_addr_4_rep2, B => m42, C => Kt_addr_0_rep2, 
        D => Kt_addr(1), Y => m83_am);
    
    \next_rout_31_0_.m70\ : CFG3
      generic map(INIT => x"79")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m70);
    
    \next_rout_31_0_.m104_am\ : CFG4
      generic map(INIT => x"1D0C")

      port map(A => Kt_addr_0_rep2, B => Kt_addr_3_rep1, C => m98, 
        D => m42, Y => m104_am);
    
    \next_rout_31_0_.m308_ns\ : CFG4
      generic map(INIT => x"B964")

      port map(A => Kt_addr(3), B => Kt_addr(4), C => m117, D => 
        m308_ns_1, Y => i3_mux_1);
    
    \next_rout_31_0_.m83_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m83_bm, C => m83_am, Y => 
        m83_ns);
    
    \next_rout_31_0_.m281_am\ : CFG4
      generic map(INIT => x"A2B3")

      port map(A => Kt_addr(0), B => Kt_addr(4), C => m42, D => 
        m15, Y => m281_am);
    
    \next_rout_31_0_.m230\ : CFG4
      generic map(INIT => x"F0F7")

      port map(A => Kt_addr(4), B => Kt_addr(2), C => m230_0, D
         => m230_1_1, Y => m230);
    
    \next_rout_31_0_.m137_bm_1\ : CFG3
      generic map(INIT => x"47")

      port map(A => m133, B => Kt_addr_fast(4), C => m132, Y => 
        m137_bm_1);
    
    \next_rout_31_0_.m310\ : CFG4
      generic map(INIT => x"607C")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m310);
    
    \next_rout_31_0_.m188_1_2\ : CFG4
      generic map(INIT => x"3726")

      port map(A => Kt_addr_5_rep1, B => Kt_addr_3_rep2, C => 
        m181, D => m180, Y => m188_1_2);
    
    \next_rout_31_0_.m133\ : CFG3
      generic map(INIT => x"29")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m133);
    
    \next_rout_31_0_.m110_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m110_bm, B => Kt_addr(3), C => m110_am, Y => 
        m110_ns);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \next_rout_31_0_.m325_1_0\ : CFG4
      generic map(INIT => x"8F85")

      port map(A => Kt_addr_3_rep1, B => m318, C => m325_1_0_1, D
         => hash_control_st_reg_ns_i_0_a2_0(4), Y => m325_1_0);
    
    \next_rout_31_0_.m250_bm_1_0\ : CFG3
      generic map(INIT => x"CB")

      port map(A => Kt_addr_3_rep1, B => Kt_addr_1_rep2, C => 
        m250_bm_1_0_1, Y => m250_bm_1_0);
    
    \next_rout_31_0_.m49_am\ : CFG4
      generic map(INIT => x"0A0D")

      port map(A => Kt_addr_3_rep1, B => Kt_addr_0_rep2, C => 
        m78_1, D => m49_am_1_0, Y => m49_am);
    
    \next_rout_31_0_.m292_bm\ : CFG4
      generic map(INIT => x"280C")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m292_bm);
    
    \next_rout_31_0_.m186\ : CFG4
      generic map(INIT => x"6133")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m186);
    
    \next_rout_31_0_.m60\ : CFG4
      generic map(INIT => x"2B0E")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m60);
    
    \next_rout_31_0_.m49_bm\ : CFG4
      generic map(INIT => x"FFAB")

      port map(A => m48_2, B => m49_bm_1, C => Kt_addr_3_rep1, D
         => m48_1, Y => m49_bm);
    
    \next_rout_31_0_.m177_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_4_rep2, B => m22, C => Kt_addr_3_rep2, 
        Y => m177_2);
    
    \next_rout_31_0_.m15\ : CFG2
      generic map(INIT => x"2")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, Y => m15);
    
    \next_rout_31_0_.m132\ : CFG3
      generic map(INIT => x"3B")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m132);
    
    \next_rout_31_0_.m273_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => Kt_addr_4_rep1, B => m68, C => Kt_addr_3_rep1, 
        Y => m73);
    
    \next_rout_31_0_.m48_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_fast(4), B => m46, C => 
        Kt_addr_fast(3), Y => m48_2);
    
    \next_rout_31_0_.m114_1\ : CFG3
      generic map(INIT => x"02")

      port map(A => Kt_addr_4_rep1, B => m111, C => 
        Kt_addr_3_rep1, Y => m230_0);
    
    \next_rout_31_0_.m258_bm\ : CFG4
      generic map(INIT => x"72FA")

      port map(A => Kt_addr(4), B => Kt_addr(2), C => m120, D => 
        Kt_addr(0), Y => m258_bm);
    
    \next_rout_31_0_.m237\ : CFG3
      generic map(INIT => x"3E")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m237);
    
    \next_rout_31_0_.m157\ : CFG4
      generic map(INIT => x"38F8")

      port map(A => m155, B => Kt_addr_5_rep1, C => m157_1_2, D
         => m153, Y => m157);
    
    \next_rout_31_0_.m126\ : CFG3
      generic map(INIT => x"6E")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m126);
    
    \next_rout_31_0_.m318\ : CFG3
      generic map(INIT => x"36")

      port map(A => Kt_addr_fast(0), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, Y => m318);
    
    \next_rout_31_0_.m151\ : CFG4
      generic map(INIT => x"7B06")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_fast(4), C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m151);
    
    \next_rout_31_0_.m117\ : CFG3
      generic map(INIT => x"19")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m117);
    
    \next_rout_31_0_.m111\ : CFG3
      generic map(INIT => x"7A")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m111);
    
    \next_rout_31_0_.m219_1_2\ : CFG4
      generic map(INIT => x"2367")

      port map(A => Kt_addr_3_rep2, B => Kt_addr_4_rep2, C => m68, 
        D => m216, Y => m219_1_2);
    
    \next_rout_31_0_.m155\ : CFG4
      generic map(INIT => x"69DF")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m155);
    
    \next_rout_31_0_.m45\ : CFG3
      generic map(INIT => x"28")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m45);
    
    \next_rout_31_0_.m137_bm\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m137_bm_1_0, B => Kt_addr_3_rep2, C => 
        m137_bm_1, Y => m137_bm);
    
    \next_rout_31_0_.m304_2\ : CFG4
      generic map(INIT => x"0002")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(4), C => 
        Kt_addr(0), D => m1, Y => m304_1);
    
    \next_rout_31_0_.m35\ : CFG3
      generic map(INIT => x"5E")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m35);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \next_rout_31_0_.m103_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_fast(4), B => m29, C => 
        Kt_addr_fast(3), Y => m304_2);
    
    \next_rout_31_0_.m239\ : CFG4
      generic map(INIT => x"3E32")

      port map(A => m237, B => m239_1_2, C => Kt_addr(4), D => 
        m81, Y => m239);
    
    \next_rout_31_0_.m172_bm\ : CFG4
      generic map(INIT => x"6C1E")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m172_bm);
    
    \next_rout_31_0_.m93\ : CFG4
      generic map(INIT => x"3465")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m93);
    
    \next_rout_31_0_.m76\ : CFG3
      generic map(INIT => x"6D")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m76);
    
    \next_rout_31_0_.m197_1_0\ : CFG4
      generic map(INIT => x"41EB")

      port map(A => Kt_addr_3_rep2, B => Kt_addr_4_rep2, C => 
        m185, D => m191, Y => m197_1_0);
    
    \next_rout_31_0_.m17\ : CFG3
      generic map(INIT => x"38")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m17);
    
    \next_rout_31_0_.m10_bm\ : CFG4
      generic map(INIT => x"4427")

      port map(A => Kt_addr(4), B => Kt_addr(2), C => 
        hash_control_st_reg_ns_i_0_a2_0(4), D => Kt_addr(0), Y
         => \m10_bm\);
    
    \next_rout_31_0_.m215_bm_1_0\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr_4_rep1, B => m90, C => m22, Y => 
        m215_bm_1_0);
    
    \next_rout_31_0_.m266\ : CFG4
      generic map(INIT => x"3733")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m266);
    
    \next_rout_31_0_.m119_bm\ : CFG3
      generic map(INIT => x"E4")

      port map(A => Kt_addr_4_rep2, B => m117, C => m35, Y => 
        m119_bm);
    
    \next_rout_31_0_.m235_bm\ : CFG4
      generic map(INIT => x"7E45")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m235_bm);
    
    \next_rout_31_0_.m292_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m292_bm, C => m292_am, Y => 
        m292_ns);
    
    \next_rout_31_0_.m244_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_4_rep1, B => m242, C => 
        Kt_addr_3_rep1, Y => m273_2);
    
    \next_rout_31_0_.m215_bm\ : CFG3
      generic map(INIT => x"74")

      port map(A => m215_bm_1_0, B => Kt_addr_3_rep2, C => 
        m215_bm_1, Y => m215_bm);
    
    \next_rout_31_0_.m276_am\ : CFG4
      generic map(INIT => x"8827")

      port map(A => Kt_addr(4), B => Kt_addr(1), C => 
        pad_one_reg_0_0_a2_0, D => Kt_addr(0), Y => m276_am);
    
    \next_rout_31_0_.m188\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => m186, B => Kt_addr(5), C => m188_1_2, D => 
        m184, Y => Kt_data_15);
    
    \next_rout_31_0_.m177\ : CFG4
      generic map(INIT => x"FFAB")

      port map(A => m177_2, B => Kt_addr(3), C => m177_1_0, D => 
        m177_1, Y => m177);
    
    \next_rout_31_0_.m141_1_0\ : CFG4
      generic map(INIT => x"6E7F")

      port map(A => Kt_addr_4_rep2, B => Kt_addr_3_rep2, C => m79, 
        D => m138, Y => m141_1);
    
    \next_rout_31_0_.m197_1_1\ : CFG3
      generic map(INIT => x"74")

      port map(A => m195, B => Kt_addr_3_rep2, C => m193, Y => 
        m197_1_1);
    
    \next_rout_31_0_.m300_bm\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(4), B => m146, C => Kt_addr(2), Y => 
        m300_bm);
    
    \next_rout_31_0_.m261\ : CFG4
      generic map(INIT => x"573C")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m261);
    
    \next_rout_31_0_.m258_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m258_bm, C => m258_am, Y => 
        m258_ns);
    
    \next_rout_31_0_.m168_1_1\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr_3_rep2, B => m166, C => m163, Y => 
        m168_1_1);
    
    \next_rout_31_0_.m153\ : CFG4
      generic map(INIT => x"0A10")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m153);
    
    \next_rout_31_0_.m79\ : CFG3
      generic map(INIT => x"3D")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m79);
    
    \next_rout_31_0_.m273\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => m273_1, B => m273_0, C => m273_2, D => m73, Y
         => m273);
    
    \next_rout_31_0_.m141_1\ : CFG4
      generic map(INIT => x"0200")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_3_rep1, C => 
        hash_control_st_reg_ns_i_0_a2_0(4), D => Kt_addr_0_rep1, 
        Y => m211_0);
    
    \next_rout_31_0_.m34_1_2\ : CFG4
      generic map(INIT => x"2637")

      port map(A => Kt_addr_5_rep1, B => Kt_addr_3_rep1, C => 
        i2_mux, D => m23, Y => m34_1_2);
    
    \next_rout_31_0_.m119_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m119_bm, B => Kt_addr(3), C => m119_am, Y => 
        m119_ns);
    
    \next_rout_31_0_.m110_am\ : CFG4
      generic map(INIT => x"E170")

      port map(A => Kt_addr(1), B => Kt_addr_4_rep2, C => 
        Kt_addr(2), D => Kt_addr_0_rep2, Y => m110_am);
    
    \next_rout_31_0_.m296\ : CFG4
      generic map(INIT => x"AEEE")

      port map(A => m296_2, B => m296_1_1, C => Kt_addr(3), D => 
        m16, Y => m296);
    
    \next_rout_31_0_.m321\ : CFG2
      generic map(INIT => x"2")

      port map(A => hash_control_st_reg_ns_i_0_a2_0(4), B => 
        Kt_addr(4), Y => \hash_control_st_reg_ns_i_0_a2_2[4]\);
    
    \next_rout_31_0_.m114\ : CFG4
      generic map(INIT => x"FAFB")

      port map(A => m230_0, B => Kt_addr(4), C => m296_2, D => 
        m114_1_0, Y => m114);
    
    \next_rout_31_0_.m103_2\ : CFG3
      generic map(INIT => x"10")

      port map(A => Kt_addr_fast(4), B => m22, C => 
        Kt_addr_fast(3), Y => m103_1);
    
    \next_rout_31_0_.m67_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m67_bm, C => m67_am, Y => 
        m67_ns);
    
    \next_rout_31_0_.m95_1_0\ : CFG4
      generic map(INIT => x"7520")

      port map(A => Kt_addr_3_rep1, B => Kt_addr_4_rep2, C => m46, 
        D => m87, Y => m95_1_0);
    
    \next_rout_31_0_.m78\ : CFG4
      generic map(INIT => x"FFCD")

      port map(A => Kt_addr(3), B => m78_2, C => m78_1_0, D => 
        m78_1, Y => m78);
    
    \next_rout_31_0_.m37\ : CFG3
      generic map(INIT => x"51")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m37);
    
    \next_rout_31_0_.m207_1_0\ : CFG4
      generic map(INIT => x"67C2")

      port map(A => Kt_addr_4_rep2, B => m207_1_0_1, C => 
        Kt_addr(2), D => Kt_addr(1), Y => m207_1_0);
    
    \next_rout_31_0_.m105\ : CFG3
      generic map(INIT => x"65")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m105);
    
    \next_rout_31_0_.m19_1_0\ : CFG4
      generic map(INIT => x"1B4E")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_0_rep2, C => m13, 
        D => pad_one_reg_0_0_a2_0, Y => m19_1_0);
    
    \next_rout_31_0_.m250_am_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => Kt_addr_4_rep1, B => m194, C => m85, Y => 
        m250_am_1);
    
    \next_rout_31_0_.m20\ : CFG4
      generic map(INIT => x"C1CD")

      port map(A => \m10_bm\, B => \m20_1\, C => Kt_addr(5), D
         => \m10_am\, Y => Kt_data_0);
    
    \next_rout_31_0_.m30\ : CFG4
      generic map(INIT => x"6335")

      port map(A => Kt_addr_4_rep1, B => Kt_addr(2), C => 
        Kt_addr_0_rep2, D => Kt_addr(1), Y => m30);
    
    \next_rout_31_0_.m276_bm\ : CFG4
      generic map(INIT => x"5ABE")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m276_bm);
    
    \next_rout_31_0_.m83_bm\ : CFG4
      generic map(INIT => x"0938")

      port map(A => Kt_addr(1), B => Kt_addr_4_rep2, C => 
        Kt_addr(2), D => Kt_addr_0_rep2, Y => m83_bm);
    
    \next_rout_31_0_.m323\ : CFG4
      generic map(INIT => x"2044")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_4_rep1, C => 
        Kt_addr_0_rep2, D => Kt_addr(2), Y => m323);
    
    \next_rout_31_0_.m95_1_1\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr_3_rep1, B => m93, C => m91, Y => 
        m95_1_1);
    
    \next_rout_31_0_.m270\ : CFG4
      generic map(INIT => x"EBAB")

      port map(A => m270_2, B => m270_1_1, C => Kt_addr(5), D => 
        m266, Y => Kt_data_24);
    
    \next_rout_31_0_.m174\ : CFG3
      generic map(INIT => x"64")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep1, Y => m174);
    
    \next_rout_31_0_.m146\ : CFG3
      generic map(INIT => x"1B")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m146);
    
    \next_rout_31_0_.m273_1\ : CFG4
      generic map(INIT => x"0440")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(4), C => 
        Kt_addr(0), D => m15, Y => m273_0);
    
    \next_rout_31_0_.m68\ : CFG3
      generic map(INIT => x"3E")

      port map(A => Kt_addr_fast(0), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, Y => m68);
    
    \next_rout_31_0_.m114_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_4_rep1, B => m81, C => Kt_addr_3_rep1, 
        Y => m296_2);
    
    \next_rout_31_0_.m62_am_1_0\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr_fast(4), B => m54, C => m53, Y => 
        m62_am_1_0);
    
    \next_rout_31_0_.m144_bm\ : CFG4
      generic map(INIT => x"F5E4")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => m85, D
         => hash_control_st_reg_ns_i_0_a2_0(4), Y => m144_bm);
    
    \next_rout_31_0_.m316_1_1\ : CFG4
      generic map(INIT => x"3726")

      port map(A => Kt_addr_5_rep1, B => Kt_addr(3), C => m311, D
         => m310, Y => m316_1_1);
    
    \next_rout_31_0_.m304\ : CFG4
      generic map(INIT => x"FFDC")

      port map(A => Kt_addr(3), B => m304_2, C => m304_1_0, D => 
        m304_1, Y => m304);
    
    \next_rout_31_0_.m215_bm_1\ : CFG4
      generic map(INIT => x"01AB")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep2, D => m164, Y => m215_bm_1);
    
    \next_rout_31_0_.m325\ : CFG4
      generic map(INIT => x"04BF")

      port map(A => Kt_addr(3), B => Kt_addr(5), C => 
        \hash_control_st_reg_ns_i_0_a2_2[4]\, D => m325_1_1, Y
         => m325);
    
    \next_rout_31_0_.m254_1_1\ : CFG3
      generic map(INIT => x"72")

      port map(A => Kt_addr(4), B => m252, C => m232, Y => 
        m254_1_1);
    
    \next_rout_31_0_.m219\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => m127, B => Kt_addr(3), C => m219_1_2, D => 
        m51, Y => m219);
    
    \next_rout_31_0_.m91\ : CFG4
      generic map(INIT => x"774B")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m91);
    
    \next_rout_31_0_.m273_2\ : CFG3
      generic map(INIT => x"20")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(4), C => m81, Y
         => m273_1);
    
    \next_rout_31_0_.m16\ : CFG3
      generic map(INIT => x"67")

      port map(A => Kt_addr_fast(0), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, Y => m16);
    
    \next_rout_31_0_.m78_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_4_rep2, B => m76, C => Kt_addr_3_rep1, 
        Y => m78_2);
    
    \next_rout_31_0_.m110_bm\ : CFG3
      generic map(INIT => x"64")

      port map(A => Kt_addr_4_rep2, B => m2, C => 
        pad_one_reg_0_0_a2_0, Y => m110_bm);
    
    \next_rout_31_0_.m48_2\ : CFG3
      generic map(INIT => x"40")

      port map(A => Kt_addr_fast(4), B => m45, C => 
        Kt_addr_fast(3), Y => m48_1);
    
    \next_rout_31_0_.m85\ : CFG3
      generic map(INIT => x"59")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m85);
    
    \next_rout_31_0_.m325_1_0_1\ : CFG4
      generic map(INIT => x"5456")

      port map(A => Kt_addr_fast(4), B => Kt_addr_fast(3), C => 
        Kt_addr_1_rep1, D => Kt_addr_2_rep1, Y => m325_1_0_1);
    
    \next_rout_31_0_.m250_bm_1_0_1\ : CFG4
      generic map(INIT => x"523F")

      port map(A => Kt_addr_fast(4), B => Kt_addr_fast(0), C => 
        Kt_addr_2_rep1, D => Kt_addr_1_rep1, Y => m250_bm_1_0_1);
    
    \next_rout_31_0_.m81\ : CFG3
      generic map(INIT => x"1A")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m81);
    
    \next_rout_31_0_.m276_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m276_bm, C => m276_am, Y => 
        m276_ns);
    
    \next_rout_31_0_.m172_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m172_bm, C => m172_am, Y => 
        m172_ns);
    
    \next_rout_31_0_.m285_1_1_1\ : CFG4
      generic map(INIT => x"100E")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_3_rep1, C => 
        Kt_addr_0_rep2, D => Kt_addr_1_rep2, Y => m285_1_1_1);
    
    \next_rout_31_0_.m104_bm\ : CFG4
      generic map(INIT => x"FFAB")

      port map(A => m304_2, B => Kt_addr_3_rep2, C => m104_bm_1, 
        D => m103_1, Y => m104_bm);
    
    \next_rout_31_0_.m168_1_0_1\ : CFG4
      generic map(INIT => x"058B")

      port map(A => Kt_addr_fast(3), B => Kt_addr_4_rep1, C => 
        Kt_addr_2_rep2, D => Kt_addr_1_rep2, Y => m168_1_0_1);
    
    \next_rout_31_0_.m263\ : CFG4
      generic map(INIT => x"7840")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m263);
    
    \next_rout_31_0_.m300_am\ : CFG4
      generic map(INIT => x"6C6A")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m300_am);
    
    \next_rout_31_0_.m205\ : CFG4
      generic map(INIT => x"615F")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m205);
    
    \next_rout_31_0_.m46\ : CFG3
      generic map(INIT => x"1D")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m46);
    
    \next_rout_31_0_.m207_1_0_1\ : CFG4
      generic map(INIT => x"1C3A")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_3_rep1, C => 
        Kt_addr_0_rep2, D => Kt_addr_1_rep2, Y => m207_1_0_1);
    
    \next_rout_31_0_.m26\ : CFG4
      generic map(INIT => x"43A5")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => i2_mux);
    
    \next_rout_31_0_.m235_am\ : CFG4
      generic map(INIT => x"E4B1")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => m232, D
         => hash_control_st_reg_ns_i_0_a2_0(4), Y => m235_am);
    
    \next_rout_31_0_.m230_1_0\ : CFG4
      generic map(INIT => x"0B5B")

      port map(A => Kt_addr_4_rep2, B => m227, C => 
        Kt_addr_3_rep2, D => Kt_addr(1), Y => m230_1_1);
    
    \next_rout_31_0_.m316\ : CFG4
      generic map(INIT => x"EEAE")

      port map(A => m316_2, B => m316_1_1, C => Kt_addr(5), D => 
        m313, Y => m316);
    
    \next_rout_31_0_.m222_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m222_bm, B => Kt_addr(3), C => m222_am, Y => 
        m222_ns);
    
    \next_rout_31_0_.m191\ : CFG4
      generic map(INIT => x"14CE")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m191);
    
    \next_rout_31_0_.m148\ : CFG4
      generic map(INIT => x"3250")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_fast(4), C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m148);
    
    \next_rout_31_0_.m144_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m144_bm, B => Kt_addr(3), C => m144_am, Y => 
        m144_ns);
    
    \next_rout_31_0_.m296_1_1\ : CFG4
      generic map(INIT => x"4567")

      port map(A => Kt_addr(4), B => Kt_addr_3_rep2, C => m237, D
         => hash_control_st_reg_ns_i_0_a2_0(4), Y => m296_1_1);
    
    \next_rout_31_0_.m215_am\ : CFG4
      generic map(INIT => x"DDCD")

      port map(A => m215_am_1_0, B => m211_0, C => Kt_addr_4_rep2, 
        D => m209, Y => m215_am);
    
    \next_rout_31_0_.m138\ : CFG3
      generic map(INIT => x"5C")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep1, Y => m138);
    
    \next_rout_31_0_.m49_am_1_0\ : CFG4
      generic map(INIT => x"4657")

      port map(A => Kt_addr_fast(4), B => Kt_addr_fast(3), C => 
        m35, D => Kt_addr_1_rep1, Y => m49_am_1_0);
    
    \next_rout_31_0_.m222_am\ : CFG4
      generic map(INIT => x"A7F4")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m222_am);
    
    \next_rout_31_0_.m209\ : CFG3
      generic map(INIT => x"21")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m209);
    
    \next_rout_31_0_.m325_1_1\ : CFG3
      generic map(INIT => x"1D")

      port map(A => m325_1_0, B => Kt_addr_5_rep1, C => m323, Y
         => m325_1_1);
    
    \next_rout_31_0_.m90\ : CFG3
      generic map(INIT => x"53")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m90);
    
    \next_rout_31_0_.m195\ : CFG4
      generic map(INIT => x"596C")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m195);
    
    \next_rout_31_0_.m87\ : CFG4
      generic map(INIT => x"1B41")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m87);
    
    \next_rout_31_0_.m254_1_0\ : CFG4
      generic map(INIT => x"058D")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => m105, D => 
        m1, Y => m254_1_0);
    
    \next_rout_31_0_.m250_bm\ : CFG4
      generic map(INIT => x"20FD")

      port map(A => Kt_addr_3_rep2, B => Kt_addr_4_rep2, C => 
        m132, D => m250_bm_1_0, Y => m250_bm);
    
    \next_rout_31_0_.m181\ : CFG4
      generic map(INIT => x"2E11")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_4_rep1, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m181);
    
    \next_rout_31_0_.m129\ : CFG3
      generic map(INIT => x"72")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_0_rep1, C => 
        Kt_addr_1_rep1, Y => m129);
    
    \next_rout_31_0_.m29\ : CFG3
      generic map(INIT => x"54")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m29);
    
    \next_rout_31_0_.m242\ : CFG3
      generic map(INIT => x"38")

      port map(A => Kt_addr_fast(1), B => Kt_addr_fast(0), C => 
        Kt_addr_2_rep1, Y => m242);
    
    \next_rout_31_0_.m232\ : CFG3
      generic map(INIT => x"45")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m232);
    
    \next_rout_31_0_.m172_am\ : CFG4
      generic map(INIT => x"111B")

      port map(A => Kt_addr_4_rep2, B => m133, C => Kt_addr(2), D
         => Kt_addr(1), Y => m172_am);
    
    \next_rout_31_0_.m163\ : CFG4
      generic map(INIT => x"12AD")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_4_rep1, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m163);
    
    \next_rout_31_0_.m73\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => m73_1, B => Kt_addr(4), C => m73_1_0, D => 
        m73, Y => m73_0);
    
    \next_rout_31_0_.m215_am_1_0\ : CFG4
      generic map(INIT => x"3276")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_3_rep1, C => m53, 
        D => m92, Y => m215_am_1_0);
    
    \next_rout_31_0_.m185\ : CFG3
      generic map(INIT => x"87")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep1, Y => m185);
    
    \next_rout_31_0_.m164\ : CFG3
      generic map(INIT => x"4A")

      port map(A => Kt_addr_fast(1), B => Kt_addr_fast(0), C => 
        Kt_addr_2_rep1, Y => m164);
    
    \next_rout_31_0_.m300_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m300_bm, B => Kt_addr(3), C => m300_am, Y => 
        m300_ns);
    
    \next_rout_31_0_.m78_1_0\ : CFG4
      generic map(INIT => x"44E4")

      port map(A => Kt_addr_4_rep2, B => m28, C => Kt_addr(2), D
         => Kt_addr(1), Y => m78_1_0);
    
    \next_rout_31_0_.m127\ : CFG3
      generic map(INIT => x"36")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m127);
    
    \next_rout_31_0_.m270_3\ : CFG4
      generic map(INIT => x"0800")

      port map(A => Kt_addr_5_rep1, B => Kt_addr_3_rep2, C => 
        Kt_addr(4), D => m267, Y => m270_2);
    
    \next_rout_31_0_.m226_am\ : CFG4
      generic map(INIT => x"F4DE")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m226_am);
    
    \next_rout_31_0_.m28\ : CFG3
      generic map(INIT => x"68")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m28);
    
    \next_rout_31_0_.m304_1_0\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr(4), B => m216, C => m133, Y => 
        m304_1_0);
    
    \next_rout_31_0_.m137_am_1_0\ : CFG4
      generic map(INIT => x"3276")

      port map(A => Kt_addr_fast(3), B => Kt_addr_fast(4), C => 
        m126, D => m127, Y => m137_am_1_0);
    
    \next_rout_31_0_.m254\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr(3), B => m254_1_1, C => m254_1_0, Y
         => m254);
    
    \next_rout_31_0_.m62_bm\ : CFG4
      generic map(INIT => x"BE14")

      port map(A => Kt_addr_3_rep1, B => Kt_addr_0_rep2, C => 
        Kt_addr(1), D => m60, Y => m62_bm);
    
    \next_rout_31_0_.m258_am\ : CFG3
      generic map(INIT => x"38")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => m1, Y => 
        m258_am);
    
    \next_rout_31_0_.m222_bm\ : CFG3
      generic map(INIT => x"67")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => m42, Y
         => m222_bm);
    
    \next_rout_31_0_.m193\ : CFG4
      generic map(INIT => x"0301")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m193);
    
    \next_rout_31_0_.m141_2\ : CFG3
      generic map(INIT => x"10")

      port map(A => Kt_addr_4_rep2, B => m90, C => Kt_addr_3_rep1, 
        Y => m177_1);
    
    \next_rout_31_0_.m42\ : CFG2
      generic map(INIT => x"4")

      port map(A => Kt_addr_1_rep1, B => Kt_addr_2_rep1, Y => m42);
    
    \next_rout_31_0_.m194\ : CFG3
      generic map(INIT => x"1C")

      port map(A => Kt_addr_fast(0), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, Y => m194);
    
    \next_rout_31_0_.m54\ : CFG3
      generic map(INIT => x"14")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m54);
    
    \next_rout_31_0_.m53\ : CFG3
      generic map(INIT => x"25")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m53);
    
    \next_rout_31_0_.m281_bm\ : CFG3
      generic map(INIT => x"8B")

      port map(A => m51, B => Kt_addr(4), C => m15, Y => m281_bm);
    
    \next_rout_31_0_.m239_1_2\ : CFG4
      generic map(INIT => x"193B")

      port map(A => Kt_addr_4_rep2, B => Kt_addr_3_rep2, C => 
        m105, D => m227, Y => m239_1_2);
    
    \next_rout_31_0_.m267\ : CFG3
      generic map(INIT => x"42")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m267);
    
    \next_rout_31_0_.m63\ : CFG3
      generic map(INIT => x"4C")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m63);
    
    \next_rout_31_0_.m22\ : CFG3
      generic map(INIT => x"49")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m22);
    
    \next_rout_31_0_.m32\ : CFG4
      generic map(INIT => x"6745")

      port map(A => Kt_addr_4_rep1, B => Kt_addr(2), C => 
        Kt_addr_0_rep2, D => Kt_addr(1), Y => m32);
    
    \next_rout_31_0_.m73_2\ : CFG3
      generic map(INIT => x"40")

      port map(A => Kt_addr_4_rep2, B => m70, C => Kt_addr_3_rep1, 
        Y => m73_1);
    
    \next_rout_31_0_.m184\ : CFG4
      generic map(INIT => x"3882")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m184);
    
    \next_rout_31_0_.m226_bm\ : CFG4
      generic map(INIT => x"66A5")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(2), C => 
        pad_one_reg_0_0_a2_0, D => Kt_addr(0), Y => m226_bm);
    
    \next_rout_31_0_.m124_1_2\ : CFG4
      generic map(INIT => x"2367")

      port map(A => Kt_addr_4_rep2, B => Kt_addr_3_rep2, C => 
        m120, D => m122, Y => m124_1_2);
    
    \next_rout_31_0_.m180\ : CFG4
      generic map(INIT => x"270D")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_4_rep1, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m180);
    
    \next_rout_31_0_.m289_1_1\ : CFG4
      generic map(INIT => x"4E5F")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => m37, D => 
        m1, Y => m289_1_1);
    
    \next_rout_31_0_.m308_ns_1\ : CFG4
      generic map(INIT => x"33B1")

      port map(A => Kt_addr(4), B => Kt_addr(1), C => m1, D => 
        Kt_addr(0), Y => m308_ns_1);
    
    \next_rout_31_0_.m1\ : CFG2
      generic map(INIT => x"9")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, Y => m1);
    
    \next_rout_31_0_.m311\ : CFG4
      generic map(INIT => x"6521")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_4_rep1, C => 
        Kt_addr_0_rep2, D => Kt_addr(2), Y => m311);
    
    \next_rout_31_0_.m19_1_1\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr_4_rep1, B => m17, C => m16, Y => 
        m19_1_1);
    
    \next_rout_31_0_.m124\ : CFG4
      generic map(INIT => x"4F43")

      port map(A => m90, B => Kt_addr(4), C => m124_1_2, D => m16, 
        Y => m124);
    
    \next_rout_31_0_.m20_1\ : CFG4
      generic map(INIT => x"3B19")

      port map(A => Kt_addr_5_rep1, B => Kt_addr_3_rep2, C => 
        m19_1_1, D => m19_1_0, Y => \m20_1\);
    
    \next_rout_31_0_.m73_1_0\ : CFG4
      generic map(INIT => x"41EB")

      port map(A => Kt_addr_3_rep1, B => Kt_addr_0_rep2, C => 
        Kt_addr(1), D => m71, Y => m73_1_0);
    
    \next_rout_31_0_.m120\ : CFG3
      generic map(INIT => x"23")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m120);
    
    \next_rout_31_0_.m281_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m281_bm, C => m281_am, Y => 
        m281_ns);
    
    \next_rout_31_0_.m49_bm_1\ : CFG4
      generic map(INIT => x"0A4E")

      port map(A => Kt_addr_fast(4), B => Kt_addr_0_rep1, C => 
        m43, D => hash_control_st_reg_ns_i_0_a2_0(4), Y => 
        m49_bm_1);
    
    \next_rout_31_0_.m122\ : CFG3
      generic map(INIT => x"1C")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_0_rep1, C => 
        Kt_addr_1_rep1, Y => m122);
    
    \next_rout_31_0_.m285\ : CFG4
      generic map(INIT => x"02DF")

      port map(A => Kt_addr(3), B => Kt_addr(4), C => m28, D => 
        m285_1_1, Y => m285);
    
    \next_rout_31_0_.m252\ : CFG3
      generic map(INIT => x"2A")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m252);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity gv_sha256 is

    port( sha256_controller_0_bytes_o  : in    std_logic_vector(1 to 1);
          raddr_pos                    : in    std_logic_vector(3 downto 2);
          SHA256_BLOCK_0_H0_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o          : out   std_logic_vector(31 downto 0);
          state_2                      : in    std_logic;
          state_0                      : in    std_logic;
          state_3                      : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK : in    std_logic;
          SHA256_Module_0_di_req_o     : out   std_logic;
          SHA256_Module_0_do_valid_o   : out   std_logic;
          sha256_controller_0_end_o    : in    std_logic;
          last_block_0                 : in    std_logic;
          ce_i_i_2                     : in    std_logic;
          N_28                         : in    std_logic;
          SHA256_Module_0_error_o      : out   std_logic;
          N_1696                       : in    std_logic;
          N_1400                       : in    std_logic;
          N_1624                       : in    std_logic;
          N_920                        : in    std_logic;
          N_1144                       : in    std_logic;
          N_1399                       : in    std_logic;
          N_1623                       : in    std_logic;
          N_919                        : in    std_logic;
          N_1143                       : in    std_logic;
          N_1401                       : in    std_logic;
          N_1625                       : in    std_logic;
          N_921                        : in    std_logic;
          N_1145                       : in    std_logic;
          ren_pos                      : in    std_logic;
          N_1694                       : in    std_logic;
          N_1692                       : in    std_logic;
          N_1693                       : in    std_logic;
          N_1691                       : in    std_logic;
          N_1690                       : in    std_logic;
          N_89                         : in    std_logic;
          N_1695                       : in    std_logic;
          N_1708                       : in    std_logic;
          N_1709                       : in    std_logic;
          N_1707                       : in    std_logic;
          N_1706                       : in    std_logic;
          N_1705                       : in    std_logic;
          N_1704                       : in    std_logic;
          N_1703                       : in    std_logic;
          N_1700                       : in    std_logic;
          N_1701                       : in    std_logic;
          N_1697                       : in    std_logic;
          N_1699                       : in    std_logic;
          N_1698                       : in    std_logic;
          N_1717                       : in    std_logic;
          N_1712                       : in    std_logic;
          N_1716                       : in    std_logic;
          N_1715                       : in    std_logic;
          N_1711                       : in    std_logic;
          N_1713                       : in    std_logic;
          N_1714                       : in    std_logic;
          N_1718                       : in    std_logic;
          N_1702                       : in    std_logic;
          N_1710                       : in    std_logic
        );

end gv_sha256;

architecture DEF_ARCH of gv_sha256 is 

  component sha256_control
    port( hash_control_st_reg_i           : out   std_logic_vector(6 to 6);
          msg_bitlen                      : out   std_logic_vector(63 downto 3);
          Kt_addr                         : out   std_logic_vector(5 downto 0);
          st_cnt_reg                      : out   std_logic_vector(6 to 6);
          Kt_addr_fast                    : out   std_logic_vector(5 downto 0);
          sha256_controller_0_bytes_o     : in    std_logic_vector(1 to 1) := (others => 'U');
          hash_control_st_reg_ns_i_0_a2_0 : out   std_logic_vector(4 to 4);
          hash_control_st_reg_ns_i_0_a2_2 : in    std_logic_vector(4 to 4) := (others => 'U');
          hash_control_st_reg_2           : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK    : in    std_logic := 'U';
          one_insert                      : out   std_logic;
          sha_last_blk_reg                : out   std_logic;
          SHA256_Module_0_di_req_o        : out   std_logic;
          SHA256_Module_0_do_valid_o      : out   std_logic;
          Kt_addr_2_rep1                  : out   std_logic;
          Kt_addr_2_rep2                  : out   std_logic;
          Kt_addr_1_rep1                  : out   std_logic;
          Kt_addr_1_rep2                  : out   std_logic;
          Kt_addr_3_rep1                  : out   std_logic;
          Kt_addr_3_rep2                  : out   std_logic;
          Kt_addr_5_rep1                  : out   std_logic;
          Kt_addr_0_rep1                  : out   std_logic;
          Kt_addr_0_rep2                  : out   std_logic;
          Kt_addr_4_rep1                  : out   std_logic;
          Kt_addr_4_rep2                  : out   std_logic;
          sha256_controller_0_end_o       : in    std_logic := 'U';
          last_block_0                    : in    std_logic := 'U';
          N_168_i_0                       : out   std_logic;
          ce_i_i_2                        : in    std_logic := 'U';
          pad_one_reg_0_0_a2_0            : out   std_logic;
          sha_last_blk_next_0_o2_0        : out   std_logic;
          oregs_ce_i_a2_0_a2              : out   std_logic;
          N_102                           : out   std_logic;
          N_28                            : in    std_logic := 'U';
          N_387                           : out   std_logic;
          N_388                           : in    std_logic := 'U';
          W_m4_e_2                        : in    std_logic := 'U';
          N_105                           : in    std_logic := 'U';
          N_111                           : out   std_logic;
          core_ce_o_iv_i_0                : out   std_logic;
          N_244_i_0                       : out   std_logic;
          SHA256_Module_0_error_o         : out   std_logic;
          ld_i_i_3                        : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component sha256_hash_core
    port( R1_data                      : out   std_logic_vector(31 downto 0);
          R2_data                      : out   std_logic_vector(31 downto 0);
          R3_data                      : out   std_logic_vector(31 downto 0);
          R5_data                      : out   std_logic_vector(31 downto 0);
          R6_data                      : out   std_logic_vector(31 downto 0);
          R7_data                      : out   std_logic_vector(31 downto 0);
          R0_data                      : out   std_logic_vector(31 downto 0);
          R4_data                      : out   std_logic_vector(31 downto 0);
          N4_data                      : in    std_logic_vector(31 downto 1) := (others => 'U');
          N0_data                      : in    std_logic_vector(31 downto 1) := (others => 'U');
          W_out_i_0                    : in    std_logic_vector(0 to 0) := (others => 'U');
          Kt_addr                      : in    std_logic_vector(5 to 5) := (others => 'U');
          N3_data                      : in    std_logic_vector(31 downto 1) := (others => 'U');
          N2_data                      : in    std_logic_vector(31 downto 1) := (others => 'U');
          N1_data                      : in    std_logic_vector(31 downto 1) := (others => 'U');
          N7_data                      : in    std_logic_vector(31 downto 1) := (others => 'U');
          N6_data                      : in    std_logic_vector(31 downto 1) := (others => 'U');
          N5_data                      : in    std_logic_vector(31 downto 1) := (others => 'U');
          Wt_data                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          Kt_data_15                   : in    std_logic := 'U';
          Kt_data_24                   : in    std_logic := 'U';
          Kt_data_0                    : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK : in    std_logic := 'U';
          core_ce_o_iv_i_0             : in    std_logic := 'U';
          oregs_ce_i_a2_0_a2           : in    std_logic := 'U';
          next_reg_H4_cry_0_0_Y        : in    std_logic := 'U';
          next_reg_H0_cry_0_0_Y        : in    std_logic := 'U';
          next_r0_0_cry_0_Y            : in    std_logic := 'U';
          ld_i_i_3                     : in    std_logic := 'U';
          N_98                         : in    std_logic := 'U';
          m10_bm                       : in    std_logic := 'U';
          m20_1                        : in    std_logic := 'U';
          m10_am                       : in    std_logic := 'U';
          m34                          : in    std_logic := 'U';
          m49_am                       : in    std_logic := 'U';
          m49_bm                       : in    std_logic := 'U';
          Kt_addr_5_rep1               : in    std_logic := 'U';
          m62_am                       : in    std_logic := 'U';
          m62_bm                       : in    std_logic := 'U';
          m67_ns                       : in    std_logic := 'U';
          m73                          : in    std_logic := 'U';
          m78                          : in    std_logic := 'U';
          m83_ns                       : in    std_logic := 'U';
          m95_1_0                      : in    std_logic := 'U';
          m95_1_1                      : in    std_logic := 'U';
          m104_am                      : in    std_logic := 'U';
          m104_bm                      : in    std_logic := 'U';
          m110_ns                      : in    std_logic := 'U';
          m114                         : in    std_logic := 'U';
          m119_ns                      : in    std_logic := 'U';
          m124                         : in    std_logic := 'U';
          m137_am                      : in    std_logic := 'U';
          m137_bm                      : in    std_logic := 'U';
          m141                         : in    std_logic := 'U';
          m144_ns                      : in    std_logic := 'U';
          m157                         : in    std_logic := 'U';
          m168_1_0                     : in    std_logic := 'U';
          m168_1_1                     : in    std_logic := 'U';
          m172_ns                      : in    std_logic := 'U';
          m177                         : in    std_logic := 'U';
          m197_1_0                     : in    std_logic := 'U';
          m197_1_1                     : in    std_logic := 'U';
          m207_1_0                     : in    std_logic := 'U';
          m207_1_1                     : in    std_logic := 'U';
          m215_am                      : in    std_logic := 'U';
          m215_bm                      : in    std_logic := 'U';
          m219                         : in    std_logic := 'U';
          m222_ns                      : in    std_logic := 'U';
          m226_ns                      : in    std_logic := 'U';
          m230                         : in    std_logic := 'U';
          m235_ns                      : in    std_logic := 'U';
          m239                         : in    std_logic := 'U';
          m250_am                      : in    std_logic := 'U';
          m250_bm                      : in    std_logic := 'U';
          m254                         : in    std_logic := 'U';
          m258_ns                      : in    std_logic := 'U';
          m273                         : in    std_logic := 'U';
          m276_ns                      : in    std_logic := 'U';
          m281_ns                      : in    std_logic := 'U';
          m285                         : in    std_logic := 'U';
          m289                         : in    std_logic := 'U';
          m292_ns                      : in    std_logic := 'U';
          m296                         : in    std_logic := 'U';
          m300_ns                      : in    std_logic := 'U';
          m304                         : in    std_logic := 'U';
          i3_mux_1                     : in    std_logic := 'U';
          m325                         : in    std_logic := 'U';
          m316                         : in    std_logic := 'U';
          next_reg_H3_cry_0_0_Y        : in    std_logic := 'U';
          next_reg_H2_cry_0_0_Y        : in    std_logic := 'U';
          next_reg_H1_cry_0_0_Y        : in    std_logic := 'U';
          next_reg_H7_cry_0_0_Y        : in    std_logic := 'U';
          next_reg_H6_cry_0_0_Y        : in    std_logic := 'U';
          next_reg_H5_cry_0_0_Y        : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component sha256_regs
    port( SHA256_BLOCK_0_H0_o          : out   std_logic_vector(31 downto 0);
          N0_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H1_o          : out   std_logic_vector(31 downto 0);
          N1_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H2_o          : out   std_logic_vector(31 downto 0);
          N2_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H3_o          : out   std_logic_vector(31 downto 0);
          N3_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H4_o          : out   std_logic_vector(31 downto 0);
          N4_data                      : out   std_logic_vector(31 downto 1);
          N5_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H5_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o          : out   std_logic_vector(31 downto 0);
          N6_data                      : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H7_o          : out   std_logic_vector(31 downto 0);
          N7_data                      : out   std_logic_vector(31 downto 1);
          hash_control_st_reg_i        : in    std_logic_vector(6 to 6) := (others => 'U');
          R0_data                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          R1_data                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          R2_data                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          R3_data                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          R4_data                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          R5_data                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          R6_data                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          R7_data                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          sha256_system_sb_0_FIC_0_CLK : in    std_logic := 'U';
          N_168_i_0                    : in    std_logic := 'U';
          next_reg_H0_cry_0_0_Y        : out   std_logic;
          next_reg_H1_cry_0_0_Y        : out   std_logic;
          next_reg_H2_cry_0_0_Y        : out   std_logic;
          next_reg_H3_cry_0_0_Y        : out   std_logic;
          next_reg_H4_cry_0_0_Y        : out   std_logic;
          next_reg_H5_cry_0_0_Y        : out   std_logic;
          next_reg_H6_cry_0_0_Y        : out   std_logic;
          next_reg_H7_cry_0_0_Y        : out   std_logic
        );
  end component;

  component sha256_padding
    port( raddr_pos                   : in    std_logic_vector(3 downto 2) := (others => 'U');
          Kt_addr                     : in    std_logic_vector(0 to 0) := (others => 'U');
          st_cnt_reg                  : in    std_logic_vector(6 to 6) := (others => 'U');
          hash_control_st_reg         : in    std_logic_vector(2 to 2) := (others => 'U');
          Kt_addr_fast                : in    std_logic_vector(5 downto 2) := (others => 'U');
          sha256_controller_0_bytes_o : in    std_logic_vector(1 to 1) := (others => 'U');
          W_out_2_0                   : out   std_logic_vector(5 to 5);
          W_out_i_0                   : out   std_logic_vector(2 downto 0);
          W_out_i_i_1_1               : out   std_logic_vector(31 to 31);
          W_out_2_0_1                 : out   std_logic_vector(7 to 7);
          W_out_i_i_1                 : out   std_logic_vector(31 to 31);
          W_out_2_0_a4_1_0_RNIFI1DA   : out   std_logic_vector(23 to 23);
          W_out_2_0_a4_1_0_RNI32U7B   : out   std_logic_vector(23 to 23);
          msg_bitlen                  : in    std_logic_vector(63 downto 3) := (others => 'U');
          state_2                     : in    std_logic := 'U';
          state_0                     : in    std_logic := 'U';
          state_3                     : in    std_logic := 'U';
          W_out_2_0_0_20              : out   std_logic;
          W_out_2_0_0_12              : out   std_logic;
          W_out_2_0_0_4               : out   std_logic;
          W_out_2_0_0_1               : out   std_logic;
          W_out_2_0_0_3               : out   std_logic;
          W_out_2_0_0_0               : out   std_logic;
          W_out_2_i_0_22              : out   std_logic;
          W_out_2_i_0_17              : out   std_logic;
          W_out_2_i_0_21              : out   std_logic;
          W_out_2_i_0_20              : out   std_logic;
          W_out_2_i_0_16              : out   std_logic;
          W_out_2_i_0_18              : out   std_logic;
          W_out_2_i_0_19              : out   std_logic;
          W_out_2_i_2_0               : out   std_logic;
          W_out_2_i_2_5               : out   std_logic;
          W_out_2_i_2_6               : out   std_logic;
          W_out_2_i_1_1               : out   std_logic;
          W_out_2_i_1_0               : out   std_logic;
          W_out_2_i_1_22              : out   std_logic;
          W_out_2_i_1_17              : out   std_logic;
          W_out_2_i_1_21              : out   std_logic;
          W_out_2_i_1_20              : out   std_logic;
          W_out_2_i_1_16              : out   std_logic;
          W_out_2_i_1_18              : out   std_logic;
          W_out_2_i_1_19              : out   std_logic;
          W_out_2_i_1_13              : out   std_logic;
          W_out_2_i_1_10              : out   std_logic;
          W_out_2_i_1_12              : out   std_logic;
          W_out_2_i_1_14              : out   std_logic;
          W_out_2_i_1_9               : out   std_logic;
          W_out_2_i_1_11              : out   std_logic;
          W_out_2_i_1_8               : out   std_logic;
          W_out_2_i_1_2               : out   std_logic;
          W_out_2_i_1_4               : out   std_logic;
          W_out_2_i_1_3               : out   std_logic;
          N_1696                      : in    std_logic := 'U';
          SHA256_Module_0_di_req_o    : in    std_logic := 'U';
          N_1400                      : in    std_logic := 'U';
          N_1624                      : in    std_logic := 'U';
          N_920                       : in    std_logic := 'U';
          N_1144                      : in    std_logic := 'U';
          N_1399                      : in    std_logic := 'U';
          N_1623                      : in    std_logic := 'U';
          N_919                       : in    std_logic := 'U';
          N_1143                      : in    std_logic := 'U';
          N_1401                      : in    std_logic := 'U';
          N_1625                      : in    std_logic := 'U';
          N_921                       : in    std_logic := 'U';
          N_1145                      : in    std_logic := 'U';
          one_insert                  : in    std_logic := 'U';
          N_388                       : out   std_logic;
          W_m4_e_2                    : out   std_logic;
          Kt_addr_1_rep1              : in    std_logic := 'U';
          N_102                       : in    std_logic := 'U';
          N_105                       : out   std_logic;
          ren_pos                     : in    std_logic := 'U';
          sha256_controller_0_end_o   : in    std_logic := 'U';
          Kt_addr_0_rep2              : in    std_logic := 'U';
          sha_last_blk_reg            : in    std_logic := 'U';
          sha_last_blk_next_0_o2_0    : in    std_logic := 'U';
          N_387                       : in    std_logic := 'U';
          N_98                        : out   std_logic;
          N_111                       : in    std_logic := 'U';
          N_1694                      : in    std_logic := 'U';
          N_1692                      : in    std_logic := 'U';
          N_349                       : out   std_logic;
          N_1693                      : in    std_logic := 'U';
          N_251                       : out   std_logic;
          N_1691                      : in    std_logic := 'U';
          N_248                       : out   std_logic;
          N_1690                      : in    std_logic := 'U';
          N_245                       : out   std_logic;
          N_89                        : in    std_logic := 'U';
          N_1695                      : in    std_logic := 'U';
          N_1708                      : in    std_logic := 'U';
          N_1709                      : in    std_logic := 'U';
          N_1707                      : in    std_logic := 'U';
          N_1706                      : in    std_logic := 'U';
          N_1705                      : in    std_logic := 'U';
          N_1704                      : in    std_logic := 'U';
          N_1703                      : in    std_logic := 'U';
          N_1700                      : in    std_logic := 'U';
          N_1701                      : in    std_logic := 'U';
          N_1697                      : in    std_logic := 'U';
          N_1699                      : in    std_logic := 'U';
          N_1698                      : in    std_logic := 'U';
          N_1717                      : in    std_logic := 'U';
          N_1712                      : in    std_logic := 'U';
          N_1716                      : in    std_logic := 'U';
          N_1715                      : in    std_logic := 'U';
          N_1711                      : in    std_logic := 'U';
          N_1713                      : in    std_logic := 'U';
          N_1714                      : in    std_logic := 'U';
          N_1718                      : in    std_logic := 'U';
          N_1702                      : in    std_logic := 'U';
          N_1710                      : in    std_logic := 'U';
          N_263                       : out   std_logic;
          N_301                       : out   std_logic;
          N_304                       : out   std_logic;
          N_298                       : out   std_logic;
          N_295                       : out   std_logic;
          N_292                       : out   std_logic;
          N_289                       : out   std_logic;
          N_286                       : out   std_logic;
          N_278                       : out   std_logic;
          N_275                       : out   std_logic;
          N_272                       : out   std_logic;
          N_268                       : out   std_logic;
          N_265                       : out   std_logic
        );
  end component;

  component sha256_msg_sch
    port( Wt_data                      : out   std_logic_vector(31 downto 0);
          W_out_2_0                    : in    std_logic_vector(5 to 5) := (others => 'U');
          W_out_i_0                    : in    std_logic_vector(2 downto 0) := (others => 'U');
          W_out_i_i_1_1                : in    std_logic_vector(31 to 31) := (others => 'U');
          W_out_i_i_1                  : in    std_logic_vector(31 to 31) := (others => 'U');
          W_out_2_i_0                  : in    std_logic_vector(30 downto 24) := (others => 'U');
          W_out_2_0_a4_1_0_RNI32U7B    : in    std_logic_vector(23 to 23) := (others => 'U');
          W_out_2_0_a4_1_0_RNIFI1DA    : in    std_logic_vector(23 to 23) := (others => 'U');
          W_out_2_0_1                  : in    std_logic_vector(7 to 7) := (others => 'U');
          W_out_2_0_0_3                : in    std_logic := 'U';
          W_out_2_0_0_1                : in    std_logic := 'U';
          W_out_2_0_0_0                : in    std_logic := 'U';
          W_out_2_0_0_20               : in    std_logic := 'U';
          W_out_2_0_0_12               : in    std_logic := 'U';
          W_out_2_0_0_4                : in    std_logic := 'U';
          W_out_2_i_2_0                : in    std_logic := 'U';
          W_out_2_i_2_6                : in    std_logic := 'U';
          W_out_2_i_2_5                : in    std_logic := 'U';
          W_out_2_i_1_22               : in    std_logic := 'U';
          W_out_2_i_1_21               : in    std_logic := 'U';
          W_out_2_i_1_20               : in    std_logic := 'U';
          W_out_2_i_1_19               : in    std_logic := 'U';
          W_out_2_i_1_18               : in    std_logic := 'U';
          W_out_2_i_1_17               : in    std_logic := 'U';
          W_out_2_i_1_16               : in    std_logic := 'U';
          W_out_2_i_1_0                : in    std_logic := 'U';
          W_out_2_i_1_14               : in    std_logic := 'U';
          W_out_2_i_1_13               : in    std_logic := 'U';
          W_out_2_i_1_12               : in    std_logic := 'U';
          W_out_2_i_1_11               : in    std_logic := 'U';
          W_out_2_i_1_10               : in    std_logic := 'U';
          W_out_2_i_1_9                : in    std_logic := 'U';
          W_out_2_i_1_8                : in    std_logic := 'U';
          W_out_2_i_1_4                : in    std_logic := 'U';
          W_out_2_i_1_3                : in    std_logic := 'U';
          W_out_2_i_1_2                : in    std_logic := 'U';
          W_out_2_i_1_1                : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK : in    std_logic := 'U';
          N_244_i_0                    : in    std_logic := 'U';
          next_r0_0_cry_0_Y            : out   std_logic;
          N_251                        : in    std_logic := 'U';
          ld_i_i_3                     : in    std_logic := 'U';
          N_349                        : in    std_logic := 'U';
          N_248                        : in    std_logic := 'U';
          N_245                        : in    std_logic := 'U';
          N_98                         : in    std_logic := 'U';
          N_304                        : in    std_logic := 'U';
          N_301                        : in    std_logic := 'U';
          N_298                        : in    std_logic := 'U';
          N_295                        : in    std_logic := 'U';
          N_292                        : in    std_logic := 'U';
          N_289                        : in    std_logic := 'U';
          N_286                        : in    std_logic := 'U';
          N_278                        : in    std_logic := 'U';
          N_275                        : in    std_logic := 'U';
          N_272                        : in    std_logic := 'U';
          N_268                        : in    std_logic := 'U';
          N_265                        : in    std_logic := 'U';
          N_263                        : in    std_logic := 'U'
        );
  end component;

  component sha256_kt_rom
    port( hash_control_st_reg_ns_i_0_a2_0 : in    std_logic_vector(4 to 4) := (others => 'U');
          hash_control_st_reg_ns_i_0_a2_2 : out   std_logic_vector(4 to 4);
          Kt_addr                         : in    std_logic_vector(5 downto 0) := (others => 'U');
          Kt_addr_fast                    : in    std_logic_vector(4 downto 0) := (others => 'U');
          Kt_data_0                       : out   std_logic;
          Kt_data_24                      : out   std_logic;
          Kt_data_15                      : out   std_logic;
          m10_bm                          : out   std_logic;
          m20_1                           : out   std_logic;
          m10_am                          : out   std_logic;
          Kt_addr_5_rep1                  : in    std_logic := 'U';
          Kt_addr_3_rep2                  : in    std_logic := 'U';
          Kt_addr_3_rep1                  : in    std_logic := 'U';
          m62_am                          : out   std_logic;
          Kt_addr_0_rep1                  : in    std_logic := 'U';
          m104_bm                         : out   std_logic;
          Kt_addr_2_rep1                  : in    std_logic := 'U';
          Kt_addr_0_rep2                  : in    std_logic := 'U';
          m49_am                          : out   std_logic;
          Kt_addr_1_rep1                  : in    std_logic := 'U';
          m49_bm                          : out   std_logic;
          m137_am                         : out   std_logic;
          m137_bm                         : out   std_logic;
          Kt_addr_2_rep2                  : in    std_logic := 'U';
          Kt_addr_1_rep2                  : in    std_logic := 'U';
          Kt_addr_4_rep2                  : in    std_logic := 'U';
          m215_am                         : out   std_logic;
          Kt_addr_4_rep1                  : in    std_logic := 'U';
          m215_bm                         : out   std_logic;
          m250_am                         : out   std_logic;
          m250_bm                         : out   std_logic;
          m207_1_1                        : out   std_logic;
          m207_1_0                        : out   std_logic;
          m95_1_1                         : out   std_logic;
          m95_1_0                         : out   std_logic;
          m197_1_1                        : out   std_logic;
          m197_1_0                        : out   std_logic;
          m316                            : out   std_logic;
          m34                             : out   std_logic;
          m157                            : out   std_logic;
          m325                            : out   std_logic;
          m168_1_1                        : out   std_logic;
          m168_1_0                        : out   std_logic;
          m230                            : out   std_logic;
          m296                            : out   std_logic;
          m254                            : out   std_logic;
          m114                            : out   std_logic;
          m304                            : out   std_logic;
          m73_0                           : out   std_logic;
          pad_one_reg_0_0_a2_0            : in    std_logic := 'U';
          m239                            : out   std_logic;
          m219                            : out   std_logic;
          m285                            : out   std_logic;
          m177                            : out   std_logic;
          m124                            : out   std_logic;
          m289                            : out   std_logic;
          m78                             : out   std_logic;
          m141                            : out   std_logic;
          i3_mux_1                        : out   std_logic;
          m67_ns                          : out   std_logic;
          m83_ns                          : out   std_logic;
          m110_ns                         : out   std_logic;
          m119_ns                         : out   std_logic;
          m144_ns                         : out   std_logic;
          m172_ns                         : out   std_logic;
          m222_ns                         : out   std_logic;
          m226_ns                         : out   std_logic;
          m235_ns                         : out   std_logic;
          m258_ns                         : out   std_logic;
          m276_ns                         : out   std_logic;
          m281_ns                         : out   std_logic;
          m292_ns                         : out   std_logic;
          m300_ns                         : out   std_logic;
          m273                            : out   std_logic;
          m104_am                         : out   std_logic;
          m62_bm                          : out   std_logic
        );
  end component;

    signal \hash_control_st_reg_i[6]\, \msg_bitlen[3]\, 
        \msg_bitlen[4]\, \msg_bitlen[5]\, \msg_bitlen[6]\, 
        \msg_bitlen[7]\, \msg_bitlen[8]\, \msg_bitlen[9]\, 
        \msg_bitlen[10]\, \msg_bitlen[11]\, \msg_bitlen[12]\, 
        \msg_bitlen[13]\, \msg_bitlen[14]\, \msg_bitlen[15]\, 
        \msg_bitlen[16]\, \msg_bitlen[17]\, \msg_bitlen[18]\, 
        \msg_bitlen[19]\, \msg_bitlen[20]\, \msg_bitlen[21]\, 
        \msg_bitlen[22]\, \msg_bitlen[23]\, \msg_bitlen[24]\, 
        \msg_bitlen[25]\, \msg_bitlen[26]\, \msg_bitlen[27]\, 
        \msg_bitlen[28]\, \msg_bitlen[29]\, \msg_bitlen[30]\, 
        \msg_bitlen[31]\, \msg_bitlen[32]\, \msg_bitlen[33]\, 
        \msg_bitlen[34]\, \msg_bitlen[35]\, \msg_bitlen[36]\, 
        \msg_bitlen[37]\, \msg_bitlen[38]\, \msg_bitlen[39]\, 
        \msg_bitlen[40]\, \msg_bitlen[41]\, \msg_bitlen[42]\, 
        \msg_bitlen[43]\, \msg_bitlen[44]\, \msg_bitlen[45]\, 
        \msg_bitlen[46]\, \msg_bitlen[47]\, \msg_bitlen[48]\, 
        \msg_bitlen[49]\, \msg_bitlen[50]\, \msg_bitlen[51]\, 
        \msg_bitlen[52]\, \msg_bitlen[53]\, \msg_bitlen[54]\, 
        \msg_bitlen[55]\, \msg_bitlen[56]\, \msg_bitlen[57]\, 
        \msg_bitlen[58]\, \msg_bitlen[59]\, \msg_bitlen[60]\, 
        \msg_bitlen[61]\, \msg_bitlen[62]\, \msg_bitlen[63]\, 
        \Kt_addr[0]\, \Kt_addr[1]\, \Kt_addr[2]\, \Kt_addr[3]\, 
        \Kt_addr[4]\, \Kt_addr[5]\, \st_cnt_reg[6]\, 
        \hash_control_st_reg[2]\, \Kt_addr_fast[0]\, 
        \Kt_addr_fast[1]\, \Kt_addr_fast[2]\, \Kt_addr_fast[3]\, 
        \Kt_addr_fast[4]\, \Kt_addr_fast[5]\, 
        \hash_control_st_reg_ns_i_0_a2_0[4]\, 
        \hash_control_st_reg_ns_i_0_a2_2[4]\, one_insert, 
        sha_last_blk_reg, \SHA256_Module_0_di_req_o\, 
        Kt_addr_2_rep1, Kt_addr_2_rep2, Kt_addr_1_rep1, 
        Kt_addr_1_rep2, Kt_addr_3_rep1, Kt_addr_3_rep2, 
        Kt_addr_5_rep1, Kt_addr_0_rep1, Kt_addr_0_rep2, 
        Kt_addr_4_rep1, Kt_addr_4_rep2, N_168_i_0, 
        pad_one_reg_0_0_a2_0, sha_last_blk_next_0_o2_0, 
        oregs_ce_i_a2_0_a2, N_102, N_387, N_388, W_m4_e_2, N_105, 
        N_111, core_ce_o_iv_i_0, N_244_i_0, ld_i_i_3, 
        \W_out_2_0[5]\, \W_out_2_0_0[23]\, \W_out_2_0_0[15]\, 
        \W_out_2_0_0[7]\, \W_out_2_0_0[4]\, \W_out_2_0_0[6]\, 
        \W_out_2_0_0[3]\, \W_out_2_i_0[30]\, \W_out_2_i_0[25]\, 
        \W_out_2_i_0[29]\, \W_out_2_i_0[28]\, \W_out_2_i_0[24]\, 
        \W_out_2_i_0[26]\, \W_out_2_i_0[27]\, \W_out_i_0[0]\, 
        \W_out_i_0[1]\, \W_out_i_0[2]\, \W_out_i_i_1_1[31]\, 
        \W_out_2_0_1[7]\, \W_out_i_i_1[31]\, 
        \W_out_2_0_a4_1_0_RNIFI1DA[23]\, 
        \W_out_2_0_a4_1_0_RNI32U7B[23]\, \W_out_2_i_2[8]\, 
        \W_out_2_i_2[13]\, \W_out_2_i_2[14]\, \W_out_2_i_1[9]\, 
        \W_out_2_i_1[8]\, \W_out_2_i_1[30]\, \W_out_2_i_1[25]\, 
        \W_out_2_i_1[29]\, \W_out_2_i_1[28]\, \W_out_2_i_1[24]\, 
        \W_out_2_i_1[26]\, \W_out_2_i_1[27]\, \W_out_2_i_1[21]\, 
        \W_out_2_i_1[18]\, \W_out_2_i_1[20]\, \W_out_2_i_1[22]\, 
        \W_out_2_i_1[17]\, \W_out_2_i_1[19]\, \W_out_2_i_1[16]\, 
        \W_out_2_i_1[10]\, \W_out_2_i_1[12]\, \W_out_2_i_1[11]\, 
        N_98, N_349, N_251, N_248, N_245, N_263, N_301, N_304, 
        N_298, N_295, N_292, N_289, N_286, N_278, N_275, N_272, 
        N_268, N_265, \Wt_data[0]\, \Wt_data[1]\, \Wt_data[2]\, 
        \Wt_data[3]\, \Wt_data[4]\, \Wt_data[5]\, \Wt_data[6]\, 
        \Wt_data[7]\, \Wt_data[8]\, \Wt_data[9]\, \Wt_data[10]\, 
        \Wt_data[11]\, \Wt_data[12]\, \Wt_data[13]\, 
        \Wt_data[14]\, \Wt_data[15]\, \Wt_data[16]\, 
        \Wt_data[17]\, \Wt_data[18]\, \Wt_data[19]\, 
        \Wt_data[20]\, \Wt_data[21]\, \Wt_data[22]\, 
        \Wt_data[23]\, \Wt_data[24]\, \Wt_data[25]\, 
        \Wt_data[26]\, \Wt_data[27]\, \Wt_data[28]\, 
        \Wt_data[29]\, \Wt_data[30]\, \Wt_data[31]\, 
        next_r0_0_cry_0_Y, \R1_data[0]\, \R1_data[1]\, 
        \R1_data[2]\, \R1_data[3]\, \R1_data[4]\, \R1_data[5]\, 
        \R1_data[6]\, \R1_data[7]\, \R1_data[8]\, \R1_data[9]\, 
        \R1_data[10]\, \R1_data[11]\, \R1_data[12]\, 
        \R1_data[13]\, \R1_data[14]\, \R1_data[15]\, 
        \R1_data[16]\, \R1_data[17]\, \R1_data[18]\, 
        \R1_data[19]\, \R1_data[20]\, \R1_data[21]\, 
        \R1_data[22]\, \R1_data[23]\, \R1_data[24]\, 
        \R1_data[25]\, \R1_data[26]\, \R1_data[27]\, 
        \R1_data[28]\, \R1_data[29]\, \R1_data[30]\, 
        \R1_data[31]\, \R2_data[0]\, \R2_data[1]\, \R2_data[2]\, 
        \R2_data[3]\, \R2_data[4]\, \R2_data[5]\, \R2_data[6]\, 
        \R2_data[7]\, \R2_data[8]\, \R2_data[9]\, \R2_data[10]\, 
        \R2_data[11]\, \R2_data[12]\, \R2_data[13]\, 
        \R2_data[14]\, \R2_data[15]\, \R2_data[16]\, 
        \R2_data[17]\, \R2_data[18]\, \R2_data[19]\, 
        \R2_data[20]\, \R2_data[21]\, \R2_data[22]\, 
        \R2_data[23]\, \R2_data[24]\, \R2_data[25]\, 
        \R2_data[26]\, \R2_data[27]\, \R2_data[28]\, 
        \R2_data[29]\, \R2_data[30]\, \R2_data[31]\, \R3_data[0]\, 
        \R3_data[1]\, \R3_data[2]\, \R3_data[3]\, \R3_data[4]\, 
        \R3_data[5]\, \R3_data[6]\, \R3_data[7]\, \R3_data[8]\, 
        \R3_data[9]\, \R3_data[10]\, \R3_data[11]\, \R3_data[12]\, 
        \R3_data[13]\, \R3_data[14]\, \R3_data[15]\, 
        \R3_data[16]\, \R3_data[17]\, \R3_data[18]\, 
        \R3_data[19]\, \R3_data[20]\, \R3_data[21]\, 
        \R3_data[22]\, \R3_data[23]\, \R3_data[24]\, 
        \R3_data[25]\, \R3_data[26]\, \R3_data[27]\, 
        \R3_data[28]\, \R3_data[29]\, \R3_data[30]\, 
        \R3_data[31]\, \R5_data[0]\, \R5_data[1]\, \R5_data[2]\, 
        \R5_data[3]\, \R5_data[4]\, \R5_data[5]\, \R5_data[6]\, 
        \R5_data[7]\, \R5_data[8]\, \R5_data[9]\, \R5_data[10]\, 
        \R5_data[11]\, \R5_data[12]\, \R5_data[13]\, 
        \R5_data[14]\, \R5_data[15]\, \R5_data[16]\, 
        \R5_data[17]\, \R5_data[18]\, \R5_data[19]\, 
        \R5_data[20]\, \R5_data[21]\, \R5_data[22]\, 
        \R5_data[23]\, \R5_data[24]\, \R5_data[25]\, 
        \R5_data[26]\, \R5_data[27]\, \R5_data[28]\, 
        \R5_data[29]\, \R5_data[30]\, \R5_data[31]\, \R6_data[0]\, 
        \R6_data[1]\, \R6_data[2]\, \R6_data[3]\, \R6_data[4]\, 
        \R6_data[5]\, \R6_data[6]\, \R6_data[7]\, \R6_data[8]\, 
        \R6_data[9]\, \R6_data[10]\, \R6_data[11]\, \R6_data[12]\, 
        \R6_data[13]\, \R6_data[14]\, \R6_data[15]\, 
        \R6_data[16]\, \R6_data[17]\, \R6_data[18]\, 
        \R6_data[19]\, \R6_data[20]\, \R6_data[21]\, 
        \R6_data[22]\, \R6_data[23]\, \R6_data[24]\, 
        \R6_data[25]\, \R6_data[26]\, \R6_data[27]\, 
        \R6_data[28]\, \R6_data[29]\, \R6_data[30]\, 
        \R6_data[31]\, \R7_data[0]\, \R7_data[1]\, \R7_data[2]\, 
        \R7_data[3]\, \R7_data[4]\, \R7_data[5]\, \R7_data[6]\, 
        \R7_data[7]\, \R7_data[8]\, \R7_data[9]\, \R7_data[10]\, 
        \R7_data[11]\, \R7_data[12]\, \R7_data[13]\, 
        \R7_data[14]\, \R7_data[15]\, \R7_data[16]\, 
        \R7_data[17]\, \R7_data[18]\, \R7_data[19]\, 
        \R7_data[20]\, \R7_data[21]\, \R7_data[22]\, 
        \R7_data[23]\, \R7_data[24]\, \R7_data[25]\, 
        \R7_data[26]\, \R7_data[27]\, \R7_data[28]\, 
        \R7_data[29]\, \R7_data[30]\, \R7_data[31]\, \R0_data[0]\, 
        \R0_data[1]\, \R0_data[2]\, \R0_data[3]\, \R0_data[4]\, 
        \R0_data[5]\, \R0_data[6]\, \R0_data[7]\, \R0_data[8]\, 
        \R0_data[9]\, \R0_data[10]\, \R0_data[11]\, \R0_data[12]\, 
        \R0_data[13]\, \R0_data[14]\, \R0_data[15]\, 
        \R0_data[16]\, \R0_data[17]\, \R0_data[18]\, 
        \R0_data[19]\, \R0_data[20]\, \R0_data[21]\, 
        \R0_data[22]\, \R0_data[23]\, \R0_data[24]\, 
        \R0_data[25]\, \R0_data[26]\, \R0_data[27]\, 
        \R0_data[28]\, \R0_data[29]\, \R0_data[30]\, 
        \R0_data[31]\, \R4_data[0]\, \R4_data[1]\, \R4_data[2]\, 
        \R4_data[3]\, \R4_data[4]\, \R4_data[5]\, \R4_data[6]\, 
        \R4_data[7]\, \R4_data[8]\, \R4_data[9]\, \R4_data[10]\, 
        \R4_data[11]\, \R4_data[12]\, \R4_data[13]\, 
        \R4_data[14]\, \R4_data[15]\, \R4_data[16]\, 
        \R4_data[17]\, \R4_data[18]\, \R4_data[19]\, 
        \R4_data[20]\, \R4_data[21]\, \R4_data[22]\, 
        \R4_data[23]\, \R4_data[24]\, \R4_data[25]\, 
        \R4_data[26]\, \R4_data[27]\, \R4_data[28]\, 
        \R4_data[29]\, \R4_data[30]\, \R4_data[31]\, \N4_data[1]\, 
        \N4_data[2]\, \N4_data[3]\, \N4_data[4]\, \N4_data[5]\, 
        \N4_data[6]\, \N4_data[7]\, \N4_data[8]\, \N4_data[9]\, 
        \N4_data[10]\, \N4_data[11]\, \N4_data[12]\, 
        \N4_data[13]\, \N4_data[14]\, \N4_data[15]\, 
        \N4_data[16]\, \N4_data[17]\, \N4_data[18]\, 
        \N4_data[19]\, \N4_data[20]\, \N4_data[21]\, 
        \N4_data[22]\, \N4_data[23]\, \N4_data[24]\, 
        \N4_data[25]\, \N4_data[26]\, \N4_data[27]\, 
        \N4_data[28]\, \N4_data[29]\, \N4_data[30]\, 
        \N4_data[31]\, \N0_data[1]\, \N0_data[2]\, \N0_data[3]\, 
        \N0_data[4]\, \N0_data[5]\, \N0_data[6]\, \N0_data[7]\, 
        \N0_data[8]\, \N0_data[9]\, \N0_data[10]\, \N0_data[11]\, 
        \N0_data[12]\, \N0_data[13]\, \N0_data[14]\, 
        \N0_data[15]\, \N0_data[16]\, \N0_data[17]\, 
        \N0_data[18]\, \N0_data[19]\, \N0_data[20]\, 
        \N0_data[21]\, \N0_data[22]\, \N0_data[23]\, 
        \N0_data[24]\, \N0_data[25]\, \N0_data[26]\, 
        \N0_data[27]\, \N0_data[28]\, \N0_data[29]\, 
        \N0_data[30]\, \N0_data[31]\, \N3_data[1]\, \N3_data[2]\, 
        \N3_data[3]\, \N3_data[4]\, \N3_data[5]\, \N3_data[6]\, 
        \N3_data[7]\, \N3_data[8]\, \N3_data[9]\, \N3_data[10]\, 
        \N3_data[11]\, \N3_data[12]\, \N3_data[13]\, 
        \N3_data[14]\, \N3_data[15]\, \N3_data[16]\, 
        \N3_data[17]\, \N3_data[18]\, \N3_data[19]\, 
        \N3_data[20]\, \N3_data[21]\, \N3_data[22]\, 
        \N3_data[23]\, \N3_data[24]\, \N3_data[25]\, 
        \N3_data[26]\, \N3_data[27]\, \N3_data[28]\, 
        \N3_data[29]\, \N3_data[30]\, \N3_data[31]\, \N2_data[1]\, 
        \N2_data[2]\, \N2_data[3]\, \N2_data[4]\, \N2_data[5]\, 
        \N2_data[6]\, \N2_data[7]\, \N2_data[8]\, \N2_data[9]\, 
        \N2_data[10]\, \N2_data[11]\, \N2_data[12]\, 
        \N2_data[13]\, \N2_data[14]\, \N2_data[15]\, 
        \N2_data[16]\, \N2_data[17]\, \N2_data[18]\, 
        \N2_data[19]\, \N2_data[20]\, \N2_data[21]\, 
        \N2_data[22]\, \N2_data[23]\, \N2_data[24]\, 
        \N2_data[25]\, \N2_data[26]\, \N2_data[27]\, 
        \N2_data[28]\, \N2_data[29]\, \N2_data[30]\, 
        \N2_data[31]\, \N1_data[1]\, \N1_data[2]\, \N1_data[3]\, 
        \N1_data[4]\, \N1_data[5]\, \N1_data[6]\, \N1_data[7]\, 
        \N1_data[8]\, \N1_data[9]\, \N1_data[10]\, \N1_data[11]\, 
        \N1_data[12]\, \N1_data[13]\, \N1_data[14]\, 
        \N1_data[15]\, \N1_data[16]\, \N1_data[17]\, 
        \N1_data[18]\, \N1_data[19]\, \N1_data[20]\, 
        \N1_data[21]\, \N1_data[22]\, \N1_data[23]\, 
        \N1_data[24]\, \N1_data[25]\, \N1_data[26]\, 
        \N1_data[27]\, \N1_data[28]\, \N1_data[29]\, 
        \N1_data[30]\, \N1_data[31]\, \N7_data[1]\, \N7_data[2]\, 
        \N7_data[3]\, \N7_data[4]\, \N7_data[5]\, \N7_data[6]\, 
        \N7_data[7]\, \N7_data[8]\, \N7_data[9]\, \N7_data[10]\, 
        \N7_data[11]\, \N7_data[12]\, \N7_data[13]\, 
        \N7_data[14]\, \N7_data[15]\, \N7_data[16]\, 
        \N7_data[17]\, \N7_data[18]\, \N7_data[19]\, 
        \N7_data[20]\, \N7_data[21]\, \N7_data[22]\, 
        \N7_data[23]\, \N7_data[24]\, \N7_data[25]\, 
        \N7_data[26]\, \N7_data[27]\, \N7_data[28]\, 
        \N7_data[29]\, \N7_data[30]\, \N7_data[31]\, \N6_data[1]\, 
        \N6_data[2]\, \N6_data[3]\, \N6_data[4]\, \N6_data[5]\, 
        \N6_data[6]\, \N6_data[7]\, \N6_data[8]\, \N6_data[9]\, 
        \N6_data[10]\, \N6_data[11]\, \N6_data[12]\, 
        \N6_data[13]\, \N6_data[14]\, \N6_data[15]\, 
        \N6_data[16]\, \N6_data[17]\, \N6_data[18]\, 
        \N6_data[19]\, \N6_data[20]\, \N6_data[21]\, 
        \N6_data[22]\, \N6_data[23]\, \N6_data[24]\, 
        \N6_data[25]\, \N6_data[26]\, \N6_data[27]\, 
        \N6_data[28]\, \N6_data[29]\, \N6_data[30]\, 
        \N6_data[31]\, \N5_data[1]\, \N5_data[2]\, \N5_data[3]\, 
        \N5_data[4]\, \N5_data[5]\, \N5_data[6]\, \N5_data[7]\, 
        \N5_data[8]\, \N5_data[9]\, \N5_data[10]\, \N5_data[11]\, 
        \N5_data[12]\, \N5_data[13]\, \N5_data[14]\, 
        \N5_data[15]\, \N5_data[16]\, \N5_data[17]\, 
        \N5_data[18]\, \N5_data[19]\, \N5_data[20]\, 
        \N5_data[21]\, \N5_data[22]\, \N5_data[23]\, 
        \N5_data[24]\, \N5_data[25]\, \N5_data[26]\, 
        \N5_data[27]\, \N5_data[28]\, \N5_data[29]\, 
        \N5_data[30]\, \N5_data[31]\, \Kt_data[15]\, 
        \Kt_data[24]\, \Kt_data[0]\, next_reg_H4_cry_0_0_Y, 
        next_reg_H0_cry_0_0_Y, m10_bm, m20_1, m10_am, m34, m49_am, 
        m49_bm, m62_am, m62_bm, m67_ns, m73, m78, m83_ns, m95_1_0, 
        m95_1_1, m104_am, m104_bm, m110_ns, m114, m119_ns, m124, 
        m137_am, m137_bm, m141, m144_ns, m157, m168_1_0, m168_1_1, 
        m172_ns, m177, m197_1_0, m197_1_1, m207_1_0, m207_1_1, 
        m215_am, m215_bm, m219, m222_ns, m226_ns, m230, m235_ns, 
        m239, m250_am, m250_bm, m254, m258_ns, m273, m276_ns, 
        m281_ns, m285, m289, m292_ns, m296, m300_ns, m304, 
        i3_mux_1, m325, m316, next_reg_H3_cry_0_0_Y, 
        next_reg_H2_cry_0_0_Y, next_reg_H1_cry_0_0_Y, 
        next_reg_H7_cry_0_0_Y, next_reg_H6_cry_0_0_Y, 
        next_reg_H5_cry_0_0_Y, GND_net_1, VCC_net_1 : std_logic;

    for all : sha256_control
	Use entity work.sha256_control(DEF_ARCH);
    for all : sha256_hash_core
	Use entity work.sha256_hash_core(DEF_ARCH);
    for all : sha256_regs
	Use entity work.sha256_regs(DEF_ARCH);
    for all : sha256_padding
	Use entity work.sha256_padding(DEF_ARCH);
    for all : sha256_msg_sch
	Use entity work.sha256_msg_sch(DEF_ARCH);
    for all : sha256_kt_rom
	Use entity work.sha256_kt_rom(DEF_ARCH);
begin 

    SHA256_Module_0_di_req_o <= \SHA256_Module_0_di_req_o\;

    Inst_sha256_control : sha256_control
      port map(hash_control_st_reg_i(6) => 
        \hash_control_st_reg_i[6]\, msg_bitlen(63) => 
        \msg_bitlen[63]\, msg_bitlen(62) => \msg_bitlen[62]\, 
        msg_bitlen(61) => \msg_bitlen[61]\, msg_bitlen(60) => 
        \msg_bitlen[60]\, msg_bitlen(59) => \msg_bitlen[59]\, 
        msg_bitlen(58) => \msg_bitlen[58]\, msg_bitlen(57) => 
        \msg_bitlen[57]\, msg_bitlen(56) => \msg_bitlen[56]\, 
        msg_bitlen(55) => \msg_bitlen[55]\, msg_bitlen(54) => 
        \msg_bitlen[54]\, msg_bitlen(53) => \msg_bitlen[53]\, 
        msg_bitlen(52) => \msg_bitlen[52]\, msg_bitlen(51) => 
        \msg_bitlen[51]\, msg_bitlen(50) => \msg_bitlen[50]\, 
        msg_bitlen(49) => \msg_bitlen[49]\, msg_bitlen(48) => 
        \msg_bitlen[48]\, msg_bitlen(47) => \msg_bitlen[47]\, 
        msg_bitlen(46) => \msg_bitlen[46]\, msg_bitlen(45) => 
        \msg_bitlen[45]\, msg_bitlen(44) => \msg_bitlen[44]\, 
        msg_bitlen(43) => \msg_bitlen[43]\, msg_bitlen(42) => 
        \msg_bitlen[42]\, msg_bitlen(41) => \msg_bitlen[41]\, 
        msg_bitlen(40) => \msg_bitlen[40]\, msg_bitlen(39) => 
        \msg_bitlen[39]\, msg_bitlen(38) => \msg_bitlen[38]\, 
        msg_bitlen(37) => \msg_bitlen[37]\, msg_bitlen(36) => 
        \msg_bitlen[36]\, msg_bitlen(35) => \msg_bitlen[35]\, 
        msg_bitlen(34) => \msg_bitlen[34]\, msg_bitlen(33) => 
        \msg_bitlen[33]\, msg_bitlen(32) => \msg_bitlen[32]\, 
        msg_bitlen(31) => \msg_bitlen[31]\, msg_bitlen(30) => 
        \msg_bitlen[30]\, msg_bitlen(29) => \msg_bitlen[29]\, 
        msg_bitlen(28) => \msg_bitlen[28]\, msg_bitlen(27) => 
        \msg_bitlen[27]\, msg_bitlen(26) => \msg_bitlen[26]\, 
        msg_bitlen(25) => \msg_bitlen[25]\, msg_bitlen(24) => 
        \msg_bitlen[24]\, msg_bitlen(23) => \msg_bitlen[23]\, 
        msg_bitlen(22) => \msg_bitlen[22]\, msg_bitlen(21) => 
        \msg_bitlen[21]\, msg_bitlen(20) => \msg_bitlen[20]\, 
        msg_bitlen(19) => \msg_bitlen[19]\, msg_bitlen(18) => 
        \msg_bitlen[18]\, msg_bitlen(17) => \msg_bitlen[17]\, 
        msg_bitlen(16) => \msg_bitlen[16]\, msg_bitlen(15) => 
        \msg_bitlen[15]\, msg_bitlen(14) => \msg_bitlen[14]\, 
        msg_bitlen(13) => \msg_bitlen[13]\, msg_bitlen(12) => 
        \msg_bitlen[12]\, msg_bitlen(11) => \msg_bitlen[11]\, 
        msg_bitlen(10) => \msg_bitlen[10]\, msg_bitlen(9) => 
        \msg_bitlen[9]\, msg_bitlen(8) => \msg_bitlen[8]\, 
        msg_bitlen(7) => \msg_bitlen[7]\, msg_bitlen(6) => 
        \msg_bitlen[6]\, msg_bitlen(5) => \msg_bitlen[5]\, 
        msg_bitlen(4) => \msg_bitlen[4]\, msg_bitlen(3) => 
        \msg_bitlen[3]\, Kt_addr(5) => \Kt_addr[5]\, Kt_addr(4)
         => \Kt_addr[4]\, Kt_addr(3) => \Kt_addr[3]\, Kt_addr(2)
         => \Kt_addr[2]\, Kt_addr(1) => \Kt_addr[1]\, Kt_addr(0)
         => \Kt_addr[0]\, st_cnt_reg(6) => \st_cnt_reg[6]\, 
        Kt_addr_fast(5) => \Kt_addr_fast[5]\, Kt_addr_fast(4) => 
        \Kt_addr_fast[4]\, Kt_addr_fast(3) => \Kt_addr_fast[3]\, 
        Kt_addr_fast(2) => \Kt_addr_fast[2]\, Kt_addr_fast(1) => 
        \Kt_addr_fast[1]\, Kt_addr_fast(0) => \Kt_addr_fast[0]\, 
        sha256_controller_0_bytes_o(1) => 
        sha256_controller_0_bytes_o(1), 
        hash_control_st_reg_ns_i_0_a2_0(4) => 
        \hash_control_st_reg_ns_i_0_a2_0[4]\, 
        hash_control_st_reg_ns_i_0_a2_2(4) => 
        \hash_control_st_reg_ns_i_0_a2_2[4]\, 
        hash_control_st_reg_2 => \hash_control_st_reg[2]\, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, one_insert => one_insert, 
        sha_last_blk_reg => sha_last_blk_reg, 
        SHA256_Module_0_di_req_o => \SHA256_Module_0_di_req_o\, 
        SHA256_Module_0_do_valid_o => SHA256_Module_0_do_valid_o, 
        Kt_addr_2_rep1 => Kt_addr_2_rep1, Kt_addr_2_rep2 => 
        Kt_addr_2_rep2, Kt_addr_1_rep1 => Kt_addr_1_rep1, 
        Kt_addr_1_rep2 => Kt_addr_1_rep2, Kt_addr_3_rep1 => 
        Kt_addr_3_rep1, Kt_addr_3_rep2 => Kt_addr_3_rep2, 
        Kt_addr_5_rep1 => Kt_addr_5_rep1, Kt_addr_0_rep1 => 
        Kt_addr_0_rep1, Kt_addr_0_rep2 => Kt_addr_0_rep2, 
        Kt_addr_4_rep1 => Kt_addr_4_rep1, Kt_addr_4_rep2 => 
        Kt_addr_4_rep2, sha256_controller_0_end_o => 
        sha256_controller_0_end_o, last_block_0 => last_block_0, 
        N_168_i_0 => N_168_i_0, ce_i_i_2 => ce_i_i_2, 
        pad_one_reg_0_0_a2_0 => pad_one_reg_0_0_a2_0, 
        sha_last_blk_next_0_o2_0 => sha_last_blk_next_0_o2_0, 
        oregs_ce_i_a2_0_a2 => oregs_ce_i_a2_0_a2, N_102 => N_102, 
        N_28 => N_28, N_387 => N_387, N_388 => N_388, W_m4_e_2
         => W_m4_e_2, N_105 => N_105, N_111 => N_111, 
        core_ce_o_iv_i_0 => core_ce_o_iv_i_0, N_244_i_0 => 
        N_244_i_0, SHA256_Module_0_error_o => 
        SHA256_Module_0_error_o, ld_i_i_3 => ld_i_i_3);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    Inst_sha256_hash_core : sha256_hash_core
      port map(R1_data(31) => \R1_data[31]\, R1_data(30) => 
        \R1_data[30]\, R1_data(29) => \R1_data[29]\, R1_data(28)
         => \R1_data[28]\, R1_data(27) => \R1_data[27]\, 
        R1_data(26) => \R1_data[26]\, R1_data(25) => 
        \R1_data[25]\, R1_data(24) => \R1_data[24]\, R1_data(23)
         => \R1_data[23]\, R1_data(22) => \R1_data[22]\, 
        R1_data(21) => \R1_data[21]\, R1_data(20) => 
        \R1_data[20]\, R1_data(19) => \R1_data[19]\, R1_data(18)
         => \R1_data[18]\, R1_data(17) => \R1_data[17]\, 
        R1_data(16) => \R1_data[16]\, R1_data(15) => 
        \R1_data[15]\, R1_data(14) => \R1_data[14]\, R1_data(13)
         => \R1_data[13]\, R1_data(12) => \R1_data[12]\, 
        R1_data(11) => \R1_data[11]\, R1_data(10) => 
        \R1_data[10]\, R1_data(9) => \R1_data[9]\, R1_data(8) => 
        \R1_data[8]\, R1_data(7) => \R1_data[7]\, R1_data(6) => 
        \R1_data[6]\, R1_data(5) => \R1_data[5]\, R1_data(4) => 
        \R1_data[4]\, R1_data(3) => \R1_data[3]\, R1_data(2) => 
        \R1_data[2]\, R1_data(1) => \R1_data[1]\, R1_data(0) => 
        \R1_data[0]\, R2_data(31) => \R2_data[31]\, R2_data(30)
         => \R2_data[30]\, R2_data(29) => \R2_data[29]\, 
        R2_data(28) => \R2_data[28]\, R2_data(27) => 
        \R2_data[27]\, R2_data(26) => \R2_data[26]\, R2_data(25)
         => \R2_data[25]\, R2_data(24) => \R2_data[24]\, 
        R2_data(23) => \R2_data[23]\, R2_data(22) => 
        \R2_data[22]\, R2_data(21) => \R2_data[21]\, R2_data(20)
         => \R2_data[20]\, R2_data(19) => \R2_data[19]\, 
        R2_data(18) => \R2_data[18]\, R2_data(17) => 
        \R2_data[17]\, R2_data(16) => \R2_data[16]\, R2_data(15)
         => \R2_data[15]\, R2_data(14) => \R2_data[14]\, 
        R2_data(13) => \R2_data[13]\, R2_data(12) => 
        \R2_data[12]\, R2_data(11) => \R2_data[11]\, R2_data(10)
         => \R2_data[10]\, R2_data(9) => \R2_data[9]\, R2_data(8)
         => \R2_data[8]\, R2_data(7) => \R2_data[7]\, R2_data(6)
         => \R2_data[6]\, R2_data(5) => \R2_data[5]\, R2_data(4)
         => \R2_data[4]\, R2_data(3) => \R2_data[3]\, R2_data(2)
         => \R2_data[2]\, R2_data(1) => \R2_data[1]\, R2_data(0)
         => \R2_data[0]\, R3_data(31) => \R3_data[31]\, 
        R3_data(30) => \R3_data[30]\, R3_data(29) => 
        \R3_data[29]\, R3_data(28) => \R3_data[28]\, R3_data(27)
         => \R3_data[27]\, R3_data(26) => \R3_data[26]\, 
        R3_data(25) => \R3_data[25]\, R3_data(24) => 
        \R3_data[24]\, R3_data(23) => \R3_data[23]\, R3_data(22)
         => \R3_data[22]\, R3_data(21) => \R3_data[21]\, 
        R3_data(20) => \R3_data[20]\, R3_data(19) => 
        \R3_data[19]\, R3_data(18) => \R3_data[18]\, R3_data(17)
         => \R3_data[17]\, R3_data(16) => \R3_data[16]\, 
        R3_data(15) => \R3_data[15]\, R3_data(14) => 
        \R3_data[14]\, R3_data(13) => \R3_data[13]\, R3_data(12)
         => \R3_data[12]\, R3_data(11) => \R3_data[11]\, 
        R3_data(10) => \R3_data[10]\, R3_data(9) => \R3_data[9]\, 
        R3_data(8) => \R3_data[8]\, R3_data(7) => \R3_data[7]\, 
        R3_data(6) => \R3_data[6]\, R3_data(5) => \R3_data[5]\, 
        R3_data(4) => \R3_data[4]\, R3_data(3) => \R3_data[3]\, 
        R3_data(2) => \R3_data[2]\, R3_data(1) => \R3_data[1]\, 
        R3_data(0) => \R3_data[0]\, R5_data(31) => \R5_data[31]\, 
        R5_data(30) => \R5_data[30]\, R5_data(29) => 
        \R5_data[29]\, R5_data(28) => \R5_data[28]\, R5_data(27)
         => \R5_data[27]\, R5_data(26) => \R5_data[26]\, 
        R5_data(25) => \R5_data[25]\, R5_data(24) => 
        \R5_data[24]\, R5_data(23) => \R5_data[23]\, R5_data(22)
         => \R5_data[22]\, R5_data(21) => \R5_data[21]\, 
        R5_data(20) => \R5_data[20]\, R5_data(19) => 
        \R5_data[19]\, R5_data(18) => \R5_data[18]\, R5_data(17)
         => \R5_data[17]\, R5_data(16) => \R5_data[16]\, 
        R5_data(15) => \R5_data[15]\, R5_data(14) => 
        \R5_data[14]\, R5_data(13) => \R5_data[13]\, R5_data(12)
         => \R5_data[12]\, R5_data(11) => \R5_data[11]\, 
        R5_data(10) => \R5_data[10]\, R5_data(9) => \R5_data[9]\, 
        R5_data(8) => \R5_data[8]\, R5_data(7) => \R5_data[7]\, 
        R5_data(6) => \R5_data[6]\, R5_data(5) => \R5_data[5]\, 
        R5_data(4) => \R5_data[4]\, R5_data(3) => \R5_data[3]\, 
        R5_data(2) => \R5_data[2]\, R5_data(1) => \R5_data[1]\, 
        R5_data(0) => \R5_data[0]\, R6_data(31) => \R6_data[31]\, 
        R6_data(30) => \R6_data[30]\, R6_data(29) => 
        \R6_data[29]\, R6_data(28) => \R6_data[28]\, R6_data(27)
         => \R6_data[27]\, R6_data(26) => \R6_data[26]\, 
        R6_data(25) => \R6_data[25]\, R6_data(24) => 
        \R6_data[24]\, R6_data(23) => \R6_data[23]\, R6_data(22)
         => \R6_data[22]\, R6_data(21) => \R6_data[21]\, 
        R6_data(20) => \R6_data[20]\, R6_data(19) => 
        \R6_data[19]\, R6_data(18) => \R6_data[18]\, R6_data(17)
         => \R6_data[17]\, R6_data(16) => \R6_data[16]\, 
        R6_data(15) => \R6_data[15]\, R6_data(14) => 
        \R6_data[14]\, R6_data(13) => \R6_data[13]\, R6_data(12)
         => \R6_data[12]\, R6_data(11) => \R6_data[11]\, 
        R6_data(10) => \R6_data[10]\, R6_data(9) => \R6_data[9]\, 
        R6_data(8) => \R6_data[8]\, R6_data(7) => \R6_data[7]\, 
        R6_data(6) => \R6_data[6]\, R6_data(5) => \R6_data[5]\, 
        R6_data(4) => \R6_data[4]\, R6_data(3) => \R6_data[3]\, 
        R6_data(2) => \R6_data[2]\, R6_data(1) => \R6_data[1]\, 
        R6_data(0) => \R6_data[0]\, R7_data(31) => \R7_data[31]\, 
        R7_data(30) => \R7_data[30]\, R7_data(29) => 
        \R7_data[29]\, R7_data(28) => \R7_data[28]\, R7_data(27)
         => \R7_data[27]\, R7_data(26) => \R7_data[26]\, 
        R7_data(25) => \R7_data[25]\, R7_data(24) => 
        \R7_data[24]\, R7_data(23) => \R7_data[23]\, R7_data(22)
         => \R7_data[22]\, R7_data(21) => \R7_data[21]\, 
        R7_data(20) => \R7_data[20]\, R7_data(19) => 
        \R7_data[19]\, R7_data(18) => \R7_data[18]\, R7_data(17)
         => \R7_data[17]\, R7_data(16) => \R7_data[16]\, 
        R7_data(15) => \R7_data[15]\, R7_data(14) => 
        \R7_data[14]\, R7_data(13) => \R7_data[13]\, R7_data(12)
         => \R7_data[12]\, R7_data(11) => \R7_data[11]\, 
        R7_data(10) => \R7_data[10]\, R7_data(9) => \R7_data[9]\, 
        R7_data(8) => \R7_data[8]\, R7_data(7) => \R7_data[7]\, 
        R7_data(6) => \R7_data[6]\, R7_data(5) => \R7_data[5]\, 
        R7_data(4) => \R7_data[4]\, R7_data(3) => \R7_data[3]\, 
        R7_data(2) => \R7_data[2]\, R7_data(1) => \R7_data[1]\, 
        R7_data(0) => \R7_data[0]\, R0_data(31) => \R0_data[31]\, 
        R0_data(30) => \R0_data[30]\, R0_data(29) => 
        \R0_data[29]\, R0_data(28) => \R0_data[28]\, R0_data(27)
         => \R0_data[27]\, R0_data(26) => \R0_data[26]\, 
        R0_data(25) => \R0_data[25]\, R0_data(24) => 
        \R0_data[24]\, R0_data(23) => \R0_data[23]\, R0_data(22)
         => \R0_data[22]\, R0_data(21) => \R0_data[21]\, 
        R0_data(20) => \R0_data[20]\, R0_data(19) => 
        \R0_data[19]\, R0_data(18) => \R0_data[18]\, R0_data(17)
         => \R0_data[17]\, R0_data(16) => \R0_data[16]\, 
        R0_data(15) => \R0_data[15]\, R0_data(14) => 
        \R0_data[14]\, R0_data(13) => \R0_data[13]\, R0_data(12)
         => \R0_data[12]\, R0_data(11) => \R0_data[11]\, 
        R0_data(10) => \R0_data[10]\, R0_data(9) => \R0_data[9]\, 
        R0_data(8) => \R0_data[8]\, R0_data(7) => \R0_data[7]\, 
        R0_data(6) => \R0_data[6]\, R0_data(5) => \R0_data[5]\, 
        R0_data(4) => \R0_data[4]\, R0_data(3) => \R0_data[3]\, 
        R0_data(2) => \R0_data[2]\, R0_data(1) => \R0_data[1]\, 
        R0_data(0) => \R0_data[0]\, R4_data(31) => \R4_data[31]\, 
        R4_data(30) => \R4_data[30]\, R4_data(29) => 
        \R4_data[29]\, R4_data(28) => \R4_data[28]\, R4_data(27)
         => \R4_data[27]\, R4_data(26) => \R4_data[26]\, 
        R4_data(25) => \R4_data[25]\, R4_data(24) => 
        \R4_data[24]\, R4_data(23) => \R4_data[23]\, R4_data(22)
         => \R4_data[22]\, R4_data(21) => \R4_data[21]\, 
        R4_data(20) => \R4_data[20]\, R4_data(19) => 
        \R4_data[19]\, R4_data(18) => \R4_data[18]\, R4_data(17)
         => \R4_data[17]\, R4_data(16) => \R4_data[16]\, 
        R4_data(15) => \R4_data[15]\, R4_data(14) => 
        \R4_data[14]\, R4_data(13) => \R4_data[13]\, R4_data(12)
         => \R4_data[12]\, R4_data(11) => \R4_data[11]\, 
        R4_data(10) => \R4_data[10]\, R4_data(9) => \R4_data[9]\, 
        R4_data(8) => \R4_data[8]\, R4_data(7) => \R4_data[7]\, 
        R4_data(6) => \R4_data[6]\, R4_data(5) => \R4_data[5]\, 
        R4_data(4) => \R4_data[4]\, R4_data(3) => \R4_data[3]\, 
        R4_data(2) => \R4_data[2]\, R4_data(1) => \R4_data[1]\, 
        R4_data(0) => \R4_data[0]\, N4_data(31) => \N4_data[31]\, 
        N4_data(30) => \N4_data[30]\, N4_data(29) => 
        \N4_data[29]\, N4_data(28) => \N4_data[28]\, N4_data(27)
         => \N4_data[27]\, N4_data(26) => \N4_data[26]\, 
        N4_data(25) => \N4_data[25]\, N4_data(24) => 
        \N4_data[24]\, N4_data(23) => \N4_data[23]\, N4_data(22)
         => \N4_data[22]\, N4_data(21) => \N4_data[21]\, 
        N4_data(20) => \N4_data[20]\, N4_data(19) => 
        \N4_data[19]\, N4_data(18) => \N4_data[18]\, N4_data(17)
         => \N4_data[17]\, N4_data(16) => \N4_data[16]\, 
        N4_data(15) => \N4_data[15]\, N4_data(14) => 
        \N4_data[14]\, N4_data(13) => \N4_data[13]\, N4_data(12)
         => \N4_data[12]\, N4_data(11) => \N4_data[11]\, 
        N4_data(10) => \N4_data[10]\, N4_data(9) => \N4_data[9]\, 
        N4_data(8) => \N4_data[8]\, N4_data(7) => \N4_data[7]\, 
        N4_data(6) => \N4_data[6]\, N4_data(5) => \N4_data[5]\, 
        N4_data(4) => \N4_data[4]\, N4_data(3) => \N4_data[3]\, 
        N4_data(2) => \N4_data[2]\, N4_data(1) => \N4_data[1]\, 
        N0_data(31) => \N0_data[31]\, N0_data(30) => 
        \N0_data[30]\, N0_data(29) => \N0_data[29]\, N0_data(28)
         => \N0_data[28]\, N0_data(27) => \N0_data[27]\, 
        N0_data(26) => \N0_data[26]\, N0_data(25) => 
        \N0_data[25]\, N0_data(24) => \N0_data[24]\, N0_data(23)
         => \N0_data[23]\, N0_data(22) => \N0_data[22]\, 
        N0_data(21) => \N0_data[21]\, N0_data(20) => 
        \N0_data[20]\, N0_data(19) => \N0_data[19]\, N0_data(18)
         => \N0_data[18]\, N0_data(17) => \N0_data[17]\, 
        N0_data(16) => \N0_data[16]\, N0_data(15) => 
        \N0_data[15]\, N0_data(14) => \N0_data[14]\, N0_data(13)
         => \N0_data[13]\, N0_data(12) => \N0_data[12]\, 
        N0_data(11) => \N0_data[11]\, N0_data(10) => 
        \N0_data[10]\, N0_data(9) => \N0_data[9]\, N0_data(8) => 
        \N0_data[8]\, N0_data(7) => \N0_data[7]\, N0_data(6) => 
        \N0_data[6]\, N0_data(5) => \N0_data[5]\, N0_data(4) => 
        \N0_data[4]\, N0_data(3) => \N0_data[3]\, N0_data(2) => 
        \N0_data[2]\, N0_data(1) => \N0_data[1]\, W_out_i_0(0)
         => \W_out_i_0[0]\, Kt_addr(5) => \Kt_addr[5]\, 
        N3_data(31) => \N3_data[31]\, N3_data(30) => 
        \N3_data[30]\, N3_data(29) => \N3_data[29]\, N3_data(28)
         => \N3_data[28]\, N3_data(27) => \N3_data[27]\, 
        N3_data(26) => \N3_data[26]\, N3_data(25) => 
        \N3_data[25]\, N3_data(24) => \N3_data[24]\, N3_data(23)
         => \N3_data[23]\, N3_data(22) => \N3_data[22]\, 
        N3_data(21) => \N3_data[21]\, N3_data(20) => 
        \N3_data[20]\, N3_data(19) => \N3_data[19]\, N3_data(18)
         => \N3_data[18]\, N3_data(17) => \N3_data[17]\, 
        N3_data(16) => \N3_data[16]\, N3_data(15) => 
        \N3_data[15]\, N3_data(14) => \N3_data[14]\, N3_data(13)
         => \N3_data[13]\, N3_data(12) => \N3_data[12]\, 
        N3_data(11) => \N3_data[11]\, N3_data(10) => 
        \N3_data[10]\, N3_data(9) => \N3_data[9]\, N3_data(8) => 
        \N3_data[8]\, N3_data(7) => \N3_data[7]\, N3_data(6) => 
        \N3_data[6]\, N3_data(5) => \N3_data[5]\, N3_data(4) => 
        \N3_data[4]\, N3_data(3) => \N3_data[3]\, N3_data(2) => 
        \N3_data[2]\, N3_data(1) => \N3_data[1]\, N2_data(31) => 
        \N2_data[31]\, N2_data(30) => \N2_data[30]\, N2_data(29)
         => \N2_data[29]\, N2_data(28) => \N2_data[28]\, 
        N2_data(27) => \N2_data[27]\, N2_data(26) => 
        \N2_data[26]\, N2_data(25) => \N2_data[25]\, N2_data(24)
         => \N2_data[24]\, N2_data(23) => \N2_data[23]\, 
        N2_data(22) => \N2_data[22]\, N2_data(21) => 
        \N2_data[21]\, N2_data(20) => \N2_data[20]\, N2_data(19)
         => \N2_data[19]\, N2_data(18) => \N2_data[18]\, 
        N2_data(17) => \N2_data[17]\, N2_data(16) => 
        \N2_data[16]\, N2_data(15) => \N2_data[15]\, N2_data(14)
         => \N2_data[14]\, N2_data(13) => \N2_data[13]\, 
        N2_data(12) => \N2_data[12]\, N2_data(11) => 
        \N2_data[11]\, N2_data(10) => \N2_data[10]\, N2_data(9)
         => \N2_data[9]\, N2_data(8) => \N2_data[8]\, N2_data(7)
         => \N2_data[7]\, N2_data(6) => \N2_data[6]\, N2_data(5)
         => \N2_data[5]\, N2_data(4) => \N2_data[4]\, N2_data(3)
         => \N2_data[3]\, N2_data(2) => \N2_data[2]\, N2_data(1)
         => \N2_data[1]\, N1_data(31) => \N1_data[31]\, 
        N1_data(30) => \N1_data[30]\, N1_data(29) => 
        \N1_data[29]\, N1_data(28) => \N1_data[28]\, N1_data(27)
         => \N1_data[27]\, N1_data(26) => \N1_data[26]\, 
        N1_data(25) => \N1_data[25]\, N1_data(24) => 
        \N1_data[24]\, N1_data(23) => \N1_data[23]\, N1_data(22)
         => \N1_data[22]\, N1_data(21) => \N1_data[21]\, 
        N1_data(20) => \N1_data[20]\, N1_data(19) => 
        \N1_data[19]\, N1_data(18) => \N1_data[18]\, N1_data(17)
         => \N1_data[17]\, N1_data(16) => \N1_data[16]\, 
        N1_data(15) => \N1_data[15]\, N1_data(14) => 
        \N1_data[14]\, N1_data(13) => \N1_data[13]\, N1_data(12)
         => \N1_data[12]\, N1_data(11) => \N1_data[11]\, 
        N1_data(10) => \N1_data[10]\, N1_data(9) => \N1_data[9]\, 
        N1_data(8) => \N1_data[8]\, N1_data(7) => \N1_data[7]\, 
        N1_data(6) => \N1_data[6]\, N1_data(5) => \N1_data[5]\, 
        N1_data(4) => \N1_data[4]\, N1_data(3) => \N1_data[3]\, 
        N1_data(2) => \N1_data[2]\, N1_data(1) => \N1_data[1]\, 
        N7_data(31) => \N7_data[31]\, N7_data(30) => 
        \N7_data[30]\, N7_data(29) => \N7_data[29]\, N7_data(28)
         => \N7_data[28]\, N7_data(27) => \N7_data[27]\, 
        N7_data(26) => \N7_data[26]\, N7_data(25) => 
        \N7_data[25]\, N7_data(24) => \N7_data[24]\, N7_data(23)
         => \N7_data[23]\, N7_data(22) => \N7_data[22]\, 
        N7_data(21) => \N7_data[21]\, N7_data(20) => 
        \N7_data[20]\, N7_data(19) => \N7_data[19]\, N7_data(18)
         => \N7_data[18]\, N7_data(17) => \N7_data[17]\, 
        N7_data(16) => \N7_data[16]\, N7_data(15) => 
        \N7_data[15]\, N7_data(14) => \N7_data[14]\, N7_data(13)
         => \N7_data[13]\, N7_data(12) => \N7_data[12]\, 
        N7_data(11) => \N7_data[11]\, N7_data(10) => 
        \N7_data[10]\, N7_data(9) => \N7_data[9]\, N7_data(8) => 
        \N7_data[8]\, N7_data(7) => \N7_data[7]\, N7_data(6) => 
        \N7_data[6]\, N7_data(5) => \N7_data[5]\, N7_data(4) => 
        \N7_data[4]\, N7_data(3) => \N7_data[3]\, N7_data(2) => 
        \N7_data[2]\, N7_data(1) => \N7_data[1]\, N6_data(31) => 
        \N6_data[31]\, N6_data(30) => \N6_data[30]\, N6_data(29)
         => \N6_data[29]\, N6_data(28) => \N6_data[28]\, 
        N6_data(27) => \N6_data[27]\, N6_data(26) => 
        \N6_data[26]\, N6_data(25) => \N6_data[25]\, N6_data(24)
         => \N6_data[24]\, N6_data(23) => \N6_data[23]\, 
        N6_data(22) => \N6_data[22]\, N6_data(21) => 
        \N6_data[21]\, N6_data(20) => \N6_data[20]\, N6_data(19)
         => \N6_data[19]\, N6_data(18) => \N6_data[18]\, 
        N6_data(17) => \N6_data[17]\, N6_data(16) => 
        \N6_data[16]\, N6_data(15) => \N6_data[15]\, N6_data(14)
         => \N6_data[14]\, N6_data(13) => \N6_data[13]\, 
        N6_data(12) => \N6_data[12]\, N6_data(11) => 
        \N6_data[11]\, N6_data(10) => \N6_data[10]\, N6_data(9)
         => \N6_data[9]\, N6_data(8) => \N6_data[8]\, N6_data(7)
         => \N6_data[7]\, N6_data(6) => \N6_data[6]\, N6_data(5)
         => \N6_data[5]\, N6_data(4) => \N6_data[4]\, N6_data(3)
         => \N6_data[3]\, N6_data(2) => \N6_data[2]\, N6_data(1)
         => \N6_data[1]\, N5_data(31) => \N5_data[31]\, 
        N5_data(30) => \N5_data[30]\, N5_data(29) => 
        \N5_data[29]\, N5_data(28) => \N5_data[28]\, N5_data(27)
         => \N5_data[27]\, N5_data(26) => \N5_data[26]\, 
        N5_data(25) => \N5_data[25]\, N5_data(24) => 
        \N5_data[24]\, N5_data(23) => \N5_data[23]\, N5_data(22)
         => \N5_data[22]\, N5_data(21) => \N5_data[21]\, 
        N5_data(20) => \N5_data[20]\, N5_data(19) => 
        \N5_data[19]\, N5_data(18) => \N5_data[18]\, N5_data(17)
         => \N5_data[17]\, N5_data(16) => \N5_data[16]\, 
        N5_data(15) => \N5_data[15]\, N5_data(14) => 
        \N5_data[14]\, N5_data(13) => \N5_data[13]\, N5_data(12)
         => \N5_data[12]\, N5_data(11) => \N5_data[11]\, 
        N5_data(10) => \N5_data[10]\, N5_data(9) => \N5_data[9]\, 
        N5_data(8) => \N5_data[8]\, N5_data(7) => \N5_data[7]\, 
        N5_data(6) => \N5_data[6]\, N5_data(5) => \N5_data[5]\, 
        N5_data(4) => \N5_data[4]\, N5_data(3) => \N5_data[3]\, 
        N5_data(2) => \N5_data[2]\, N5_data(1) => \N5_data[1]\, 
        Wt_data(31) => \Wt_data[31]\, Wt_data(30) => 
        \Wt_data[30]\, Wt_data(29) => \Wt_data[29]\, Wt_data(28)
         => \Wt_data[28]\, Wt_data(27) => \Wt_data[27]\, 
        Wt_data(26) => \Wt_data[26]\, Wt_data(25) => 
        \Wt_data[25]\, Wt_data(24) => \Wt_data[24]\, Wt_data(23)
         => \Wt_data[23]\, Wt_data(22) => \Wt_data[22]\, 
        Wt_data(21) => \Wt_data[21]\, Wt_data(20) => 
        \Wt_data[20]\, Wt_data(19) => \Wt_data[19]\, Wt_data(18)
         => \Wt_data[18]\, Wt_data(17) => \Wt_data[17]\, 
        Wt_data(16) => \Wt_data[16]\, Wt_data(15) => 
        \Wt_data[15]\, Wt_data(14) => \Wt_data[14]\, Wt_data(13)
         => \Wt_data[13]\, Wt_data(12) => \Wt_data[12]\, 
        Wt_data(11) => \Wt_data[11]\, Wt_data(10) => 
        \Wt_data[10]\, Wt_data(9) => \Wt_data[9]\, Wt_data(8) => 
        \Wt_data[8]\, Wt_data(7) => \Wt_data[7]\, Wt_data(6) => 
        \Wt_data[6]\, Wt_data(5) => \Wt_data[5]\, Wt_data(4) => 
        \Wt_data[4]\, Wt_data(3) => \Wt_data[3]\, Wt_data(2) => 
        \Wt_data[2]\, Wt_data(1) => \Wt_data[1]\, Wt_data(0) => 
        \Wt_data[0]\, Kt_data_15 => \Kt_data[15]\, Kt_data_24 => 
        \Kt_data[24]\, Kt_data_0 => \Kt_data[0]\, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, core_ce_o_iv_i_0 => 
        core_ce_o_iv_i_0, oregs_ce_i_a2_0_a2 => 
        oregs_ce_i_a2_0_a2, next_reg_H4_cry_0_0_Y => 
        next_reg_H4_cry_0_0_Y, next_reg_H0_cry_0_0_Y => 
        next_reg_H0_cry_0_0_Y, next_r0_0_cry_0_Y => 
        next_r0_0_cry_0_Y, ld_i_i_3 => ld_i_i_3, N_98 => N_98, 
        m10_bm => m10_bm, m20_1 => m20_1, m10_am => m10_am, m34
         => m34, m49_am => m49_am, m49_bm => m49_bm, 
        Kt_addr_5_rep1 => Kt_addr_5_rep1, m62_am => m62_am, 
        m62_bm => m62_bm, m67_ns => m67_ns, m73 => m73, m78 => 
        m78, m83_ns => m83_ns, m95_1_0 => m95_1_0, m95_1_1 => 
        m95_1_1, m104_am => m104_am, m104_bm => m104_bm, m110_ns
         => m110_ns, m114 => m114, m119_ns => m119_ns, m124 => 
        m124, m137_am => m137_am, m137_bm => m137_bm, m141 => 
        m141, m144_ns => m144_ns, m157 => m157, m168_1_0 => 
        m168_1_0, m168_1_1 => m168_1_1, m172_ns => m172_ns, m177
         => m177, m197_1_0 => m197_1_0, m197_1_1 => m197_1_1, 
        m207_1_0 => m207_1_0, m207_1_1 => m207_1_1, m215_am => 
        m215_am, m215_bm => m215_bm, m219 => m219, m222_ns => 
        m222_ns, m226_ns => m226_ns, m230 => m230, m235_ns => 
        m235_ns, m239 => m239, m250_am => m250_am, m250_bm => 
        m250_bm, m254 => m254, m258_ns => m258_ns, m273 => m273, 
        m276_ns => m276_ns, m281_ns => m281_ns, m285 => m285, 
        m289 => m289, m292_ns => m292_ns, m296 => m296, m300_ns
         => m300_ns, m304 => m304, i3_mux_1 => i3_mux_1, m325 => 
        m325, m316 => m316, next_reg_H3_cry_0_0_Y => 
        next_reg_H3_cry_0_0_Y, next_reg_H2_cry_0_0_Y => 
        next_reg_H2_cry_0_0_Y, next_reg_H1_cry_0_0_Y => 
        next_reg_H1_cry_0_0_Y, next_reg_H7_cry_0_0_Y => 
        next_reg_H7_cry_0_0_Y, next_reg_H6_cry_0_0_Y => 
        next_reg_H6_cry_0_0_Y, next_reg_H5_cry_0_0_Y => 
        next_reg_H5_cry_0_0_Y);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    Inst_sha256_regs : sha256_regs
      port map(SHA256_BLOCK_0_H0_o(31) => SHA256_BLOCK_0_H0_o(31), 
        SHA256_BLOCK_0_H0_o(30) => SHA256_BLOCK_0_H0_o(30), 
        SHA256_BLOCK_0_H0_o(29) => SHA256_BLOCK_0_H0_o(29), 
        SHA256_BLOCK_0_H0_o(28) => SHA256_BLOCK_0_H0_o(28), 
        SHA256_BLOCK_0_H0_o(27) => SHA256_BLOCK_0_H0_o(27), 
        SHA256_BLOCK_0_H0_o(26) => SHA256_BLOCK_0_H0_o(26), 
        SHA256_BLOCK_0_H0_o(25) => SHA256_BLOCK_0_H0_o(25), 
        SHA256_BLOCK_0_H0_o(24) => SHA256_BLOCK_0_H0_o(24), 
        SHA256_BLOCK_0_H0_o(23) => SHA256_BLOCK_0_H0_o(23), 
        SHA256_BLOCK_0_H0_o(22) => SHA256_BLOCK_0_H0_o(22), 
        SHA256_BLOCK_0_H0_o(21) => SHA256_BLOCK_0_H0_o(21), 
        SHA256_BLOCK_0_H0_o(20) => SHA256_BLOCK_0_H0_o(20), 
        SHA256_BLOCK_0_H0_o(19) => SHA256_BLOCK_0_H0_o(19), 
        SHA256_BLOCK_0_H0_o(18) => SHA256_BLOCK_0_H0_o(18), 
        SHA256_BLOCK_0_H0_o(17) => SHA256_BLOCK_0_H0_o(17), 
        SHA256_BLOCK_0_H0_o(16) => SHA256_BLOCK_0_H0_o(16), 
        SHA256_BLOCK_0_H0_o(15) => SHA256_BLOCK_0_H0_o(15), 
        SHA256_BLOCK_0_H0_o(14) => SHA256_BLOCK_0_H0_o(14), 
        SHA256_BLOCK_0_H0_o(13) => SHA256_BLOCK_0_H0_o(13), 
        SHA256_BLOCK_0_H0_o(12) => SHA256_BLOCK_0_H0_o(12), 
        SHA256_BLOCK_0_H0_o(11) => SHA256_BLOCK_0_H0_o(11), 
        SHA256_BLOCK_0_H0_o(10) => SHA256_BLOCK_0_H0_o(10), 
        SHA256_BLOCK_0_H0_o(9) => SHA256_BLOCK_0_H0_o(9), 
        SHA256_BLOCK_0_H0_o(8) => SHA256_BLOCK_0_H0_o(8), 
        SHA256_BLOCK_0_H0_o(7) => SHA256_BLOCK_0_H0_o(7), 
        SHA256_BLOCK_0_H0_o(6) => SHA256_BLOCK_0_H0_o(6), 
        SHA256_BLOCK_0_H0_o(5) => SHA256_BLOCK_0_H0_o(5), 
        SHA256_BLOCK_0_H0_o(4) => SHA256_BLOCK_0_H0_o(4), 
        SHA256_BLOCK_0_H0_o(3) => SHA256_BLOCK_0_H0_o(3), 
        SHA256_BLOCK_0_H0_o(2) => SHA256_BLOCK_0_H0_o(2), 
        SHA256_BLOCK_0_H0_o(1) => SHA256_BLOCK_0_H0_o(1), 
        SHA256_BLOCK_0_H0_o(0) => SHA256_BLOCK_0_H0_o(0), 
        N0_data(31) => \N0_data[31]\, N0_data(30) => 
        \N0_data[30]\, N0_data(29) => \N0_data[29]\, N0_data(28)
         => \N0_data[28]\, N0_data(27) => \N0_data[27]\, 
        N0_data(26) => \N0_data[26]\, N0_data(25) => 
        \N0_data[25]\, N0_data(24) => \N0_data[24]\, N0_data(23)
         => \N0_data[23]\, N0_data(22) => \N0_data[22]\, 
        N0_data(21) => \N0_data[21]\, N0_data(20) => 
        \N0_data[20]\, N0_data(19) => \N0_data[19]\, N0_data(18)
         => \N0_data[18]\, N0_data(17) => \N0_data[17]\, 
        N0_data(16) => \N0_data[16]\, N0_data(15) => 
        \N0_data[15]\, N0_data(14) => \N0_data[14]\, N0_data(13)
         => \N0_data[13]\, N0_data(12) => \N0_data[12]\, 
        N0_data(11) => \N0_data[11]\, N0_data(10) => 
        \N0_data[10]\, N0_data(9) => \N0_data[9]\, N0_data(8) => 
        \N0_data[8]\, N0_data(7) => \N0_data[7]\, N0_data(6) => 
        \N0_data[6]\, N0_data(5) => \N0_data[5]\, N0_data(4) => 
        \N0_data[4]\, N0_data(3) => \N0_data[3]\, N0_data(2) => 
        \N0_data[2]\, N0_data(1) => \N0_data[1]\, 
        SHA256_BLOCK_0_H1_o(31) => SHA256_BLOCK_0_H1_o(31), 
        SHA256_BLOCK_0_H1_o(30) => SHA256_BLOCK_0_H1_o(30), 
        SHA256_BLOCK_0_H1_o(29) => SHA256_BLOCK_0_H1_o(29), 
        SHA256_BLOCK_0_H1_o(28) => SHA256_BLOCK_0_H1_o(28), 
        SHA256_BLOCK_0_H1_o(27) => SHA256_BLOCK_0_H1_o(27), 
        SHA256_BLOCK_0_H1_o(26) => SHA256_BLOCK_0_H1_o(26), 
        SHA256_BLOCK_0_H1_o(25) => SHA256_BLOCK_0_H1_o(25), 
        SHA256_BLOCK_0_H1_o(24) => SHA256_BLOCK_0_H1_o(24), 
        SHA256_BLOCK_0_H1_o(23) => SHA256_BLOCK_0_H1_o(23), 
        SHA256_BLOCK_0_H1_o(22) => SHA256_BLOCK_0_H1_o(22), 
        SHA256_BLOCK_0_H1_o(21) => SHA256_BLOCK_0_H1_o(21), 
        SHA256_BLOCK_0_H1_o(20) => SHA256_BLOCK_0_H1_o(20), 
        SHA256_BLOCK_0_H1_o(19) => SHA256_BLOCK_0_H1_o(19), 
        SHA256_BLOCK_0_H1_o(18) => SHA256_BLOCK_0_H1_o(18), 
        SHA256_BLOCK_0_H1_o(17) => SHA256_BLOCK_0_H1_o(17), 
        SHA256_BLOCK_0_H1_o(16) => SHA256_BLOCK_0_H1_o(16), 
        SHA256_BLOCK_0_H1_o(15) => SHA256_BLOCK_0_H1_o(15), 
        SHA256_BLOCK_0_H1_o(14) => SHA256_BLOCK_0_H1_o(14), 
        SHA256_BLOCK_0_H1_o(13) => SHA256_BLOCK_0_H1_o(13), 
        SHA256_BLOCK_0_H1_o(12) => SHA256_BLOCK_0_H1_o(12), 
        SHA256_BLOCK_0_H1_o(11) => SHA256_BLOCK_0_H1_o(11), 
        SHA256_BLOCK_0_H1_o(10) => SHA256_BLOCK_0_H1_o(10), 
        SHA256_BLOCK_0_H1_o(9) => SHA256_BLOCK_0_H1_o(9), 
        SHA256_BLOCK_0_H1_o(8) => SHA256_BLOCK_0_H1_o(8), 
        SHA256_BLOCK_0_H1_o(7) => SHA256_BLOCK_0_H1_o(7), 
        SHA256_BLOCK_0_H1_o(6) => SHA256_BLOCK_0_H1_o(6), 
        SHA256_BLOCK_0_H1_o(5) => SHA256_BLOCK_0_H1_o(5), 
        SHA256_BLOCK_0_H1_o(4) => SHA256_BLOCK_0_H1_o(4), 
        SHA256_BLOCK_0_H1_o(3) => SHA256_BLOCK_0_H1_o(3), 
        SHA256_BLOCK_0_H1_o(2) => SHA256_BLOCK_0_H1_o(2), 
        SHA256_BLOCK_0_H1_o(1) => SHA256_BLOCK_0_H1_o(1), 
        SHA256_BLOCK_0_H1_o(0) => SHA256_BLOCK_0_H1_o(0), 
        N1_data(31) => \N1_data[31]\, N1_data(30) => 
        \N1_data[30]\, N1_data(29) => \N1_data[29]\, N1_data(28)
         => \N1_data[28]\, N1_data(27) => \N1_data[27]\, 
        N1_data(26) => \N1_data[26]\, N1_data(25) => 
        \N1_data[25]\, N1_data(24) => \N1_data[24]\, N1_data(23)
         => \N1_data[23]\, N1_data(22) => \N1_data[22]\, 
        N1_data(21) => \N1_data[21]\, N1_data(20) => 
        \N1_data[20]\, N1_data(19) => \N1_data[19]\, N1_data(18)
         => \N1_data[18]\, N1_data(17) => \N1_data[17]\, 
        N1_data(16) => \N1_data[16]\, N1_data(15) => 
        \N1_data[15]\, N1_data(14) => \N1_data[14]\, N1_data(13)
         => \N1_data[13]\, N1_data(12) => \N1_data[12]\, 
        N1_data(11) => \N1_data[11]\, N1_data(10) => 
        \N1_data[10]\, N1_data(9) => \N1_data[9]\, N1_data(8) => 
        \N1_data[8]\, N1_data(7) => \N1_data[7]\, N1_data(6) => 
        \N1_data[6]\, N1_data(5) => \N1_data[5]\, N1_data(4) => 
        \N1_data[4]\, N1_data(3) => \N1_data[3]\, N1_data(2) => 
        \N1_data[2]\, N1_data(1) => \N1_data[1]\, 
        SHA256_BLOCK_0_H2_o(31) => SHA256_BLOCK_0_H2_o(31), 
        SHA256_BLOCK_0_H2_o(30) => SHA256_BLOCK_0_H2_o(30), 
        SHA256_BLOCK_0_H2_o(29) => SHA256_BLOCK_0_H2_o(29), 
        SHA256_BLOCK_0_H2_o(28) => SHA256_BLOCK_0_H2_o(28), 
        SHA256_BLOCK_0_H2_o(27) => SHA256_BLOCK_0_H2_o(27), 
        SHA256_BLOCK_0_H2_o(26) => SHA256_BLOCK_0_H2_o(26), 
        SHA256_BLOCK_0_H2_o(25) => SHA256_BLOCK_0_H2_o(25), 
        SHA256_BLOCK_0_H2_o(24) => SHA256_BLOCK_0_H2_o(24), 
        SHA256_BLOCK_0_H2_o(23) => SHA256_BLOCK_0_H2_o(23), 
        SHA256_BLOCK_0_H2_o(22) => SHA256_BLOCK_0_H2_o(22), 
        SHA256_BLOCK_0_H2_o(21) => SHA256_BLOCK_0_H2_o(21), 
        SHA256_BLOCK_0_H2_o(20) => SHA256_BLOCK_0_H2_o(20), 
        SHA256_BLOCK_0_H2_o(19) => SHA256_BLOCK_0_H2_o(19), 
        SHA256_BLOCK_0_H2_o(18) => SHA256_BLOCK_0_H2_o(18), 
        SHA256_BLOCK_0_H2_o(17) => SHA256_BLOCK_0_H2_o(17), 
        SHA256_BLOCK_0_H2_o(16) => SHA256_BLOCK_0_H2_o(16), 
        SHA256_BLOCK_0_H2_o(15) => SHA256_BLOCK_0_H2_o(15), 
        SHA256_BLOCK_0_H2_o(14) => SHA256_BLOCK_0_H2_o(14), 
        SHA256_BLOCK_0_H2_o(13) => SHA256_BLOCK_0_H2_o(13), 
        SHA256_BLOCK_0_H2_o(12) => SHA256_BLOCK_0_H2_o(12), 
        SHA256_BLOCK_0_H2_o(11) => SHA256_BLOCK_0_H2_o(11), 
        SHA256_BLOCK_0_H2_o(10) => SHA256_BLOCK_0_H2_o(10), 
        SHA256_BLOCK_0_H2_o(9) => SHA256_BLOCK_0_H2_o(9), 
        SHA256_BLOCK_0_H2_o(8) => SHA256_BLOCK_0_H2_o(8), 
        SHA256_BLOCK_0_H2_o(7) => SHA256_BLOCK_0_H2_o(7), 
        SHA256_BLOCK_0_H2_o(6) => SHA256_BLOCK_0_H2_o(6), 
        SHA256_BLOCK_0_H2_o(5) => SHA256_BLOCK_0_H2_o(5), 
        SHA256_BLOCK_0_H2_o(4) => SHA256_BLOCK_0_H2_o(4), 
        SHA256_BLOCK_0_H2_o(3) => SHA256_BLOCK_0_H2_o(3), 
        SHA256_BLOCK_0_H2_o(2) => SHA256_BLOCK_0_H2_o(2), 
        SHA256_BLOCK_0_H2_o(1) => SHA256_BLOCK_0_H2_o(1), 
        SHA256_BLOCK_0_H2_o(0) => SHA256_BLOCK_0_H2_o(0), 
        N2_data(31) => \N2_data[31]\, N2_data(30) => 
        \N2_data[30]\, N2_data(29) => \N2_data[29]\, N2_data(28)
         => \N2_data[28]\, N2_data(27) => \N2_data[27]\, 
        N2_data(26) => \N2_data[26]\, N2_data(25) => 
        \N2_data[25]\, N2_data(24) => \N2_data[24]\, N2_data(23)
         => \N2_data[23]\, N2_data(22) => \N2_data[22]\, 
        N2_data(21) => \N2_data[21]\, N2_data(20) => 
        \N2_data[20]\, N2_data(19) => \N2_data[19]\, N2_data(18)
         => \N2_data[18]\, N2_data(17) => \N2_data[17]\, 
        N2_data(16) => \N2_data[16]\, N2_data(15) => 
        \N2_data[15]\, N2_data(14) => \N2_data[14]\, N2_data(13)
         => \N2_data[13]\, N2_data(12) => \N2_data[12]\, 
        N2_data(11) => \N2_data[11]\, N2_data(10) => 
        \N2_data[10]\, N2_data(9) => \N2_data[9]\, N2_data(8) => 
        \N2_data[8]\, N2_data(7) => \N2_data[7]\, N2_data(6) => 
        \N2_data[6]\, N2_data(5) => \N2_data[5]\, N2_data(4) => 
        \N2_data[4]\, N2_data(3) => \N2_data[3]\, N2_data(2) => 
        \N2_data[2]\, N2_data(1) => \N2_data[1]\, 
        SHA256_BLOCK_0_H3_o(31) => SHA256_BLOCK_0_H3_o(31), 
        SHA256_BLOCK_0_H3_o(30) => SHA256_BLOCK_0_H3_o(30), 
        SHA256_BLOCK_0_H3_o(29) => SHA256_BLOCK_0_H3_o(29), 
        SHA256_BLOCK_0_H3_o(28) => SHA256_BLOCK_0_H3_o(28), 
        SHA256_BLOCK_0_H3_o(27) => SHA256_BLOCK_0_H3_o(27), 
        SHA256_BLOCK_0_H3_o(26) => SHA256_BLOCK_0_H3_o(26), 
        SHA256_BLOCK_0_H3_o(25) => SHA256_BLOCK_0_H3_o(25), 
        SHA256_BLOCK_0_H3_o(24) => SHA256_BLOCK_0_H3_o(24), 
        SHA256_BLOCK_0_H3_o(23) => SHA256_BLOCK_0_H3_o(23), 
        SHA256_BLOCK_0_H3_o(22) => SHA256_BLOCK_0_H3_o(22), 
        SHA256_BLOCK_0_H3_o(21) => SHA256_BLOCK_0_H3_o(21), 
        SHA256_BLOCK_0_H3_o(20) => SHA256_BLOCK_0_H3_o(20), 
        SHA256_BLOCK_0_H3_o(19) => SHA256_BLOCK_0_H3_o(19), 
        SHA256_BLOCK_0_H3_o(18) => SHA256_BLOCK_0_H3_o(18), 
        SHA256_BLOCK_0_H3_o(17) => SHA256_BLOCK_0_H3_o(17), 
        SHA256_BLOCK_0_H3_o(16) => SHA256_BLOCK_0_H3_o(16), 
        SHA256_BLOCK_0_H3_o(15) => SHA256_BLOCK_0_H3_o(15), 
        SHA256_BLOCK_0_H3_o(14) => SHA256_BLOCK_0_H3_o(14), 
        SHA256_BLOCK_0_H3_o(13) => SHA256_BLOCK_0_H3_o(13), 
        SHA256_BLOCK_0_H3_o(12) => SHA256_BLOCK_0_H3_o(12), 
        SHA256_BLOCK_0_H3_o(11) => SHA256_BLOCK_0_H3_o(11), 
        SHA256_BLOCK_0_H3_o(10) => SHA256_BLOCK_0_H3_o(10), 
        SHA256_BLOCK_0_H3_o(9) => SHA256_BLOCK_0_H3_o(9), 
        SHA256_BLOCK_0_H3_o(8) => SHA256_BLOCK_0_H3_o(8), 
        SHA256_BLOCK_0_H3_o(7) => SHA256_BLOCK_0_H3_o(7), 
        SHA256_BLOCK_0_H3_o(6) => SHA256_BLOCK_0_H3_o(6), 
        SHA256_BLOCK_0_H3_o(5) => SHA256_BLOCK_0_H3_o(5), 
        SHA256_BLOCK_0_H3_o(4) => SHA256_BLOCK_0_H3_o(4), 
        SHA256_BLOCK_0_H3_o(3) => SHA256_BLOCK_0_H3_o(3), 
        SHA256_BLOCK_0_H3_o(2) => SHA256_BLOCK_0_H3_o(2), 
        SHA256_BLOCK_0_H3_o(1) => SHA256_BLOCK_0_H3_o(1), 
        SHA256_BLOCK_0_H3_o(0) => SHA256_BLOCK_0_H3_o(0), 
        N3_data(31) => \N3_data[31]\, N3_data(30) => 
        \N3_data[30]\, N3_data(29) => \N3_data[29]\, N3_data(28)
         => \N3_data[28]\, N3_data(27) => \N3_data[27]\, 
        N3_data(26) => \N3_data[26]\, N3_data(25) => 
        \N3_data[25]\, N3_data(24) => \N3_data[24]\, N3_data(23)
         => \N3_data[23]\, N3_data(22) => \N3_data[22]\, 
        N3_data(21) => \N3_data[21]\, N3_data(20) => 
        \N3_data[20]\, N3_data(19) => \N3_data[19]\, N3_data(18)
         => \N3_data[18]\, N3_data(17) => \N3_data[17]\, 
        N3_data(16) => \N3_data[16]\, N3_data(15) => 
        \N3_data[15]\, N3_data(14) => \N3_data[14]\, N3_data(13)
         => \N3_data[13]\, N3_data(12) => \N3_data[12]\, 
        N3_data(11) => \N3_data[11]\, N3_data(10) => 
        \N3_data[10]\, N3_data(9) => \N3_data[9]\, N3_data(8) => 
        \N3_data[8]\, N3_data(7) => \N3_data[7]\, N3_data(6) => 
        \N3_data[6]\, N3_data(5) => \N3_data[5]\, N3_data(4) => 
        \N3_data[4]\, N3_data(3) => \N3_data[3]\, N3_data(2) => 
        \N3_data[2]\, N3_data(1) => \N3_data[1]\, 
        SHA256_BLOCK_0_H4_o(31) => SHA256_BLOCK_0_H4_o(31), 
        SHA256_BLOCK_0_H4_o(30) => SHA256_BLOCK_0_H4_o(30), 
        SHA256_BLOCK_0_H4_o(29) => SHA256_BLOCK_0_H4_o(29), 
        SHA256_BLOCK_0_H4_o(28) => SHA256_BLOCK_0_H4_o(28), 
        SHA256_BLOCK_0_H4_o(27) => SHA256_BLOCK_0_H4_o(27), 
        SHA256_BLOCK_0_H4_o(26) => SHA256_BLOCK_0_H4_o(26), 
        SHA256_BLOCK_0_H4_o(25) => SHA256_BLOCK_0_H4_o(25), 
        SHA256_BLOCK_0_H4_o(24) => SHA256_BLOCK_0_H4_o(24), 
        SHA256_BLOCK_0_H4_o(23) => SHA256_BLOCK_0_H4_o(23), 
        SHA256_BLOCK_0_H4_o(22) => SHA256_BLOCK_0_H4_o(22), 
        SHA256_BLOCK_0_H4_o(21) => SHA256_BLOCK_0_H4_o(21), 
        SHA256_BLOCK_0_H4_o(20) => SHA256_BLOCK_0_H4_o(20), 
        SHA256_BLOCK_0_H4_o(19) => SHA256_BLOCK_0_H4_o(19), 
        SHA256_BLOCK_0_H4_o(18) => SHA256_BLOCK_0_H4_o(18), 
        SHA256_BLOCK_0_H4_o(17) => SHA256_BLOCK_0_H4_o(17), 
        SHA256_BLOCK_0_H4_o(16) => SHA256_BLOCK_0_H4_o(16), 
        SHA256_BLOCK_0_H4_o(15) => SHA256_BLOCK_0_H4_o(15), 
        SHA256_BLOCK_0_H4_o(14) => SHA256_BLOCK_0_H4_o(14), 
        SHA256_BLOCK_0_H4_o(13) => SHA256_BLOCK_0_H4_o(13), 
        SHA256_BLOCK_0_H4_o(12) => SHA256_BLOCK_0_H4_o(12), 
        SHA256_BLOCK_0_H4_o(11) => SHA256_BLOCK_0_H4_o(11), 
        SHA256_BLOCK_0_H4_o(10) => SHA256_BLOCK_0_H4_o(10), 
        SHA256_BLOCK_0_H4_o(9) => SHA256_BLOCK_0_H4_o(9), 
        SHA256_BLOCK_0_H4_o(8) => SHA256_BLOCK_0_H4_o(8), 
        SHA256_BLOCK_0_H4_o(7) => SHA256_BLOCK_0_H4_o(7), 
        SHA256_BLOCK_0_H4_o(6) => SHA256_BLOCK_0_H4_o(6), 
        SHA256_BLOCK_0_H4_o(5) => SHA256_BLOCK_0_H4_o(5), 
        SHA256_BLOCK_0_H4_o(4) => SHA256_BLOCK_0_H4_o(4), 
        SHA256_BLOCK_0_H4_o(3) => SHA256_BLOCK_0_H4_o(3), 
        SHA256_BLOCK_0_H4_o(2) => SHA256_BLOCK_0_H4_o(2), 
        SHA256_BLOCK_0_H4_o(1) => SHA256_BLOCK_0_H4_o(1), 
        SHA256_BLOCK_0_H4_o(0) => SHA256_BLOCK_0_H4_o(0), 
        N4_data(31) => \N4_data[31]\, N4_data(30) => 
        \N4_data[30]\, N4_data(29) => \N4_data[29]\, N4_data(28)
         => \N4_data[28]\, N4_data(27) => \N4_data[27]\, 
        N4_data(26) => \N4_data[26]\, N4_data(25) => 
        \N4_data[25]\, N4_data(24) => \N4_data[24]\, N4_data(23)
         => \N4_data[23]\, N4_data(22) => \N4_data[22]\, 
        N4_data(21) => \N4_data[21]\, N4_data(20) => 
        \N4_data[20]\, N4_data(19) => \N4_data[19]\, N4_data(18)
         => \N4_data[18]\, N4_data(17) => \N4_data[17]\, 
        N4_data(16) => \N4_data[16]\, N4_data(15) => 
        \N4_data[15]\, N4_data(14) => \N4_data[14]\, N4_data(13)
         => \N4_data[13]\, N4_data(12) => \N4_data[12]\, 
        N4_data(11) => \N4_data[11]\, N4_data(10) => 
        \N4_data[10]\, N4_data(9) => \N4_data[9]\, N4_data(8) => 
        \N4_data[8]\, N4_data(7) => \N4_data[7]\, N4_data(6) => 
        \N4_data[6]\, N4_data(5) => \N4_data[5]\, N4_data(4) => 
        \N4_data[4]\, N4_data(3) => \N4_data[3]\, N4_data(2) => 
        \N4_data[2]\, N4_data(1) => \N4_data[1]\, N5_data(31) => 
        \N5_data[31]\, N5_data(30) => \N5_data[30]\, N5_data(29)
         => \N5_data[29]\, N5_data(28) => \N5_data[28]\, 
        N5_data(27) => \N5_data[27]\, N5_data(26) => 
        \N5_data[26]\, N5_data(25) => \N5_data[25]\, N5_data(24)
         => \N5_data[24]\, N5_data(23) => \N5_data[23]\, 
        N5_data(22) => \N5_data[22]\, N5_data(21) => 
        \N5_data[21]\, N5_data(20) => \N5_data[20]\, N5_data(19)
         => \N5_data[19]\, N5_data(18) => \N5_data[18]\, 
        N5_data(17) => \N5_data[17]\, N5_data(16) => 
        \N5_data[16]\, N5_data(15) => \N5_data[15]\, N5_data(14)
         => \N5_data[14]\, N5_data(13) => \N5_data[13]\, 
        N5_data(12) => \N5_data[12]\, N5_data(11) => 
        \N5_data[11]\, N5_data(10) => \N5_data[10]\, N5_data(9)
         => \N5_data[9]\, N5_data(8) => \N5_data[8]\, N5_data(7)
         => \N5_data[7]\, N5_data(6) => \N5_data[6]\, N5_data(5)
         => \N5_data[5]\, N5_data(4) => \N5_data[4]\, N5_data(3)
         => \N5_data[3]\, N5_data(2) => \N5_data[2]\, N5_data(1)
         => \N5_data[1]\, SHA256_BLOCK_0_H5_o(31) => 
        SHA256_BLOCK_0_H5_o(31), SHA256_BLOCK_0_H5_o(30) => 
        SHA256_BLOCK_0_H5_o(30), SHA256_BLOCK_0_H5_o(29) => 
        SHA256_BLOCK_0_H5_o(29), SHA256_BLOCK_0_H5_o(28) => 
        SHA256_BLOCK_0_H5_o(28), SHA256_BLOCK_0_H5_o(27) => 
        SHA256_BLOCK_0_H5_o(27), SHA256_BLOCK_0_H5_o(26) => 
        SHA256_BLOCK_0_H5_o(26), SHA256_BLOCK_0_H5_o(25) => 
        SHA256_BLOCK_0_H5_o(25), SHA256_BLOCK_0_H5_o(24) => 
        SHA256_BLOCK_0_H5_o(24), SHA256_BLOCK_0_H5_o(23) => 
        SHA256_BLOCK_0_H5_o(23), SHA256_BLOCK_0_H5_o(22) => 
        SHA256_BLOCK_0_H5_o(22), SHA256_BLOCK_0_H5_o(21) => 
        SHA256_BLOCK_0_H5_o(21), SHA256_BLOCK_0_H5_o(20) => 
        SHA256_BLOCK_0_H5_o(20), SHA256_BLOCK_0_H5_o(19) => 
        SHA256_BLOCK_0_H5_o(19), SHA256_BLOCK_0_H5_o(18) => 
        SHA256_BLOCK_0_H5_o(18), SHA256_BLOCK_0_H5_o(17) => 
        SHA256_BLOCK_0_H5_o(17), SHA256_BLOCK_0_H5_o(16) => 
        SHA256_BLOCK_0_H5_o(16), SHA256_BLOCK_0_H5_o(15) => 
        SHA256_BLOCK_0_H5_o(15), SHA256_BLOCK_0_H5_o(14) => 
        SHA256_BLOCK_0_H5_o(14), SHA256_BLOCK_0_H5_o(13) => 
        SHA256_BLOCK_0_H5_o(13), SHA256_BLOCK_0_H5_o(12) => 
        SHA256_BLOCK_0_H5_o(12), SHA256_BLOCK_0_H5_o(11) => 
        SHA256_BLOCK_0_H5_o(11), SHA256_BLOCK_0_H5_o(10) => 
        SHA256_BLOCK_0_H5_o(10), SHA256_BLOCK_0_H5_o(9) => 
        SHA256_BLOCK_0_H5_o(9), SHA256_BLOCK_0_H5_o(8) => 
        SHA256_BLOCK_0_H5_o(8), SHA256_BLOCK_0_H5_o(7) => 
        SHA256_BLOCK_0_H5_o(7), SHA256_BLOCK_0_H5_o(6) => 
        SHA256_BLOCK_0_H5_o(6), SHA256_BLOCK_0_H5_o(5) => 
        SHA256_BLOCK_0_H5_o(5), SHA256_BLOCK_0_H5_o(4) => 
        SHA256_BLOCK_0_H5_o(4), SHA256_BLOCK_0_H5_o(3) => 
        SHA256_BLOCK_0_H5_o(3), SHA256_BLOCK_0_H5_o(2) => 
        SHA256_BLOCK_0_H5_o(2), SHA256_BLOCK_0_H5_o(1) => 
        SHA256_BLOCK_0_H5_o(1), SHA256_BLOCK_0_H5_o(0) => 
        SHA256_BLOCK_0_H5_o(0), SHA256_BLOCK_0_H6_o(31) => 
        SHA256_BLOCK_0_H6_o(31), SHA256_BLOCK_0_H6_o(30) => 
        SHA256_BLOCK_0_H6_o(30), SHA256_BLOCK_0_H6_o(29) => 
        SHA256_BLOCK_0_H6_o(29), SHA256_BLOCK_0_H6_o(28) => 
        SHA256_BLOCK_0_H6_o(28), SHA256_BLOCK_0_H6_o(27) => 
        SHA256_BLOCK_0_H6_o(27), SHA256_BLOCK_0_H6_o(26) => 
        SHA256_BLOCK_0_H6_o(26), SHA256_BLOCK_0_H6_o(25) => 
        SHA256_BLOCK_0_H6_o(25), SHA256_BLOCK_0_H6_o(24) => 
        SHA256_BLOCK_0_H6_o(24), SHA256_BLOCK_0_H6_o(23) => 
        SHA256_BLOCK_0_H6_o(23), SHA256_BLOCK_0_H6_o(22) => 
        SHA256_BLOCK_0_H6_o(22), SHA256_BLOCK_0_H6_o(21) => 
        SHA256_BLOCK_0_H6_o(21), SHA256_BLOCK_0_H6_o(20) => 
        SHA256_BLOCK_0_H6_o(20), SHA256_BLOCK_0_H6_o(19) => 
        SHA256_BLOCK_0_H6_o(19), SHA256_BLOCK_0_H6_o(18) => 
        SHA256_BLOCK_0_H6_o(18), SHA256_BLOCK_0_H6_o(17) => 
        SHA256_BLOCK_0_H6_o(17), SHA256_BLOCK_0_H6_o(16) => 
        SHA256_BLOCK_0_H6_o(16), SHA256_BLOCK_0_H6_o(15) => 
        SHA256_BLOCK_0_H6_o(15), SHA256_BLOCK_0_H6_o(14) => 
        SHA256_BLOCK_0_H6_o(14), SHA256_BLOCK_0_H6_o(13) => 
        SHA256_BLOCK_0_H6_o(13), SHA256_BLOCK_0_H6_o(12) => 
        SHA256_BLOCK_0_H6_o(12), SHA256_BLOCK_0_H6_o(11) => 
        SHA256_BLOCK_0_H6_o(11), SHA256_BLOCK_0_H6_o(10) => 
        SHA256_BLOCK_0_H6_o(10), SHA256_BLOCK_0_H6_o(9) => 
        SHA256_BLOCK_0_H6_o(9), SHA256_BLOCK_0_H6_o(8) => 
        SHA256_BLOCK_0_H6_o(8), SHA256_BLOCK_0_H6_o(7) => 
        SHA256_BLOCK_0_H6_o(7), SHA256_BLOCK_0_H6_o(6) => 
        SHA256_BLOCK_0_H6_o(6), SHA256_BLOCK_0_H6_o(5) => 
        SHA256_BLOCK_0_H6_o(5), SHA256_BLOCK_0_H6_o(4) => 
        SHA256_BLOCK_0_H6_o(4), SHA256_BLOCK_0_H6_o(3) => 
        SHA256_BLOCK_0_H6_o(3), SHA256_BLOCK_0_H6_o(2) => 
        SHA256_BLOCK_0_H6_o(2), SHA256_BLOCK_0_H6_o(1) => 
        SHA256_BLOCK_0_H6_o(1), SHA256_BLOCK_0_H6_o(0) => 
        SHA256_BLOCK_0_H6_o(0), N6_data(31) => \N6_data[31]\, 
        N6_data(30) => \N6_data[30]\, N6_data(29) => 
        \N6_data[29]\, N6_data(28) => \N6_data[28]\, N6_data(27)
         => \N6_data[27]\, N6_data(26) => \N6_data[26]\, 
        N6_data(25) => \N6_data[25]\, N6_data(24) => 
        \N6_data[24]\, N6_data(23) => \N6_data[23]\, N6_data(22)
         => \N6_data[22]\, N6_data(21) => \N6_data[21]\, 
        N6_data(20) => \N6_data[20]\, N6_data(19) => 
        \N6_data[19]\, N6_data(18) => \N6_data[18]\, N6_data(17)
         => \N6_data[17]\, N6_data(16) => \N6_data[16]\, 
        N6_data(15) => \N6_data[15]\, N6_data(14) => 
        \N6_data[14]\, N6_data(13) => \N6_data[13]\, N6_data(12)
         => \N6_data[12]\, N6_data(11) => \N6_data[11]\, 
        N6_data(10) => \N6_data[10]\, N6_data(9) => \N6_data[9]\, 
        N6_data(8) => \N6_data[8]\, N6_data(7) => \N6_data[7]\, 
        N6_data(6) => \N6_data[6]\, N6_data(5) => \N6_data[5]\, 
        N6_data(4) => \N6_data[4]\, N6_data(3) => \N6_data[3]\, 
        N6_data(2) => \N6_data[2]\, N6_data(1) => \N6_data[1]\, 
        SHA256_BLOCK_0_H7_o(31) => SHA256_BLOCK_0_H7_o(31), 
        SHA256_BLOCK_0_H7_o(30) => SHA256_BLOCK_0_H7_o(30), 
        SHA256_BLOCK_0_H7_o(29) => SHA256_BLOCK_0_H7_o(29), 
        SHA256_BLOCK_0_H7_o(28) => SHA256_BLOCK_0_H7_o(28), 
        SHA256_BLOCK_0_H7_o(27) => SHA256_BLOCK_0_H7_o(27), 
        SHA256_BLOCK_0_H7_o(26) => SHA256_BLOCK_0_H7_o(26), 
        SHA256_BLOCK_0_H7_o(25) => SHA256_BLOCK_0_H7_o(25), 
        SHA256_BLOCK_0_H7_o(24) => SHA256_BLOCK_0_H7_o(24), 
        SHA256_BLOCK_0_H7_o(23) => SHA256_BLOCK_0_H7_o(23), 
        SHA256_BLOCK_0_H7_o(22) => SHA256_BLOCK_0_H7_o(22), 
        SHA256_BLOCK_0_H7_o(21) => SHA256_BLOCK_0_H7_o(21), 
        SHA256_BLOCK_0_H7_o(20) => SHA256_BLOCK_0_H7_o(20), 
        SHA256_BLOCK_0_H7_o(19) => SHA256_BLOCK_0_H7_o(19), 
        SHA256_BLOCK_0_H7_o(18) => SHA256_BLOCK_0_H7_o(18), 
        SHA256_BLOCK_0_H7_o(17) => SHA256_BLOCK_0_H7_o(17), 
        SHA256_BLOCK_0_H7_o(16) => SHA256_BLOCK_0_H7_o(16), 
        SHA256_BLOCK_0_H7_o(15) => SHA256_BLOCK_0_H7_o(15), 
        SHA256_BLOCK_0_H7_o(14) => SHA256_BLOCK_0_H7_o(14), 
        SHA256_BLOCK_0_H7_o(13) => SHA256_BLOCK_0_H7_o(13), 
        SHA256_BLOCK_0_H7_o(12) => SHA256_BLOCK_0_H7_o(12), 
        SHA256_BLOCK_0_H7_o(11) => SHA256_BLOCK_0_H7_o(11), 
        SHA256_BLOCK_0_H7_o(10) => SHA256_BLOCK_0_H7_o(10), 
        SHA256_BLOCK_0_H7_o(9) => SHA256_BLOCK_0_H7_o(9), 
        SHA256_BLOCK_0_H7_o(8) => SHA256_BLOCK_0_H7_o(8), 
        SHA256_BLOCK_0_H7_o(7) => SHA256_BLOCK_0_H7_o(7), 
        SHA256_BLOCK_0_H7_o(6) => SHA256_BLOCK_0_H7_o(6), 
        SHA256_BLOCK_0_H7_o(5) => SHA256_BLOCK_0_H7_o(5), 
        SHA256_BLOCK_0_H7_o(4) => SHA256_BLOCK_0_H7_o(4), 
        SHA256_BLOCK_0_H7_o(3) => SHA256_BLOCK_0_H7_o(3), 
        SHA256_BLOCK_0_H7_o(2) => SHA256_BLOCK_0_H7_o(2), 
        SHA256_BLOCK_0_H7_o(1) => SHA256_BLOCK_0_H7_o(1), 
        SHA256_BLOCK_0_H7_o(0) => SHA256_BLOCK_0_H7_o(0), 
        N7_data(31) => \N7_data[31]\, N7_data(30) => 
        \N7_data[30]\, N7_data(29) => \N7_data[29]\, N7_data(28)
         => \N7_data[28]\, N7_data(27) => \N7_data[27]\, 
        N7_data(26) => \N7_data[26]\, N7_data(25) => 
        \N7_data[25]\, N7_data(24) => \N7_data[24]\, N7_data(23)
         => \N7_data[23]\, N7_data(22) => \N7_data[22]\, 
        N7_data(21) => \N7_data[21]\, N7_data(20) => 
        \N7_data[20]\, N7_data(19) => \N7_data[19]\, N7_data(18)
         => \N7_data[18]\, N7_data(17) => \N7_data[17]\, 
        N7_data(16) => \N7_data[16]\, N7_data(15) => 
        \N7_data[15]\, N7_data(14) => \N7_data[14]\, N7_data(13)
         => \N7_data[13]\, N7_data(12) => \N7_data[12]\, 
        N7_data(11) => \N7_data[11]\, N7_data(10) => 
        \N7_data[10]\, N7_data(9) => \N7_data[9]\, N7_data(8) => 
        \N7_data[8]\, N7_data(7) => \N7_data[7]\, N7_data(6) => 
        \N7_data[6]\, N7_data(5) => \N7_data[5]\, N7_data(4) => 
        \N7_data[4]\, N7_data(3) => \N7_data[3]\, N7_data(2) => 
        \N7_data[2]\, N7_data(1) => \N7_data[1]\, 
        hash_control_st_reg_i(6) => \hash_control_st_reg_i[6]\, 
        R0_data(31) => \R0_data[31]\, R0_data(30) => 
        \R0_data[30]\, R0_data(29) => \R0_data[29]\, R0_data(28)
         => \R0_data[28]\, R0_data(27) => \R0_data[27]\, 
        R0_data(26) => \R0_data[26]\, R0_data(25) => 
        \R0_data[25]\, R0_data(24) => \R0_data[24]\, R0_data(23)
         => \R0_data[23]\, R0_data(22) => \R0_data[22]\, 
        R0_data(21) => \R0_data[21]\, R0_data(20) => 
        \R0_data[20]\, R0_data(19) => \R0_data[19]\, R0_data(18)
         => \R0_data[18]\, R0_data(17) => \R0_data[17]\, 
        R0_data(16) => \R0_data[16]\, R0_data(15) => 
        \R0_data[15]\, R0_data(14) => \R0_data[14]\, R0_data(13)
         => \R0_data[13]\, R0_data(12) => \R0_data[12]\, 
        R0_data(11) => \R0_data[11]\, R0_data(10) => 
        \R0_data[10]\, R0_data(9) => \R0_data[9]\, R0_data(8) => 
        \R0_data[8]\, R0_data(7) => \R0_data[7]\, R0_data(6) => 
        \R0_data[6]\, R0_data(5) => \R0_data[5]\, R0_data(4) => 
        \R0_data[4]\, R0_data(3) => \R0_data[3]\, R0_data(2) => 
        \R0_data[2]\, R0_data(1) => \R0_data[1]\, R0_data(0) => 
        \R0_data[0]\, R1_data(31) => \R1_data[31]\, R1_data(30)
         => \R1_data[30]\, R1_data(29) => \R1_data[29]\, 
        R1_data(28) => \R1_data[28]\, R1_data(27) => 
        \R1_data[27]\, R1_data(26) => \R1_data[26]\, R1_data(25)
         => \R1_data[25]\, R1_data(24) => \R1_data[24]\, 
        R1_data(23) => \R1_data[23]\, R1_data(22) => 
        \R1_data[22]\, R1_data(21) => \R1_data[21]\, R1_data(20)
         => \R1_data[20]\, R1_data(19) => \R1_data[19]\, 
        R1_data(18) => \R1_data[18]\, R1_data(17) => 
        \R1_data[17]\, R1_data(16) => \R1_data[16]\, R1_data(15)
         => \R1_data[15]\, R1_data(14) => \R1_data[14]\, 
        R1_data(13) => \R1_data[13]\, R1_data(12) => 
        \R1_data[12]\, R1_data(11) => \R1_data[11]\, R1_data(10)
         => \R1_data[10]\, R1_data(9) => \R1_data[9]\, R1_data(8)
         => \R1_data[8]\, R1_data(7) => \R1_data[7]\, R1_data(6)
         => \R1_data[6]\, R1_data(5) => \R1_data[5]\, R1_data(4)
         => \R1_data[4]\, R1_data(3) => \R1_data[3]\, R1_data(2)
         => \R1_data[2]\, R1_data(1) => \R1_data[1]\, R1_data(0)
         => \R1_data[0]\, R2_data(31) => \R2_data[31]\, 
        R2_data(30) => \R2_data[30]\, R2_data(29) => 
        \R2_data[29]\, R2_data(28) => \R2_data[28]\, R2_data(27)
         => \R2_data[27]\, R2_data(26) => \R2_data[26]\, 
        R2_data(25) => \R2_data[25]\, R2_data(24) => 
        \R2_data[24]\, R2_data(23) => \R2_data[23]\, R2_data(22)
         => \R2_data[22]\, R2_data(21) => \R2_data[21]\, 
        R2_data(20) => \R2_data[20]\, R2_data(19) => 
        \R2_data[19]\, R2_data(18) => \R2_data[18]\, R2_data(17)
         => \R2_data[17]\, R2_data(16) => \R2_data[16]\, 
        R2_data(15) => \R2_data[15]\, R2_data(14) => 
        \R2_data[14]\, R2_data(13) => \R2_data[13]\, R2_data(12)
         => \R2_data[12]\, R2_data(11) => \R2_data[11]\, 
        R2_data(10) => \R2_data[10]\, R2_data(9) => \R2_data[9]\, 
        R2_data(8) => \R2_data[8]\, R2_data(7) => \R2_data[7]\, 
        R2_data(6) => \R2_data[6]\, R2_data(5) => \R2_data[5]\, 
        R2_data(4) => \R2_data[4]\, R2_data(3) => \R2_data[3]\, 
        R2_data(2) => \R2_data[2]\, R2_data(1) => \R2_data[1]\, 
        R2_data(0) => \R2_data[0]\, R3_data(31) => \R3_data[31]\, 
        R3_data(30) => \R3_data[30]\, R3_data(29) => 
        \R3_data[29]\, R3_data(28) => \R3_data[28]\, R3_data(27)
         => \R3_data[27]\, R3_data(26) => \R3_data[26]\, 
        R3_data(25) => \R3_data[25]\, R3_data(24) => 
        \R3_data[24]\, R3_data(23) => \R3_data[23]\, R3_data(22)
         => \R3_data[22]\, R3_data(21) => \R3_data[21]\, 
        R3_data(20) => \R3_data[20]\, R3_data(19) => 
        \R3_data[19]\, R3_data(18) => \R3_data[18]\, R3_data(17)
         => \R3_data[17]\, R3_data(16) => \R3_data[16]\, 
        R3_data(15) => \R3_data[15]\, R3_data(14) => 
        \R3_data[14]\, R3_data(13) => \R3_data[13]\, R3_data(12)
         => \R3_data[12]\, R3_data(11) => \R3_data[11]\, 
        R3_data(10) => \R3_data[10]\, R3_data(9) => \R3_data[9]\, 
        R3_data(8) => \R3_data[8]\, R3_data(7) => \R3_data[7]\, 
        R3_data(6) => \R3_data[6]\, R3_data(5) => \R3_data[5]\, 
        R3_data(4) => \R3_data[4]\, R3_data(3) => \R3_data[3]\, 
        R3_data(2) => \R3_data[2]\, R3_data(1) => \R3_data[1]\, 
        R3_data(0) => \R3_data[0]\, R4_data(31) => \R4_data[31]\, 
        R4_data(30) => \R4_data[30]\, R4_data(29) => 
        \R4_data[29]\, R4_data(28) => \R4_data[28]\, R4_data(27)
         => \R4_data[27]\, R4_data(26) => \R4_data[26]\, 
        R4_data(25) => \R4_data[25]\, R4_data(24) => 
        \R4_data[24]\, R4_data(23) => \R4_data[23]\, R4_data(22)
         => \R4_data[22]\, R4_data(21) => \R4_data[21]\, 
        R4_data(20) => \R4_data[20]\, R4_data(19) => 
        \R4_data[19]\, R4_data(18) => \R4_data[18]\, R4_data(17)
         => \R4_data[17]\, R4_data(16) => \R4_data[16]\, 
        R4_data(15) => \R4_data[15]\, R4_data(14) => 
        \R4_data[14]\, R4_data(13) => \R4_data[13]\, R4_data(12)
         => \R4_data[12]\, R4_data(11) => \R4_data[11]\, 
        R4_data(10) => \R4_data[10]\, R4_data(9) => \R4_data[9]\, 
        R4_data(8) => \R4_data[8]\, R4_data(7) => \R4_data[7]\, 
        R4_data(6) => \R4_data[6]\, R4_data(5) => \R4_data[5]\, 
        R4_data(4) => \R4_data[4]\, R4_data(3) => \R4_data[3]\, 
        R4_data(2) => \R4_data[2]\, R4_data(1) => \R4_data[1]\, 
        R4_data(0) => \R4_data[0]\, R5_data(31) => \R5_data[31]\, 
        R5_data(30) => \R5_data[30]\, R5_data(29) => 
        \R5_data[29]\, R5_data(28) => \R5_data[28]\, R5_data(27)
         => \R5_data[27]\, R5_data(26) => \R5_data[26]\, 
        R5_data(25) => \R5_data[25]\, R5_data(24) => 
        \R5_data[24]\, R5_data(23) => \R5_data[23]\, R5_data(22)
         => \R5_data[22]\, R5_data(21) => \R5_data[21]\, 
        R5_data(20) => \R5_data[20]\, R5_data(19) => 
        \R5_data[19]\, R5_data(18) => \R5_data[18]\, R5_data(17)
         => \R5_data[17]\, R5_data(16) => \R5_data[16]\, 
        R5_data(15) => \R5_data[15]\, R5_data(14) => 
        \R5_data[14]\, R5_data(13) => \R5_data[13]\, R5_data(12)
         => \R5_data[12]\, R5_data(11) => \R5_data[11]\, 
        R5_data(10) => \R5_data[10]\, R5_data(9) => \R5_data[9]\, 
        R5_data(8) => \R5_data[8]\, R5_data(7) => \R5_data[7]\, 
        R5_data(6) => \R5_data[6]\, R5_data(5) => \R5_data[5]\, 
        R5_data(4) => \R5_data[4]\, R5_data(3) => \R5_data[3]\, 
        R5_data(2) => \R5_data[2]\, R5_data(1) => \R5_data[1]\, 
        R5_data(0) => \R5_data[0]\, R6_data(31) => \R6_data[31]\, 
        R6_data(30) => \R6_data[30]\, R6_data(29) => 
        \R6_data[29]\, R6_data(28) => \R6_data[28]\, R6_data(27)
         => \R6_data[27]\, R6_data(26) => \R6_data[26]\, 
        R6_data(25) => \R6_data[25]\, R6_data(24) => 
        \R6_data[24]\, R6_data(23) => \R6_data[23]\, R6_data(22)
         => \R6_data[22]\, R6_data(21) => \R6_data[21]\, 
        R6_data(20) => \R6_data[20]\, R6_data(19) => 
        \R6_data[19]\, R6_data(18) => \R6_data[18]\, R6_data(17)
         => \R6_data[17]\, R6_data(16) => \R6_data[16]\, 
        R6_data(15) => \R6_data[15]\, R6_data(14) => 
        \R6_data[14]\, R6_data(13) => \R6_data[13]\, R6_data(12)
         => \R6_data[12]\, R6_data(11) => \R6_data[11]\, 
        R6_data(10) => \R6_data[10]\, R6_data(9) => \R6_data[9]\, 
        R6_data(8) => \R6_data[8]\, R6_data(7) => \R6_data[7]\, 
        R6_data(6) => \R6_data[6]\, R6_data(5) => \R6_data[5]\, 
        R6_data(4) => \R6_data[4]\, R6_data(3) => \R6_data[3]\, 
        R6_data(2) => \R6_data[2]\, R6_data(1) => \R6_data[1]\, 
        R6_data(0) => \R6_data[0]\, R7_data(31) => \R7_data[31]\, 
        R7_data(30) => \R7_data[30]\, R7_data(29) => 
        \R7_data[29]\, R7_data(28) => \R7_data[28]\, R7_data(27)
         => \R7_data[27]\, R7_data(26) => \R7_data[26]\, 
        R7_data(25) => \R7_data[25]\, R7_data(24) => 
        \R7_data[24]\, R7_data(23) => \R7_data[23]\, R7_data(22)
         => \R7_data[22]\, R7_data(21) => \R7_data[21]\, 
        R7_data(20) => \R7_data[20]\, R7_data(19) => 
        \R7_data[19]\, R7_data(18) => \R7_data[18]\, R7_data(17)
         => \R7_data[17]\, R7_data(16) => \R7_data[16]\, 
        R7_data(15) => \R7_data[15]\, R7_data(14) => 
        \R7_data[14]\, R7_data(13) => \R7_data[13]\, R7_data(12)
         => \R7_data[12]\, R7_data(11) => \R7_data[11]\, 
        R7_data(10) => \R7_data[10]\, R7_data(9) => \R7_data[9]\, 
        R7_data(8) => \R7_data[8]\, R7_data(7) => \R7_data[7]\, 
        R7_data(6) => \R7_data[6]\, R7_data(5) => \R7_data[5]\, 
        R7_data(4) => \R7_data[4]\, R7_data(3) => \R7_data[3]\, 
        R7_data(2) => \R7_data[2]\, R7_data(1) => \R7_data[1]\, 
        R7_data(0) => \R7_data[0]\, sha256_system_sb_0_FIC_0_CLK
         => sha256_system_sb_0_FIC_0_CLK, N_168_i_0 => N_168_i_0, 
        next_reg_H0_cry_0_0_Y => next_reg_H0_cry_0_0_Y, 
        next_reg_H1_cry_0_0_Y => next_reg_H1_cry_0_0_Y, 
        next_reg_H2_cry_0_0_Y => next_reg_H2_cry_0_0_Y, 
        next_reg_H3_cry_0_0_Y => next_reg_H3_cry_0_0_Y, 
        next_reg_H4_cry_0_0_Y => next_reg_H4_cry_0_0_Y, 
        next_reg_H5_cry_0_0_Y => next_reg_H5_cry_0_0_Y, 
        next_reg_H6_cry_0_0_Y => next_reg_H6_cry_0_0_Y, 
        next_reg_H7_cry_0_0_Y => next_reg_H7_cry_0_0_Y);
    
    Inst_sha256_padding : sha256_padding
      port map(raddr_pos(3) => raddr_pos(3), raddr_pos(2) => 
        raddr_pos(2), Kt_addr(0) => \Kt_addr[0]\, st_cnt_reg(6)
         => \st_cnt_reg[6]\, hash_control_st_reg(2) => 
        \hash_control_st_reg[2]\, Kt_addr_fast(5) => 
        \Kt_addr_fast[5]\, Kt_addr_fast(4) => \Kt_addr_fast[4]\, 
        Kt_addr_fast(3) => \Kt_addr_fast[3]\, Kt_addr_fast(2) => 
        \Kt_addr_fast[2]\, sha256_controller_0_bytes_o(1) => 
        sha256_controller_0_bytes_o(1), W_out_2_0(5) => 
        \W_out_2_0[5]\, W_out_i_0(2) => \W_out_i_0[2]\, 
        W_out_i_0(1) => \W_out_i_0[1]\, W_out_i_0(0) => 
        \W_out_i_0[0]\, W_out_i_i_1_1(31) => \W_out_i_i_1_1[31]\, 
        W_out_2_0_1(7) => \W_out_2_0_1[7]\, W_out_i_i_1(31) => 
        \W_out_i_i_1[31]\, W_out_2_0_a4_1_0_RNIFI1DA(23) => 
        \W_out_2_0_a4_1_0_RNIFI1DA[23]\, 
        W_out_2_0_a4_1_0_RNI32U7B(23) => 
        \W_out_2_0_a4_1_0_RNI32U7B[23]\, msg_bitlen(63) => 
        \msg_bitlen[63]\, msg_bitlen(62) => \msg_bitlen[62]\, 
        msg_bitlen(61) => \msg_bitlen[61]\, msg_bitlen(60) => 
        \msg_bitlen[60]\, msg_bitlen(59) => \msg_bitlen[59]\, 
        msg_bitlen(58) => \msg_bitlen[58]\, msg_bitlen(57) => 
        \msg_bitlen[57]\, msg_bitlen(56) => \msg_bitlen[56]\, 
        msg_bitlen(55) => \msg_bitlen[55]\, msg_bitlen(54) => 
        \msg_bitlen[54]\, msg_bitlen(53) => \msg_bitlen[53]\, 
        msg_bitlen(52) => \msg_bitlen[52]\, msg_bitlen(51) => 
        \msg_bitlen[51]\, msg_bitlen(50) => \msg_bitlen[50]\, 
        msg_bitlen(49) => \msg_bitlen[49]\, msg_bitlen(48) => 
        \msg_bitlen[48]\, msg_bitlen(47) => \msg_bitlen[47]\, 
        msg_bitlen(46) => \msg_bitlen[46]\, msg_bitlen(45) => 
        \msg_bitlen[45]\, msg_bitlen(44) => \msg_bitlen[44]\, 
        msg_bitlen(43) => \msg_bitlen[43]\, msg_bitlen(42) => 
        \msg_bitlen[42]\, msg_bitlen(41) => \msg_bitlen[41]\, 
        msg_bitlen(40) => \msg_bitlen[40]\, msg_bitlen(39) => 
        \msg_bitlen[39]\, msg_bitlen(38) => \msg_bitlen[38]\, 
        msg_bitlen(37) => \msg_bitlen[37]\, msg_bitlen(36) => 
        \msg_bitlen[36]\, msg_bitlen(35) => \msg_bitlen[35]\, 
        msg_bitlen(34) => \msg_bitlen[34]\, msg_bitlen(33) => 
        \msg_bitlen[33]\, msg_bitlen(32) => \msg_bitlen[32]\, 
        msg_bitlen(31) => \msg_bitlen[31]\, msg_bitlen(30) => 
        \msg_bitlen[30]\, msg_bitlen(29) => \msg_bitlen[29]\, 
        msg_bitlen(28) => \msg_bitlen[28]\, msg_bitlen(27) => 
        \msg_bitlen[27]\, msg_bitlen(26) => \msg_bitlen[26]\, 
        msg_bitlen(25) => \msg_bitlen[25]\, msg_bitlen(24) => 
        \msg_bitlen[24]\, msg_bitlen(23) => \msg_bitlen[23]\, 
        msg_bitlen(22) => \msg_bitlen[22]\, msg_bitlen(21) => 
        \msg_bitlen[21]\, msg_bitlen(20) => \msg_bitlen[20]\, 
        msg_bitlen(19) => \msg_bitlen[19]\, msg_bitlen(18) => 
        \msg_bitlen[18]\, msg_bitlen(17) => \msg_bitlen[17]\, 
        msg_bitlen(16) => \msg_bitlen[16]\, msg_bitlen(15) => 
        \msg_bitlen[15]\, msg_bitlen(14) => \msg_bitlen[14]\, 
        msg_bitlen(13) => \msg_bitlen[13]\, msg_bitlen(12) => 
        \msg_bitlen[12]\, msg_bitlen(11) => \msg_bitlen[11]\, 
        msg_bitlen(10) => \msg_bitlen[10]\, msg_bitlen(9) => 
        \msg_bitlen[9]\, msg_bitlen(8) => \msg_bitlen[8]\, 
        msg_bitlen(7) => \msg_bitlen[7]\, msg_bitlen(6) => 
        \msg_bitlen[6]\, msg_bitlen(5) => \msg_bitlen[5]\, 
        msg_bitlen(4) => \msg_bitlen[4]\, msg_bitlen(3) => 
        \msg_bitlen[3]\, state_2 => state_2, state_0 => state_0, 
        state_3 => state_3, W_out_2_0_0_20 => \W_out_2_0_0[23]\, 
        W_out_2_0_0_12 => \W_out_2_0_0[15]\, W_out_2_0_0_4 => 
        \W_out_2_0_0[7]\, W_out_2_0_0_1 => \W_out_2_0_0[4]\, 
        W_out_2_0_0_3 => \W_out_2_0_0[6]\, W_out_2_0_0_0 => 
        \W_out_2_0_0[3]\, W_out_2_i_0_22 => \W_out_2_i_0[30]\, 
        W_out_2_i_0_17 => \W_out_2_i_0[25]\, W_out_2_i_0_21 => 
        \W_out_2_i_0[29]\, W_out_2_i_0_20 => \W_out_2_i_0[28]\, 
        W_out_2_i_0_16 => \W_out_2_i_0[24]\, W_out_2_i_0_18 => 
        \W_out_2_i_0[26]\, W_out_2_i_0_19 => \W_out_2_i_0[27]\, 
        W_out_2_i_2_0 => \W_out_2_i_2[8]\, W_out_2_i_2_5 => 
        \W_out_2_i_2[13]\, W_out_2_i_2_6 => \W_out_2_i_2[14]\, 
        W_out_2_i_1_1 => \W_out_2_i_1[9]\, W_out_2_i_1_0 => 
        \W_out_2_i_1[8]\, W_out_2_i_1_22 => \W_out_2_i_1[30]\, 
        W_out_2_i_1_17 => \W_out_2_i_1[25]\, W_out_2_i_1_21 => 
        \W_out_2_i_1[29]\, W_out_2_i_1_20 => \W_out_2_i_1[28]\, 
        W_out_2_i_1_16 => \W_out_2_i_1[24]\, W_out_2_i_1_18 => 
        \W_out_2_i_1[26]\, W_out_2_i_1_19 => \W_out_2_i_1[27]\, 
        W_out_2_i_1_13 => \W_out_2_i_1[21]\, W_out_2_i_1_10 => 
        \W_out_2_i_1[18]\, W_out_2_i_1_12 => \W_out_2_i_1[20]\, 
        W_out_2_i_1_14 => \W_out_2_i_1[22]\, W_out_2_i_1_9 => 
        \W_out_2_i_1[17]\, W_out_2_i_1_11 => \W_out_2_i_1[19]\, 
        W_out_2_i_1_8 => \W_out_2_i_1[16]\, W_out_2_i_1_2 => 
        \W_out_2_i_1[10]\, W_out_2_i_1_4 => \W_out_2_i_1[12]\, 
        W_out_2_i_1_3 => \W_out_2_i_1[11]\, N_1696 => N_1696, 
        SHA256_Module_0_di_req_o => \SHA256_Module_0_di_req_o\, 
        N_1400 => N_1400, N_1624 => N_1624, N_920 => N_920, 
        N_1144 => N_1144, N_1399 => N_1399, N_1623 => N_1623, 
        N_919 => N_919, N_1143 => N_1143, N_1401 => N_1401, 
        N_1625 => N_1625, N_921 => N_921, N_1145 => N_1145, 
        one_insert => one_insert, N_388 => N_388, W_m4_e_2 => 
        W_m4_e_2, Kt_addr_1_rep1 => Kt_addr_1_rep1, N_102 => 
        N_102, N_105 => N_105, ren_pos => ren_pos, 
        sha256_controller_0_end_o => sha256_controller_0_end_o, 
        Kt_addr_0_rep2 => Kt_addr_0_rep2, sha_last_blk_reg => 
        sha_last_blk_reg, sha_last_blk_next_0_o2_0 => 
        sha_last_blk_next_0_o2_0, N_387 => N_387, N_98 => N_98, 
        N_111 => N_111, N_1694 => N_1694, N_1692 => N_1692, N_349
         => N_349, N_1693 => N_1693, N_251 => N_251, N_1691 => 
        N_1691, N_248 => N_248, N_1690 => N_1690, N_245 => N_245, 
        N_89 => N_89, N_1695 => N_1695, N_1708 => N_1708, N_1709
         => N_1709, N_1707 => N_1707, N_1706 => N_1706, N_1705
         => N_1705, N_1704 => N_1704, N_1703 => N_1703, N_1700
         => N_1700, N_1701 => N_1701, N_1697 => N_1697, N_1699
         => N_1699, N_1698 => N_1698, N_1717 => N_1717, N_1712
         => N_1712, N_1716 => N_1716, N_1715 => N_1715, N_1711
         => N_1711, N_1713 => N_1713, N_1714 => N_1714, N_1718
         => N_1718, N_1702 => N_1702, N_1710 => N_1710, N_263 => 
        N_263, N_301 => N_301, N_304 => N_304, N_298 => N_298, 
        N_295 => N_295, N_292 => N_292, N_289 => N_289, N_286 => 
        N_286, N_278 => N_278, N_275 => N_275, N_272 => N_272, 
        N_268 => N_268, N_265 => N_265);
    
    Inst_sha256_msg_sch : sha256_msg_sch
      port map(Wt_data(31) => \Wt_data[31]\, Wt_data(30) => 
        \Wt_data[30]\, Wt_data(29) => \Wt_data[29]\, Wt_data(28)
         => \Wt_data[28]\, Wt_data(27) => \Wt_data[27]\, 
        Wt_data(26) => \Wt_data[26]\, Wt_data(25) => 
        \Wt_data[25]\, Wt_data(24) => \Wt_data[24]\, Wt_data(23)
         => \Wt_data[23]\, Wt_data(22) => \Wt_data[22]\, 
        Wt_data(21) => \Wt_data[21]\, Wt_data(20) => 
        \Wt_data[20]\, Wt_data(19) => \Wt_data[19]\, Wt_data(18)
         => \Wt_data[18]\, Wt_data(17) => \Wt_data[17]\, 
        Wt_data(16) => \Wt_data[16]\, Wt_data(15) => 
        \Wt_data[15]\, Wt_data(14) => \Wt_data[14]\, Wt_data(13)
         => \Wt_data[13]\, Wt_data(12) => \Wt_data[12]\, 
        Wt_data(11) => \Wt_data[11]\, Wt_data(10) => 
        \Wt_data[10]\, Wt_data(9) => \Wt_data[9]\, Wt_data(8) => 
        \Wt_data[8]\, Wt_data(7) => \Wt_data[7]\, Wt_data(6) => 
        \Wt_data[6]\, Wt_data(5) => \Wt_data[5]\, Wt_data(4) => 
        \Wt_data[4]\, Wt_data(3) => \Wt_data[3]\, Wt_data(2) => 
        \Wt_data[2]\, Wt_data(1) => \Wt_data[1]\, Wt_data(0) => 
        \Wt_data[0]\, W_out_2_0(5) => \W_out_2_0[5]\, 
        W_out_i_0(2) => \W_out_i_0[2]\, W_out_i_0(1) => 
        \W_out_i_0[1]\, W_out_i_0(0) => \W_out_i_0[0]\, 
        W_out_i_i_1_1(31) => \W_out_i_i_1_1[31]\, W_out_i_i_1(31)
         => \W_out_i_i_1[31]\, W_out_2_i_0(30) => 
        \W_out_2_i_0[30]\, W_out_2_i_0(29) => \W_out_2_i_0[29]\, 
        W_out_2_i_0(28) => \W_out_2_i_0[28]\, W_out_2_i_0(27) => 
        \W_out_2_i_0[27]\, W_out_2_i_0(26) => \W_out_2_i_0[26]\, 
        W_out_2_i_0(25) => \W_out_2_i_0[25]\, W_out_2_i_0(24) => 
        \W_out_2_i_0[24]\, W_out_2_0_a4_1_0_RNI32U7B(23) => 
        \W_out_2_0_a4_1_0_RNI32U7B[23]\, 
        W_out_2_0_a4_1_0_RNIFI1DA(23) => 
        \W_out_2_0_a4_1_0_RNIFI1DA[23]\, W_out_2_0_1(7) => 
        \W_out_2_0_1[7]\, W_out_2_0_0_3 => \W_out_2_0_0[6]\, 
        W_out_2_0_0_1 => \W_out_2_0_0[4]\, W_out_2_0_0_0 => 
        \W_out_2_0_0[3]\, W_out_2_0_0_20 => \W_out_2_0_0[23]\, 
        W_out_2_0_0_12 => \W_out_2_0_0[15]\, W_out_2_0_0_4 => 
        \W_out_2_0_0[7]\, W_out_2_i_2_0 => \W_out_2_i_2[8]\, 
        W_out_2_i_2_6 => \W_out_2_i_2[14]\, W_out_2_i_2_5 => 
        \W_out_2_i_2[13]\, W_out_2_i_1_22 => \W_out_2_i_1[30]\, 
        W_out_2_i_1_21 => \W_out_2_i_1[29]\, W_out_2_i_1_20 => 
        \W_out_2_i_1[28]\, W_out_2_i_1_19 => \W_out_2_i_1[27]\, 
        W_out_2_i_1_18 => \W_out_2_i_1[26]\, W_out_2_i_1_17 => 
        \W_out_2_i_1[25]\, W_out_2_i_1_16 => \W_out_2_i_1[24]\, 
        W_out_2_i_1_0 => \W_out_2_i_1[8]\, W_out_2_i_1_14 => 
        \W_out_2_i_1[22]\, W_out_2_i_1_13 => \W_out_2_i_1[21]\, 
        W_out_2_i_1_12 => \W_out_2_i_1[20]\, W_out_2_i_1_11 => 
        \W_out_2_i_1[19]\, W_out_2_i_1_10 => \W_out_2_i_1[18]\, 
        W_out_2_i_1_9 => \W_out_2_i_1[17]\, W_out_2_i_1_8 => 
        \W_out_2_i_1[16]\, W_out_2_i_1_4 => \W_out_2_i_1[12]\, 
        W_out_2_i_1_3 => \W_out_2_i_1[11]\, W_out_2_i_1_2 => 
        \W_out_2_i_1[10]\, W_out_2_i_1_1 => \W_out_2_i_1[9]\, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, N_244_i_0 => N_244_i_0, 
        next_r0_0_cry_0_Y => next_r0_0_cry_0_Y, N_251 => N_251, 
        ld_i_i_3 => ld_i_i_3, N_349 => N_349, N_248 => N_248, 
        N_245 => N_245, N_98 => N_98, N_304 => N_304, N_301 => 
        N_301, N_298 => N_298, N_295 => N_295, N_292 => N_292, 
        N_289 => N_289, N_286 => N_286, N_278 => N_278, N_275 => 
        N_275, N_272 => N_272, N_268 => N_268, N_265 => N_265, 
        N_263 => N_263);
    
    Inst_sha256_kt_rom : sha256_kt_rom
      port map(hash_control_st_reg_ns_i_0_a2_0(4) => 
        \hash_control_st_reg_ns_i_0_a2_0[4]\, 
        hash_control_st_reg_ns_i_0_a2_2(4) => 
        \hash_control_st_reg_ns_i_0_a2_2[4]\, Kt_addr(5) => 
        \Kt_addr[5]\, Kt_addr(4) => \Kt_addr[4]\, Kt_addr(3) => 
        \Kt_addr[3]\, Kt_addr(2) => \Kt_addr[2]\, Kt_addr(1) => 
        \Kt_addr[1]\, Kt_addr(0) => \Kt_addr[0]\, Kt_addr_fast(4)
         => \Kt_addr_fast[4]\, Kt_addr_fast(3) => 
        \Kt_addr_fast[3]\, Kt_addr_fast(2) => \Kt_addr_fast[2]\, 
        Kt_addr_fast(1) => \Kt_addr_fast[1]\, Kt_addr_fast(0) => 
        \Kt_addr_fast[0]\, Kt_data_0 => \Kt_data[0]\, Kt_data_24
         => \Kt_data[24]\, Kt_data_15 => \Kt_data[15]\, m10_bm
         => m10_bm, m20_1 => m20_1, m10_am => m10_am, 
        Kt_addr_5_rep1 => Kt_addr_5_rep1, Kt_addr_3_rep2 => 
        Kt_addr_3_rep2, Kt_addr_3_rep1 => Kt_addr_3_rep1, m62_am
         => m62_am, Kt_addr_0_rep1 => Kt_addr_0_rep1, m104_bm => 
        m104_bm, Kt_addr_2_rep1 => Kt_addr_2_rep1, Kt_addr_0_rep2
         => Kt_addr_0_rep2, m49_am => m49_am, Kt_addr_1_rep1 => 
        Kt_addr_1_rep1, m49_bm => m49_bm, m137_am => m137_am, 
        m137_bm => m137_bm, Kt_addr_2_rep2 => Kt_addr_2_rep2, 
        Kt_addr_1_rep2 => Kt_addr_1_rep2, Kt_addr_4_rep2 => 
        Kt_addr_4_rep2, m215_am => m215_am, Kt_addr_4_rep1 => 
        Kt_addr_4_rep1, m215_bm => m215_bm, m250_am => m250_am, 
        m250_bm => m250_bm, m207_1_1 => m207_1_1, m207_1_0 => 
        m207_1_0, m95_1_1 => m95_1_1, m95_1_0 => m95_1_0, 
        m197_1_1 => m197_1_1, m197_1_0 => m197_1_0, m316 => m316, 
        m34 => m34, m157 => m157, m325 => m325, m168_1_1 => 
        m168_1_1, m168_1_0 => m168_1_0, m230 => m230, m296 => 
        m296, m254 => m254, m114 => m114, m304 => m304, m73_0 => 
        m73, pad_one_reg_0_0_a2_0 => pad_one_reg_0_0_a2_0, m239
         => m239, m219 => m219, m285 => m285, m177 => m177, m124
         => m124, m289 => m289, m78 => m78, m141 => m141, 
        i3_mux_1 => i3_mux_1, m67_ns => m67_ns, m83_ns => m83_ns, 
        m110_ns => m110_ns, m119_ns => m119_ns, m144_ns => 
        m144_ns, m172_ns => m172_ns, m222_ns => m222_ns, m226_ns
         => m226_ns, m235_ns => m235_ns, m258_ns => m258_ns, 
        m276_ns => m276_ns, m281_ns => m281_ns, m292_ns => 
        m292_ns, m300_ns => m300_ns, m273 => m273, m104_am => 
        m104_am, m62_bm => m62_bm);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity limiter_1cycle_0 is

    port( prev_sig                     : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK : in    std_logic;
          first_block                  : in    std_logic
        );

end limiter_1cycle_0;

architecture DEF_ARCH of limiter_1cycle_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \prev_sig\ : SLE
      port map(D => first_block, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => prev_sig);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity limiter_1cycle_1 is

    port( prev_sig                       : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic;
          SHA256_Module_0_data_out_ready : in    std_logic
        );

end limiter_1cycle_1;

architecture DEF_ARCH of limiter_1cycle_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \prev_sig\ : SLE
      port map(D => SHA256_Module_0_data_out_ready, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => prev_sig);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_17x32 is

    port( AHB_slave_dummy_0_mem_wdata     : in    std_logic_vector(31 downto 0);
          sha256_controller_0_read_addr_0 : in    std_logic_vector(3 downto 0);
          waddr_in_net_0                  : in    std_logic_vector(4 downto 0);
          raddr_pos_3                     : out   std_logic;
          raddr_pos_2                     : out   std_logic;
          SHA256_Module_0_data_out_ready  : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK    : in    std_logic;
          sha256_system_sb_0_GPIO_9_M2F   : in    std_logic;
          SHA256_Module_0_data_available  : out   std_logic;
          ren_pos                         : out   std_logic;
          last_block                      : out   std_logic;
          first_block                     : out   std_logic;
          N_1717                          : out   std_logic;
          N_1716                          : out   std_logic;
          N_1711                          : out   std_logic;
          N_1710                          : out   std_logic;
          N_1708                          : out   std_logic;
          N_1705                          : out   std_logic;
          N_1704                          : out   std_logic;
          N_1701                          : out   std_logic;
          N_1690                          : out   std_logic;
          N_1691                          : out   std_logic;
          N_1707                          : out   std_logic;
          N_1703                          : out   std_logic;
          N_1715                          : out   std_logic;
          N_1700                          : out   std_logic;
          N_1714                          : out   std_logic;
          N_1697                          : out   std_logic;
          N_1693                          : out   std_logic;
          N_1706                          : out   std_logic;
          N_1696                          : out   std_logic;
          N_1709                          : out   std_logic;
          N_1698                          : out   std_logic;
          N_1699                          : out   std_logic;
          N_1694                          : out   std_logic;
          N_1702                          : out   std_logic;
          N_1712                          : out   std_logic;
          N_1695                          : out   std_logic;
          N_1692                          : out   std_logic;
          N_1718                          : out   std_logic;
          N_1713                          : out   std_logic;
          N_1144                          : out   std_logic;
          N_921                           : out   std_logic;
          N_1401                          : out   std_logic;
          N_1145                          : out   std_logic;
          N_919                           : out   std_logic;
          N_1400                          : out   std_logic;
          N_1623                          : out   std_logic;
          N_920                           : out   std_logic;
          N_1143                          : out   std_logic;
          N_1624                          : out   std_logic;
          N_1625                          : out   std_logic;
          N_1399                          : out   std_logic;
          sha256_system_sb_0_GPIO_1_M2F   : in    std_logic;
          AHB_slave_dummy_0_write_en      : in    std_logic
        );

end reg_17x32;

architecture DEF_ARCH of reg_17x32 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \SHA256_Module_0_data_out_ready\, VCC_net_1, 
        \data_out_ready_1\, GND_net_1, 
        \SHA256_Module_0_data_available\, N_12_0_i_0, 
        data_out_ready_0_sqmuxa, \line8_or[0]_net_1\, line8_0_62, 
        \line7[63]_net_1\, \line7_or[32]_net_1\, 
        \line7[62]_net_1\, \line7[61]_net_1\, \line7[60]_net_1\, 
        \line7[59]_net_1\, \line7[58]_net_1\, \line7[57]_net_1\, 
        \line7[56]_net_1\, \line7[55]_net_1\, \line7[54]_net_1\, 
        \line7[53]_net_1\, \line7[52]_net_1\, \line7[51]_net_1\, 
        \line7[50]_net_1\, \line7[49]_net_1\, \line7[48]_net_1\, 
        \line7[47]_net_1\, \line7[46]_net_1\, \line7[45]_net_1\, 
        \line7[44]_net_1\, \line7[43]_net_1\, \line7[42]_net_1\, 
        \line7[41]_net_1\, \line7[40]_net_1\, \line7[39]_net_1\, 
        \line7[38]_net_1\, \line7[37]_net_1\, \line7[36]_net_1\, 
        \line7[35]_net_1\, \line7[34]_net_1\, \line7[33]_net_1\, 
        \line7[32]_net_1\, line7_0, \line7[31]_net_1\, 
        \line7_or[0]_net_1\, \line7[30]_net_1\, \line7[29]_net_1\, 
        \line7[28]_net_1\, \line7[27]_net_1\, \line7[26]_net_1\, 
        \line7[25]_net_1\, \line7[24]_net_1\, \line7[23]_net_1\, 
        \line7[22]_net_1\, \line7[21]_net_1\, \line7[20]_net_1\, 
        \line7[19]_net_1\, \line7[18]_net_1\, \line7[17]_net_1\, 
        \line7[16]_net_1\, \line7[15]_net_1\, \line7[14]_net_1\, 
        \line7[13]_net_1\, \line7[12]_net_1\, \line7[11]_net_1\, 
        \line7[10]_net_1\, \line7[9]_net_1\, \line7[8]_net_1\, 
        \line7[7]_net_1\, \line7[6]_net_1\, \line7[5]_net_1\, 
        \line7[4]_net_1\, \line7[3]_net_1\, \line7[2]_net_1\, 
        \line7[1]_net_1\, \line7[0]_net_1\, line7_0_62, 
        \line6[63]_net_1\, \line6_or[32]_net_1\, 
        \line6[62]_net_1\, \line6[61]_net_1\, \line6[60]_net_1\, 
        \line6[59]_net_1\, \line6[58]_net_1\, \line6[57]_net_1\, 
        \line6[56]_net_1\, \line6[55]_net_1\, \line6[54]_net_1\, 
        \line6[53]_net_1\, \line6[52]_net_1\, \line6[51]_net_1\, 
        \line6[50]_net_1\, \line6[49]_net_1\, \line6[48]_net_1\, 
        \line6[47]_net_1\, \line6[46]_net_1\, \line6[45]_net_1\, 
        \line6[44]_net_1\, \line6[43]_net_1\, \line6[42]_net_1\, 
        \line6[41]_net_1\, \line6[40]_net_1\, \line6[39]_net_1\, 
        \line6[38]_net_1\, \line6[37]_net_1\, \line6[36]_net_1\, 
        \line6[35]_net_1\, \line6[34]_net_1\, \line6[33]_net_1\, 
        \line6[32]_net_1\, line6_0, \line6[31]_net_1\, 
        \line6_or[0]_net_1\, \line6[30]_net_1\, \line6[29]_net_1\, 
        \line6[28]_net_1\, \line6[27]_net_1\, \line6[26]_net_1\, 
        \line6[25]_net_1\, \line6[24]_net_1\, \line6[23]_net_1\, 
        \line6[22]_net_1\, \line6[21]_net_1\, \line6[20]_net_1\, 
        \line6[19]_net_1\, \line6[18]_net_1\, \line6[17]_net_1\, 
        \line6[16]_net_1\, \line6[15]_net_1\, \line6[14]_net_1\, 
        \line6[13]_net_1\, \line6[12]_net_1\, \line6[11]_net_1\, 
        \line6[10]_net_1\, \line6[9]_net_1\, \line6[8]_net_1\, 
        \line6[7]_net_1\, \line6[6]_net_1\, \line6[5]_net_1\, 
        \line6[4]_net_1\, \line6[3]_net_1\, \line6[2]_net_1\, 
        \line6[1]_net_1\, \line6[0]_net_1\, line6_0_62, 
        \line5[63]_net_1\, \line5_or[32]_net_1\, 
        \line5[62]_net_1\, \line5[61]_net_1\, \line5[60]_net_1\, 
        \line5[59]_net_1\, \line5[58]_net_1\, \line5[57]_net_1\, 
        \line5[56]_net_1\, \line5[55]_net_1\, \line5[54]_net_1\, 
        \line5[53]_net_1\, \line5[52]_net_1\, \line5[51]_net_1\, 
        \line5[50]_net_1\, \line5[49]_net_1\, \line5[48]_net_1\, 
        \line5[47]_net_1\, \line5[46]_net_1\, \line5[45]_net_1\, 
        \line5[44]_net_1\, \line5[43]_net_1\, \line5[42]_net_1\, 
        \line5[41]_net_1\, \line5[40]_net_1\, \line5[39]_net_1\, 
        \line5[38]_net_1\, \line5[37]_net_1\, \line5[36]_net_1\, 
        \line5[35]_net_1\, \line5[34]_net_1\, \line5[33]_net_1\, 
        \line5[32]_net_1\, line5_0, \line5[31]_net_1\, 
        \line5_or[0]_net_1\, \line5[30]_net_1\, \line5[29]_net_1\, 
        \line5[28]_net_1\, \line5[27]_net_1\, \line5[26]_net_1\, 
        \line5[25]_net_1\, \line5[24]_net_1\, \line5[23]_net_1\, 
        \line5[22]_net_1\, \line5[21]_net_1\, \line5[20]_net_1\, 
        \line5[19]_net_1\, \line5[18]_net_1\, \line5[17]_net_1\, 
        \line5[16]_net_1\, \line5[15]_net_1\, \line5[14]_net_1\, 
        \line5[13]_net_1\, \line5[12]_net_1\, \line5[11]_net_1\, 
        \line5[10]_net_1\, \line5[9]_net_1\, \line5[8]_net_1\, 
        \line5[7]_net_1\, \line5[6]_net_1\, \line5[5]_net_1\, 
        \line5[4]_net_1\, \line5[3]_net_1\, \line5[2]_net_1\, 
        \line5[1]_net_1\, \line5[0]_net_1\, line5_0_62, 
        \line4[63]_net_1\, \line4_or[32]_net_1\, 
        \line4[62]_net_1\, \line4[61]_net_1\, \line4[60]_net_1\, 
        \line4[59]_net_1\, \line4[58]_net_1\, \line4[57]_net_1\, 
        \line4[56]_net_1\, \line4[55]_net_1\, \line4[54]_net_1\, 
        \line4[53]_net_1\, \line4[52]_net_1\, \line4[51]_net_1\, 
        \line4[50]_net_1\, \line4[49]_net_1\, \line4[48]_net_1\, 
        \line4[47]_net_1\, \line4[46]_net_1\, \line4[45]_net_1\, 
        \line4[44]_net_1\, \line4[43]_net_1\, \line4[42]_net_1\, 
        \line4[41]_net_1\, \line4[40]_net_1\, \line4[39]_net_1\, 
        \line4[38]_net_1\, \line4[37]_net_1\, \line4[36]_net_1\, 
        \line4[35]_net_1\, \line4[34]_net_1\, \line4[33]_net_1\, 
        \line4[32]_net_1\, line4_0, \line4[31]_net_1\, 
        \line4_or[0]_net_1\, \line4[30]_net_1\, \line4[29]_net_1\, 
        \line4[28]_net_1\, \line4[27]_net_1\, \line4[26]_net_1\, 
        \line4[25]_net_1\, \line4[24]_net_1\, \line4[23]_net_1\, 
        \line4[22]_net_1\, \line4[21]_net_1\, \line4[20]_net_1\, 
        \line4[19]_net_1\, \line4[18]_net_1\, \line4[17]_net_1\, 
        \line4[16]_net_1\, \line4[15]_net_1\, \line4[14]_net_1\, 
        \line4[13]_net_1\, \line4[12]_net_1\, \line4[11]_net_1\, 
        \line4[10]_net_1\, \line4[9]_net_1\, \line4[8]_net_1\, 
        \line4[7]_net_1\, \line4[6]_net_1\, \line4[5]_net_1\, 
        \line4[4]_net_1\, \line4[3]_net_1\, \line4[2]_net_1\, 
        \line4[1]_net_1\, \line4[0]_net_1\, line4_0_62, 
        \line3[63]_net_1\, \line3_or[32]_net_1\, 
        \line3[62]_net_1\, \line3[61]_net_1\, \line3[60]_net_1\, 
        \line3[59]_net_1\, \line3[58]_net_1\, \line3[57]_net_1\, 
        \line3[56]_net_1\, \line3[55]_net_1\, \line3[54]_net_1\, 
        \line3[53]_net_1\, \line3[52]_net_1\, \line3[51]_net_1\, 
        \line3[50]_net_1\, \line3[49]_net_1\, \line3[48]_net_1\, 
        \line3[47]_net_1\, \line3[46]_net_1\, \line3[45]_net_1\, 
        \line3[44]_net_1\, \line3[43]_net_1\, \line3[42]_net_1\, 
        \line3[41]_net_1\, \line3[40]_net_1\, \line3[39]_net_1\, 
        \line3[38]_net_1\, \line3[37]_net_1\, \line3[36]_net_1\, 
        \line3[35]_net_1\, \line3[34]_net_1\, \line3[33]_net_1\, 
        \line3[32]_net_1\, line3_0, \line3[31]_net_1\, 
        \line3_or[0]_net_1\, \line3[30]_net_1\, \line3[29]_net_1\, 
        \line3[28]_net_1\, \line3[27]_net_1\, \line3[26]_net_1\, 
        \line3[25]_net_1\, \line3[24]_net_1\, \line3[23]_net_1\, 
        \line3[22]_net_1\, \line3[21]_net_1\, \line3[20]_net_1\, 
        \line3[19]_net_1\, \line3[18]_net_1\, \line3[17]_net_1\, 
        \line3[16]_net_1\, \line3[15]_net_1\, \line3[14]_net_1\, 
        \line3[13]_net_1\, \line3[12]_net_1\, \line3[11]_net_1\, 
        \line3[10]_net_1\, \line3[9]_net_1\, \line3[8]_net_1\, 
        \line3[7]_net_1\, \line3[6]_net_1\, \line3[5]_net_1\, 
        \line3[4]_net_1\, \line3[3]_net_1\, \line3[2]_net_1\, 
        \line3[1]_net_1\, \line3[0]_net_1\, line3_0_62, 
        \line2[63]_net_1\, \line2_or[32]_net_1\, 
        \line2[62]_net_1\, \line2[61]_net_1\, \line2[60]_net_1\, 
        \line2[59]_net_1\, \line2[58]_net_1\, \line2[57]_net_1\, 
        \line2[56]_net_1\, \line2[55]_net_1\, \line2[54]_net_1\, 
        \line2[53]_net_1\, \line2[52]_net_1\, \line2[51]_net_1\, 
        \line2[50]_net_1\, \line2[49]_net_1\, \line2[48]_net_1\, 
        \line2[47]_net_1\, \line2[46]_net_1\, \line2[45]_net_1\, 
        \line2[44]_net_1\, \line2[43]_net_1\, \line2[42]_net_1\, 
        \line2[41]_net_1\, \line2[40]_net_1\, \line2[39]_net_1\, 
        \line2[38]_net_1\, \line2[37]_net_1\, \line2[36]_net_1\, 
        \line2[35]_net_1\, \line2[34]_net_1\, \line2[33]_net_1\, 
        \line2[32]_net_1\, line2_0, \line2[31]_net_1\, 
        \line2_or[0]_net_1\, \line2[30]_net_1\, \line2[29]_net_1\, 
        \line2[28]_net_1\, \line2[27]_net_1\, \line2[26]_net_1\, 
        \line2[25]_net_1\, \line2[24]_net_1\, \line2[23]_net_1\, 
        \line2[22]_net_1\, \line2[21]_net_1\, \line2[20]_net_1\, 
        \line2[19]_net_1\, \line2[18]_net_1\, \line2[17]_net_1\, 
        \line2[16]_net_1\, \line2[15]_net_1\, \line2[14]_net_1\, 
        \line2[13]_net_1\, \line2[12]_net_1\, \line2[11]_net_1\, 
        \line2[10]_net_1\, \line2[9]_net_1\, \line2[8]_net_1\, 
        \line2[7]_net_1\, \line2[6]_net_1\, \line2[5]_net_1\, 
        \line2[4]_net_1\, \line2[3]_net_1\, \line2[2]_net_1\, 
        \line2[1]_net_1\, \line2[0]_net_1\, line2_0_62, 
        \line1[63]_net_1\, \line1_or[32]_net_1\, 
        \line1[62]_net_1\, \line1[61]_net_1\, \line1[60]_net_1\, 
        \line1[59]_net_1\, \line1[58]_net_1\, \line1[57]_net_1\, 
        \line1[56]_net_1\, \line1[55]_net_1\, \line1[54]_net_1\, 
        \line1[53]_net_1\, \line1[52]_net_1\, \line1[51]_net_1\, 
        \line1[50]_net_1\, \line1[49]_net_1\, \line1[48]_net_1\, 
        \line1[47]_net_1\, \line1[46]_net_1\, \line1[45]_net_1\, 
        \line1[44]_net_1\, \line1[43]_net_1\, \line1[42]_net_1\, 
        \line1[41]_net_1\, \line1[40]_net_1\, \line1[39]_net_1\, 
        \line1[38]_net_1\, \line1[37]_net_1\, \line1[36]_net_1\, 
        \line1[35]_net_1\, \line1[34]_net_1\, \line1[33]_net_1\, 
        \line1[32]_net_1\, line1_0, \line1[31]_net_1\, 
        \line1_or[0]_net_1\, \line1[30]_net_1\, \line1[29]_net_1\, 
        \line1[28]_net_1\, \line1[27]_net_1\, \line1[26]_net_1\, 
        \line1[25]_net_1\, \line1[24]_net_1\, \line1[23]_net_1\, 
        \line1[22]_net_1\, \line1[21]_net_1\, \line1[20]_net_1\, 
        \line1[19]_net_1\, \line1[18]_net_1\, \line1[17]_net_1\, 
        \line1[16]_net_1\, \line1[15]_net_1\, \line1[14]_net_1\, 
        \line1[13]_net_1\, \line1[12]_net_1\, \line1[11]_net_1\, 
        \line1[10]_net_1\, \line1[9]_net_1\, \line1[8]_net_1\, 
        \line1[7]_net_1\, \line1[6]_net_1\, \line1[5]_net_1\, 
        \line1[4]_net_1\, \line1[3]_net_1\, \line1[2]_net_1\, 
        \line1[1]_net_1\, \line1[0]_net_1\, line1_0_62, 
        \line0[63]_net_1\, \line0_or[32]_net_1\, 
        \line0[62]_net_1\, \line0[61]_net_1\, \line0[60]_net_1\, 
        \line0[59]_net_1\, \line0[58]_net_1\, \line0[57]_net_1\, 
        \line0[56]_net_1\, \line0[55]_net_1\, \line0[54]_net_1\, 
        \line0[53]_net_1\, \line0[52]_net_1\, \line0[51]_net_1\, 
        \line0[50]_net_1\, \line0[49]_net_1\, \line0[48]_net_1\, 
        \line0[47]_net_1\, \line0[46]_net_1\, \line0[45]_net_1\, 
        \line0[44]_net_1\, \line0[43]_net_1\, \line0[42]_net_1\, 
        \line0[41]_net_1\, \line0[40]_net_1\, \line0[39]_net_1\, 
        \line0[38]_net_1\, \line0[37]_net_1\, \line0[36]_net_1\, 
        \line0[35]_net_1\, \line0[34]_net_1\, \line0[33]_net_1\, 
        \line0[32]_net_1\, line0_0, \line0[31]_net_1\, 
        \line0_or[0]_net_1\, \line0[30]_net_1\, \line0[29]_net_1\, 
        \line0[28]_net_1\, \line0[27]_net_1\, \line0[26]_net_1\, 
        \line0[25]_net_1\, \line0[24]_net_1\, \line0[23]_net_1\, 
        \line0[22]_net_1\, \line0[21]_net_1\, \line0[20]_net_1\, 
        \line0[19]_net_1\, \line0[18]_net_1\, \line0[17]_net_1\, 
        \line0[16]_net_1\, \line0[15]_net_1\, \line0[14]_net_1\, 
        \line0[13]_net_1\, \line0[12]_net_1\, \line0[11]_net_1\, 
        \line0[10]_net_1\, \line0[9]_net_1\, \line0[8]_net_1\, 
        \line0[7]_net_1\, \line0[6]_net_1\, \line0[5]_net_1\, 
        \line0[4]_net_1\, \line0[3]_net_1\, \line0[2]_net_1\, 
        \line0[1]_net_1\, \line0[0]_net_1\, line0_0_62, 
        \raddr_pos_3\, N_3_0, \raddr_pos_2\, \raddr_pos[1]_net_1\, 
        \raddr_pos[0]_net_1\, \raddr_pos_fast[0]_net_1\, 
        \raddr_pos_0_rep1\, \raddr_pos_0_rep2\, 
        \raddr_pos_fast[1]_net_1\, \raddr_pos_1_rep1\, 
        \raddr_pos_1_rep2\, \raddr_pos_fast_fast[0]_net_1\, 
        \raddr_pos_fast_0_rep1\, \raddr_pos_fast_0_rep2\, N_1653, 
        \data_out_31_1_1[30]\, N_1429, N_949, N_1173, N_1652, 
        \data_out_31_1_1[29]\, N_1428, N_948, N_1172, N_1647, 
        \data_out_31_1_1[24]\, N_1423, N_943, N_1167, N_1646, 
        \data_out_31_1_1[23]\, N_1422, N_942, N_1166, N_1644, 
        \data_out_31_1_1[21]\, N_1420, N_940, N_1164, N_1641, 
        \data_out_31_1_1[18]\, N_1417, N_937, N_1161, N_1640, 
        \data_out_31_1_1[17]\, N_1416, N_936, N_1160, N_1637, 
        \data_out_31_1_1[14]\, N_1413, N_933, N_1157, N_1626, 
        \data_out_31_1_1[3]\, N_1402, N_922, N_1146, N_1627, 
        \data_out_31_1_1[4]\, N_1403, N_923, N_1147, N_1643, 
        \data_out_31_1_1[20]\, N_1419, N_939, N_1163, N_1639, 
        \data_out_31_1_1[16]\, N_1415, N_935, N_1159, N_1651, 
        \data_out_31_1_1[28]\, N_1427, N_947, N_1171, N_1636, 
        \data_out_31_1_1[13]\, N_1412, N_932, N_1156, N_1650, 
        \data_out_31_1_1[27]\, N_1426, N_946, N_1170, N_1633, 
        \data_out_31_1_1[10]\, N_1409, N_929, N_1153, N_1629, 
        \data_out_31_1_1[6]\, N_1405, N_925, N_1149, N_1642, 
        \data_out_31_1_1[19]\, N_1418, N_938, N_1162, N_1632, 
        \data_out_31_1_1[9]\, N_1408, N_928, N_1152, N_1645, 
        \data_out_31_1_1[22]\, N_1421, N_941, N_1165, N_1634, 
        \data_out_31_1_1[11]\, N_1410, N_930, N_1154, N_1635, 
        \data_out_31_1_1[12]\, N_1411, N_931, N_1155, N_1630, 
        \data_out_31_1_1[7]\, N_1406, N_926, N_1150, N_1638, 
        \data_out_31_1_1[15]\, N_1414, N_934, N_1158, N_1648, 
        \data_out_31_1_1[25]\, N_1424, N_944, N_1168, N_1631, 
        \data_out_31_1_1[8]\, N_1407, N_927, N_1151, N_1628, 
        \data_out_31_1_1[5]\, N_1404, N_924, N_1148, N_1654, 
        \data_out_31_1_1[31]\, N_1430, N_950, N_1174, N_1649, 
        \data_out_31_1_1[26]\, N_1425, N_945, N_1169, 
        \data_out_14_1_1[17]\, \data_out_22_1_1[30]\, 
        \data_out_14_1_1[7]\, \data_out_14_1_1[18]\, 
        \data_out_29_1_1[19]\, \data_out_22_1_1[19]\, 
        \data_out_22_1_1[24]\, \data_out_14_1_1[21]\, 
        \data_out_22_1_1[8]\, \data_out_7_1_1[15]\, 
        \data_out_29_1_1[6]\, \data_out_22_1_1[6]\, 
        \data_out_14_1_1[25]\, \data_out_14_1_1[1]\, 
        \data_out_7_1_1[7]\, \data_out_14_1_1[10]\, 
        \data_out_14_1_1[19]\, \data_out_14_1_1[30]\, 
        \data_out_29_1_1[7]\, \data_out_22_1_1[25]\, 
        \data_out_7_1_1[21]\, \data_out_7_1_1[20]\, 
        \data_out_7_1_1[18]\, \data_out_29_1_1[20]\, 
        \data_out_22_1_1[27]\, \data_out_7_1_1[23]\, 
        \data_out_7_1_1[22]\, \data_out_22_1_1[29]\, 
        \data_out_14_1_1[20]\, \data_out_7_1_1[14]\, 
        \data_out_7_1_1[29]\, \data_out_7_1_1[28]\, 
        \data_out_7_1_1[10]\, \data_out_7_1_1[2]\, 
        \data_out_14_1_1[27]\, \data_out_22_1_1[2]\, 
        \data_out_29_1_1[9]\, \data_out_14_1_1[2]\, 
        \data_out_14_1_1[29]\, \data_out_14_1_1[16]\, 
        \data_out_7_1_1[27]\, \data_out_29_1_1[13]\, 
        \data_out_14_1_1[28]\, \data_out_14_1_1[12]\, 
        \data_out_14_1_1[11]\, \data_out_7_1_1[8]\, 
        \data_out_14_1_1[14]\, \data_out_22_1_1[5]\, 
        \data_out_29_1_1[28]\, \data_out_7_1_1[16]\, 
        \data_out_29_1_1[14]\, \data_out_14_1_1[13]\, 
        \data_out_14_1_1[3]\, \data_out_22_1_1[22]\, 
        \data_out_22_1_1[21]\, \data_out_7_1_1[0]\, 
        \data_out_22_1_1[17]\, \data_out_22_1_1[15]\, 
        \data_out_14_1_1[31]\, \data_out_22_1_1[28]\, 
        \data_out_22_1_1[23]\, \data_out_22_1_1[1]\, 
        \data_out_7_1_1[6]\, \data_out_29_1_1[22]\, 
        \data_out_29_1_1[21]\, \data_out_7_1_1[30]\, 
        \data_out_7_1_1[26]\, \data_out_7_1_1[17]\, 
        \data_out_29_1_1[0]\, \data_out_7_1_1[19]\, 
        \data_out_7_1_1[24]\, \data_out_7_1_1[31]\, 
        \data_out_7_1_1[9]\, \data_out_7_1_1[1]\, 
        \data_out_14_1_1[8]\, \data_out_14_1_1[0]\, 
        \data_out_22_1_1[13]\, \data_out_22_1_1[12]\, 
        \data_out_29_1_1[31]\, \data_out_29_1_1[27]\, 
        \data_out_29_1_1[26]\, \data_out_29_1_1[23]\, 
        \data_out_14_1_1[6]\, \data_out_29_1_1[18]\, 
        \data_out_29_1_1[16]\, \data_out_29_1_1[12]\, 
        \data_out_14_1_1[4]\, \data_out_14_1_1[23]\, 
        \data_out_14_1_1[22]\, \data_out_14_1_1[15]\, 
        \data_out_29_1_1[8]\, \data_out_29_1_1[29]\, 
        \data_out_29_1_1[30]\, \data_out_22_1_1[16]\, 
        \data_out_29_1_1[3]\, \data_out_29_1_1[5]\, 
        \data_out_7_1_1[5]\, \data_out_22_1_1[7]\, 
        \data_out_29_1_1[4]\, \data_out_22_1_1[31]\, 
        \data_out_22_1_1[11]\, \data_out_7_1_1[11]\, 
        \data_out_22_1_1[4]\, \data_out_29_1_1[15]\, 
        \data_out_29_1_1[1]\, \data_out_22_1_1[9]\, 
        \data_out_22_1_1[20]\, \data_out_22_1_1[18]\, 
        \data_out_14_1_1[24]\, \data_out_7_1_1[13]\, 
        \data_out_29_1_1[17]\, \data_out_29_1_1[24]\, 
        \data_out_29_1_1[11]\, \data_out_29_1_1[10]\, 
        \data_out_7_1_1[12]\, \data_out_29_1_1[2]\, 
        \data_out_14_1_1[26]\, \data_out_7_1_1[3]\, 
        \data_out_22_1_1[0]\, \data_out_22_1_1[3]\, 
        \data_out_14_1_1[5]\, \data_out_14_1_1[9]\, 
        \data_out_7_1_1[25]\, \data_out_22_1_1[10]\, 
        \data_out_29_1_1[25]\, \data_out_7_1_1[4]\, 
        \data_out_22_1_1[26]\, \data_out_22_1_1[14]\, N_49, 
        N_49_mux, N_13_0, N_39, N_30, N_23_0, N_15_0 : std_logic;

begin 

    raddr_pos_3 <= \raddr_pos_3\;
    raddr_pos_2 <= \raddr_pos_2\;
    SHA256_Module_0_data_out_ready <= 
        \SHA256_Module_0_data_out_ready\;
    SHA256_Module_0_data_available <= 
        \SHA256_Module_0_data_available\;

    \line6_RNIT2FG1[63]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[31]\, C => \line7[63]_net_1\, D => 
        \line6[63]_net_1\, Y => N_1654);
    
    m43 : CFG4
      generic map(INIT => x"1302")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_39, Y => 
        line6_0_62);
    
    \line3[15]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[15]_net_1\);
    
    \raddr_pos_RNIMPIB8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1646, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[23]\, D => N_1422, Y => N_1710);
    
    \line5[19]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[19]_net_1\);
    
    \line3[41]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[41]_net_1\);
    
    \line1[30]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[30]_net_1\);
    
    \line1[16]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[16]_net_1\);
    
    \line6_RNIRK9N[7]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line7[7]_net_1\, B => \line6[7]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_29_1_1[7]\);
    
    \line6[17]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[17]_net_1\);
    
    \line1[22]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[22]_net_1\);
    
    \raddr_pos_RNIO2PV6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1641, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[18]\, D => N_1417, Y => N_1705);
    
    \line7[61]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[61]_net_1\);
    
    \line0_RNIAIA32[35]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[3]\, 
        C => \line1[35]_net_1\, D => \line0[35]_net_1\, Y => 
        N_922);
    
    \line5[33]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[33]_net_1\);
    
    \line3[0]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[0]_net_1\);
    
    \line6[45]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[45]_net_1\);
    
    \line1[14]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[14]_net_1\);
    
    \line0_RNI9Q422[47]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[15]\, 
        C => \line1[47]_net_1\, D => \line0[47]_net_1\, Y => 
        N_934);
    
    \raddr_pos_fast[1]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_fast[1]_net_1\);
    
    \line0_RNI5FUU1[39]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_7_1_1[7]\, C => \line1[39]_net_1\, D => 
        \line0[39]_net_1\, Y => N_926);
    
    \line7[27]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[27]_net_1\);
    
    \raddr_pos_RNIO4C07[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1630, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[7]\, D => N_1406, Y => N_1694);
    
    \line4_RNI9JQE2[59]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[27]\, C => \line5[59]_net_1\, D => 
        \line4[59]_net_1\, Y => N_1426);
    
    \line1[11]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[11]_net_1\);
    
    \line7[47]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[47]_net_1\);
    
    \line2_RNIJ6151[9]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[9]_net_1\, B => \line2[9]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[9]\);
    
    \raddr_pos_RNIKSDB3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_939, 
        D => N_1163, Y => \data_out_31_1_1[20]\);
    
    \line2[50]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[50]_net_1\);
    
    \raddr_pos_RNIBD6B3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_933, 
        D => N_1157, Y => \data_out_31_1_1[14]\);
    
    \line0[32]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[32]_net_1\);
    
    m40 : CFG4
      generic map(INIT => x"2301")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_39, Y => 
        line7_0_62);
    
    m14 : CFG4
      generic map(INIT => x"2F0D")

      port map(A => waddr_in_net_0(3), B => waddr_in_net_0(2), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_13_0, Y => 
        N_15_0);
    
    \line6[20]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[20]_net_1\);
    
    \line1[56]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[56]_net_1\);
    
    \line3[36]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[36]_net_1\);
    
    \line3[4]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[4]_net_1\);
    
    \line0[20]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[20]_net_1\);
    
    \line6[55]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[55]_net_1\);
    
    \line0[56]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[56]_net_1\);
    
    \line0_RNIV9O01[10]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[10]_net_1\, B => \line0[10]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[10]\);
    
    \line0_RNITND31[31]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line0[31]_net_1\, B => \line1[31]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_7_1_1[31]\);
    
    \line2[49]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[49]_net_1\);
    
    \raddr_pos_RNIFQRB8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1652, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[29]\, D => N_1428, Y => N_1716);
    
    \line2_RNIHQL31[47]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_14_1_1[15]\, C => \line3[47]_net_1\, D => 
        \line2[47]_net_1\, Y => N_1158);
    
    \line2[20]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[20]_net_1\);
    
    \line7[12]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[12]_net_1\);
    
    \line5[22]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[22]_net_1\);
    
    \line4_RNIKC4F1[36]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[4]\, C => \line5[36]_net_1\, D => 
        \line4[36]_net_1\, Y => N_1403);
    
    \line3[61]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[61]_net_1\);
    
    \line3[29]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[29]_net_1\);
    
    \line1[54]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[54]_net_1\);
    
    \line5[38]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[38]_net_1\);
    
    \line3[34]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[34]_net_1\);
    
    \line3[7]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[7]_net_1\);
    
    \line4[61]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[61]_net_1\);
    
    \line0[54]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[54]_net_1\);
    
    \line0[8]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[8]_net_1\);
    
    \line0[49]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[49]_net_1\);
    
    \line7[52]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[52]_net_1\);
    
    \raddr_pos_RNIJ0AG4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_924, 
        D => N_1148, Y => \data_out_31_1_1[5]\);
    
    \line2_RNICUP61[63]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[31]\, C => \line3[63]_net_1\, D => 
        \line2[63]_net_1\, Y => N_1174);
    
    \line1[51]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[51]_net_1\);
    
    \line4[50]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[50]_net_1\);
    
    \line3[31]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[31]_net_1\);
    
    \line2_RNIDB3K1[39]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_14_1_1[7]\, C => \line3[39]_net_1\, D => 
        \line2[39]_net_1\, Y => N_1150);
    
    \line0[51]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[51]_net_1\);
    
    \line5[42]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[42]_net_1\);
    
    \line0_RNI6UR82[55]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[23]\, C => \line1[55]_net_1\, D => 
        \line0[55]_net_1\, Y => N_942);
    
    \line2[16]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[16]_net_1\);
    
    \raddr_pos_RNI6AJB8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1647, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[24]\, D => N_1423, Y => N_1711);
    
    \ren_pos\ : SLE
      port map(D => data_out_ready_0_sqmuxa, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ren_pos);
    
    \line6[60]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[60]_net_1\);
    
    m16 : CFG4
      generic map(INIT => x"2301")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_15_0, Y => 
        line5_0_62);
    
    \line1[23]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[23]_net_1\);
    
    \line4[8]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[8]_net_1\);
    
    \line3[55]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[55]_net_1\);
    
    \line7[30]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[30]_net_1\);
    
    \line0_RNIR60V1[41]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_7_1_1[9]\, C => \line1[41]_net_1\, D => 
        \line0[41]_net_1\, Y => N_928);
    
    \line6[2]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[2]_net_1\);
    
    \line4[0]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[0]_net_1\);
    
    \line4[42]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[42]_net_1\);
    
    \line2[14]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[14]_net_1\);
    
    \line7[4]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[4]_net_1\);
    
    \line0_RNI6ASR1[44]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[12]\, 
        C => \line1[44]_net_1\, D => \line0[44]_net_1\, Y => 
        N_931);
    
    \line0_RNI26SR1[43]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[11]\, 
        C => \line1[43]_net_1\, D => \line0[43]_net_1\, Y => 
        N_930);
    
    \raddr_pos_RNIU9RB8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1651, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[28]\, D => N_1427, Y => N_1715);
    
    \line1[49]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[49]_net_1\);
    
    \raddr_pos_RNI2AMG7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1638, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[15]\, D => N_1414, Y => N_1702);
    
    \line2[11]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[11]_net_1\);
    
    raddr_pos_fast_0_rep1 : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_fast_0_rep1\);
    
    \line3[2]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[2]_net_1\);
    
    \line0_RNIN20V1[40]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_7_1_1[8]\, C => \line1[40]_net_1\, D => 
        \line0[40]_net_1\, Y => N_927);
    
    \line4[32]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[32]_net_1\);
    
    \line4[16]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[16]_net_1\);
    
    \line2[32]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[32]_net_1\);
    
    \line6_RNIHEAP[18]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[18]_net_1\, B => \line6[18]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[18]\);
    
    \line4[7]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[7]_net_1\);
    
    \line6_RNIOO8S[29]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[29]_net_1\, B => \line6[29]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[29]\);
    
    \line5[17]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[17]_net_1\);
    
    \line3[9]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[9]_net_1\);
    
    \line0[33]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[33]_net_1\);
    
    \line4[1]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[1]_net_1\);
    
    \line1[35]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[35]_net_1\);
    
    \line3[49]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[49]_net_1\);
    
    \raddr_pos_RNIA8EE4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_923, 
        D => N_1147, Y => \data_out_31_1_1[4]\);
    
    \line0[12]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[12]_net_1\);
    
    \raddr_pos_RNIV3JM3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_934, 
        D => N_1158, Y => \data_out_31_1_1[15]\);
    
    \raddr_pos_RNILBRS3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_950, 
        D => N_1174, Y => \data_out_31_1_1[31]\);
    
    \line2_RNI4UKC1[0]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[0]_net_1\, B => \line2[0]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[0]\);
    
    \line4[14]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[14]_net_1\);
    
    \line2_RNICC7P[22]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[22]_net_1\, B => \line2[22]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[22]\);
    
    \line7[13]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[13]_net_1\);
    
    \line2_RNI0B3U[53]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[21]\, C => \line3[53]_net_1\, D => 
        \line2[53]_net_1\, Y => N_1164);
    
    \line1[28]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[28]_net_1\);
    
    \line5[23]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[23]_net_1\);
    
    m2 : CFG2
      generic map(INIT => x"D")

      port map(A => sha256_system_sb_0_GPIO_9_M2F, B => 
        sha256_system_sb_0_GPIO_1_M2F, Y => N_3_0);
    
    \line2[4]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[4]_net_1\);
    
    \line6_RNI54CP[21]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[21]_net_1\, B => \line6[21]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[21]\);
    
    \line6[1]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[1]_net_1\);
    
    \line0_RNI2PA11[19]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[19]_net_1\, B => \line0[19]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[19]\);
    
    \line4[11]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[11]_net_1\);
    
    \line6[30]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[30]_net_1\);
    
    \line2_RNI82LC1[2]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[2]_net_1\, B => \line2[2]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[2]\);
    
    \line6_RNIPUEG1[62]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[30]\, C => \line7[62]_net_1\, D => 
        \line6[62]_net_1\, Y => N_1653);
    
    \line7[53]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[53]_net_1\);
    
    \line0_RNIJ6IS1[52]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[20]\, 
        C => \line1[52]_net_1\, D => \line0[52]_net_1\, Y => 
        N_939);
    
    \line6_RNI7BDG1[61]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[29]\, C => \line7[61]_net_1\, D => 
        \line6[61]_net_1\, Y => N_1652);
    
    \line7[7]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[7]_net_1\);
    
    \line1[19]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[19]_net_1\);
    
    \line1[0]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[0]_net_1\);
    
    \line0_RNIUKA11[17]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[17]_net_1\, B => \line0[17]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[17]\);
    
    \line5[43]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[43]_net_1\);
    
    \line4[20]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[20]_net_1\);
    
    \line2[55]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[55]_net_1\);
    
    \line0_RNIVEES1[46]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[14]\, 
        C => \line1[46]_net_1\, D => \line0[46]_net_1\, Y => 
        N_933);
    
    \line5[50]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[50]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line6[25]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[25]_net_1\);
    
    \line3[1]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[1]_net_1\);
    
    \line0[38]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[38]_net_1\);
    
    \line2[47]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[47]_net_1\);
    
    \raddr_pos_RNIN9Q34[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_926, 
        D => N_1150, Y => \data_out_31_1_1[7]\);
    
    \line7_or[32]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line7_0, B => sha256_system_sb_0_GPIO_9_M2F, 
        Y => \line7_or[32]_net_1\);
    
    \line4_RNI9QH81[16]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[16]_net_1\, B => \line4[16]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[16]\);
    
    \line0_RNIUPV82[62]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[30]\, C => \line1[62]_net_1\, D => 
        \line0[62]_net_1\, Y => N_949);
    
    \line0[25]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[25]_net_1\);
    
    \line0_RNINE652[38]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[6]\, 
        C => \line1[38]_net_1\, D => \line0[38]_net_1\, Y => 
        N_925);
    
    \line3[27]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[27]_net_1\);
    
    \line2[25]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[25]_net_1\);
    
    \line6_RNI20AP[11]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[11]_net_1\, B => \line6[11]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[11]\);
    
    \line4[43]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[43]_net_1\);
    
    \line7[18]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[18]_net_1\);
    
    \line3[12]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[12]_net_1\);
    
    \line5[28]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[28]_net_1\);
    
    \line0[47]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[47]_net_1\);
    
    \line4_RNI6SHB1[31]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[31]_net_1\, B => \line4[31]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[31]\);
    
    \line5[36]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[36]_net_1\);
    
    \line4[33]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[33]_net_1\);
    
    \line6_RNIKEN61[44]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[12]\, C => \line7[44]_net_1\, D => 
        \line6[44]_net_1\, Y => N_1635);
    
    \line2[33]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[33]_net_1\);
    
    \line7[58]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[58]_net_1\);
    
    \line4[55]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[55]_net_1\);
    
    \line1[59]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[59]_net_1\);
    
    \line3[39]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[39]_net_1\);
    
    \raddr_pos_RNI04IV6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1639, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[16]\, D => N_1415, Y => N_1703);
    
    \line0[59]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[59]_net_1\);
    
    \line4_RNIRCTI[9]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line5[9]_net_1\, B => \line4[9]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_22_1_1[9]\);
    
    \line5[48]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[48]_net_1\);
    
    \line0[13]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[13]_net_1\);
    
    \line6[42]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[42]_net_1\);
    
    \line6_RNIKK8S[27]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[27]_net_1\, B => \line6[27]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[27]\);
    
    \line5[34]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[34]_net_1\);
    
    \line4_RNISDH81[10]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[10]_net_1\, B => \line4[10]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[10]\);
    
    \line1[9]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[9]_net_1\);
    
    \line1_or[32]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line1_0, B => sha256_system_sb_0_GPIO_9_M2F, 
        Y => \line1_or[32]_net_1\);
    
    \line4_RNIBSH81[17]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[17]_net_1\, B => \line4[17]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[17]\);
    
    \line3[5]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[5]_net_1\);
    
    \line3[8]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[8]_net_1\);
    
    \raddr_pos_RNIFLAB3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_938, 
        D => N_1162, Y => \data_out_31_1_1[19]\);
    
    \line6_RNIO4941[35]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[3]\, C => \line7[35]_net_1\, D => 
        \line6[35]_net_1\, Y => N_1626);
    
    \line2_RNI7FVT[46]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[14]\, C => \line3[46]_net_1\, D => 
        \line2[46]_net_1\, Y => N_1157);
    
    \line7[35]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[35]_net_1\);
    
    \line5[31]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[31]_net_1\);
    
    \line4_RNI1KJ81[21]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[21]_net_1\, B => \line4[21]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[21]\);
    
    \line1[47]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[47]_net_1\);
    
    \line6[10]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[10]_net_1\);
    
    \line1[7]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[7]_net_1\);
    
    \line1[60]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[60]_net_1\);
    
    \line4[48]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[48]_net_1\);
    
    \line0[62]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[62]_net_1\);
    
    \raddr_pos_RNIT4EB3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_940, 
        D => N_1164, Y => \data_out_31_1_1[21]\);
    
    \line0_RNIOAIS1[53]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[21]\, 
        C => \line1[53]_net_1\, D => \line0[53]_net_1\, Y => 
        N_940);
    
    \line0_RNIDE4A1[6]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[6]_net_1\, B => \line0[6]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[6]\);
    
    \line6_RNID8JL[15]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[15]_net_1\, B => \line7[15]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[15]\);
    
    \line2[6]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[6]_net_1\);
    
    \line6[52]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[52]_net_1\);
    
    \line2[19]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[19]_net_1\);
    
    \line6_RNI74AP[13]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[13]_net_1\, B => \line6[13]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[13]\);
    
    \line2_RNI5F1U[50]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[18]\, C => \line3[50]_net_1\, D => 
        \line2[50]_net_1\, Y => N_1161);
    
    \line2_RNIQS2I[13]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[13]_net_1\, B => \line2[13]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[13]\);
    
    \line4[38]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[38]_net_1\);
    
    \line3[47]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[47]_net_1\);
    
    \line2[38]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[38]_net_1\);
    
    \line7[20]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[20]_net_1\);
    
    \line6_RNIBQAG[5]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[5]_net_1\, B => \line7[5]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[5]\);
    
    \line7[40]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[40]_net_1\);
    
    \line2_RNIBIRN[28]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[28]_net_1\, B => \line2[28]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_14_1_1[28]\);
    
    \line0[18]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[18]_net_1\);
    
    \line2_RNI335K1[41]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_14_1_1[9]\, C => \line3[41]_net_1\, D => 
        \line2[41]_net_1\, Y => N_1152);
    
    \line2_RNIEKRN[29]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[29]_net_1\, B => \line2[29]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep2\, Y => 
        \data_out_14_1_1[29]\);
    
    \line2[3]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[3]_net_1\);
    
    \line3[13]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[13]_net_1\);
    
    \line7[0]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[0]_net_1\);
    
    \line1[26]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[26]_net_1\);
    
    \line4_RNIK8GB1[29]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[29]_net_1\, B => \line4[29]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[29]\);
    
    \line4[19]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[19]_net_1\);
    
    \line2_RNINQ4I[20]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[20]_net_1\, B => \line2[20]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[20]\);
    
    \line7[1]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[1]_net_1\);
    
    \line6[35]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[35]_net_1\);
    
    \line1[17]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[17]_net_1\);
    
    \line5[9]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[9]_net_1\);
    
    \line4[25]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[25]_net_1\);
    
    \line3[52]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[52]_net_1\);
    
    \line5[62]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[62]_net_1\);
    
    \line1[24]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[24]_net_1\);
    
    \line5[55]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[55]_net_1\);
    
    \line6[43]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[43]_net_1\);
    
    \line0_RNILCC11[21]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[21]_net_1\, B => \line0[21]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[21]\);
    
    \line0_RNIMES82[59]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[27]\, C => \line1[59]_net_1\, D => 
        \line0[59]_net_1\, Y => N_946);
    
    m27 : CFG4
      generic map(INIT => x"1302")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_23_0, Y => 
        line2_0_62);
    
    \line6[5]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[5]_net_1\);
    
    \line1[21]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[21]_net_1\);
    
    \line0[36]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[36]_net_1\);
    
    \line4_RNIHUTE2[62]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[30]\, C => \line5[62]_net_1\, D => 
        \line4[62]_net_1\, Y => N_1429);
    
    \line0_RNIU5A32[32]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[0]\, 
        C => \line1[32]_net_1\, D => \line0[32]_net_1\, Y => 
        N_919);
    
    \line0_RNIDSK32[54]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[22]\, 
        C => \line1[54]_net_1\, D => \line0[54]_net_1\, Y => 
        N_941);
    
    \line0_RNI6O881[3]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[3]_net_1\, B => \line0[3]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[3]\);
    
    \line7[5]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[5]_net_1\);
    
    \line1[2]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[2]_net_1\);
    
    \line6_RNI1GAG[0]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[0]_net_1\, B => \line7[0]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[0]\);
    
    \line0[63]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[63]_net_1\);
    
    \line6_RNIDAAP[16]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[16]_net_1\, B => \line6[16]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[16]\);
    
    \line3[18]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[18]_net_1\);
    
    \line7[16]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[16]_net_1\);
    
    \raddr_pos_RNI6S544[2]\ : CFG4
      generic map(INIT => x"4567")

      port map(A => \raddr_pos_2\, B => \raddr_pos_3\, C => N_948, 
        D => N_1172, Y => \data_out_31_1_1[29]\);
    
    \line5[26]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[26]_net_1\);
    
    \line1[32]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[32]_net_1\);
    
    \line1[57]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[57]_net_1\);
    
    \line6[53]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[53]_net_1\);
    
    \line0[34]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[34]_net_1\);
    
    \line3[37]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[37]_net_1\);
    
    \line0_RNIVN071[15]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[15]_net_1\, B => \line0[15]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_7_1_1[15]\);
    
    \line4_RNIBBGF1[39]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_22_1_1[7]\, 
        C => \line5[39]_net_1\, D => \line4[39]_net_1\, Y => 
        N_1406);
    
    \line6_RNI0D941[37]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[5]\, C => \line7[37]_net_1\, D => 
        \line6[37]_net_1\, Y => N_1628);
    
    \line0[57]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[57]_net_1\);
    
    \line8_or[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line8_0_62, B => 
        sha256_system_sb_0_GPIO_9_M2F, Y => \line8_or[0]_net_1\);
    
    \line6_RNI9BBG1[57]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[25]\, C => \line7[57]_net_1\, D => 
        \line6[57]_net_1\, Y => N_1648);
    
    \line0[31]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[31]_net_1\);
    
    \line7[56]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[56]_net_1\);
    
    \line2_RNIU5TN[30]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[30]_net_1\, B => \line2[30]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep2\, Y => 
        \data_out_14_1_1[30]\);
    
    \line6_or[32]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line6_0, B => sha256_system_sb_0_GPIO_9_M2F, 
        Y => \line6_or[32]_net_1\);
    
    \line0_RNI3U271[26]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[26]_net_1\, B => \line0[26]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_7_1_1[26]\);
    
    \line0_RNI4M881[2]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[2]_net_1\, B => \line0[2]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[2]\);
    
    \line7[14]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[14]_net_1\);
    
    \line5[24]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[24]_net_1\);
    
    \line8[1]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line8_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => last_block);
    
    \line6[48]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[48]_net_1\);
    
    \line5[10]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[10]_net_1\);
    
    \line5[46]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[46]_net_1\);
    
    \line2_RNIH4151[8]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[8]_net_1\, B => \line2[8]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[8]\);
    
    \line2[7]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[7]_net_1\);
    
    \line0_RNITN271[23]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[23]_net_1\, B => \line0[23]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_7_1_1[23]\);
    
    \line4_RNINQ852[51]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[19]\, C => \line5[51]_net_1\, D => 
        \line4[51]_net_1\, Y => N_1418);
    
    \raddr_pos_RNIE64C7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1628, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[5]\, D => N_1404, Y => N_1692);
    
    \line7[11]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[11]_net_1\);
    
    m32 : CFG4
      generic map(INIT => x"8C04")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_30, Y => 
        line1_0);
    
    \line5[21]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[21]_net_1\);
    
    \line4[6]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[6]_net_1\);
    
    \line7[54]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[54]_net_1\);
    
    \line4_RNI8A652[43]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[11]\, C => \line5[43]_net_1\, D => 
        \line4[43]_net_1\, Y => N_1410);
    
    \line5[39]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[39]_net_1\);
    
    \line4_RNI46652[42]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[10]\, C => \line5[42]_net_1\, D => 
        \line4[42]_net_1\, Y => N_1409);
    
    \line2[52]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[52]_net_1\);
    
    \line6[15]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[15]_net_1\);
    
    \line4_RNIDIA52[53]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[21]\, C => \line5[53]_net_1\, D => 
        \line4[53]_net_1\, Y => N_1420);
    
    \line2[17]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[17]_net_1\);
    
    \line5[44]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[44]_net_1\);
    
    \line4_RNIF0I81[19]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[19]_net_1\, B => \line4[19]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[19]\);
    
    \line7[51]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[51]_net_1\);
    
    \line6[22]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[22]_net_1\);
    
    \line4[46]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[46]_net_1\);
    
    \line4_RNIVHJ81[20]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[20]_net_1\, B => \line4[20]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[20]\);
    
    \line0[22]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[22]_net_1\);
    
    \line6[58]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[58]_net_1\);
    
    \line3[53]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[53]_net_1\);
    
    \line5[63]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[63]_net_1\);
    
    \raddr_pos_RNIPB144[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_942, 
        D => N_1166, Y => \data_out_31_1_1[23]\);
    
    \line5[41]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[41]_net_1\);
    
    \line6_RNI57BG1[56]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[24]\, C => \line7[56]_net_1\, D => 
        \line6[56]_net_1\, Y => N_1647);
    
    \line2[22]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[22]_net_1\);
    
    \line7[25]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[25]_net_1\);
    
    \line4_RNITUHF1[40]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_22_1_1[8]\, 
        C => \line5[40]_net_1\, D => \line4[40]_net_1\, Y => 
        N_1407);
    
    \line4[36]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[36]_net_1\);
    
    \line2[36]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[36]_net_1\);
    
    \line4_RNI5FQE2[58]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[26]\, C => \line5[58]_net_1\, D => 
        \line4[58]_net_1\, Y => N_1425);
    
    \line4_RNISK4F1[38]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[6]\, C => \line5[38]_net_1\, D => 
        \line4[38]_net_1\, Y => N_1405);
    
    \line2[2]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[2]_net_1\);
    
    \line4[9]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[9]_net_1\);
    
    \line2_RNI693I[19]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[19]_net_1\, B => \line2[19]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[19]\);
    
    \line7[45]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[45]_net_1\);
    
    \line4[44]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[44]_net_1\);
    
    \line0[16]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[16]_net_1\);
    
    \line4[17]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[17]_net_1\);
    
    \line4[41]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[41]_net_1\);
    
    \line2[40]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[40]_net_1\);
    
    \line6_RNIMM8S[28]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[28]_net_1\, B => \line6[28]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[28]\);
    
    \line4[52]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[52]_net_1\);
    
    \line2_RNIPS4I[21]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[21]_net_1\, B => \line2[21]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[21]\);
    
    \line4[34]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[34]_net_1\);
    
    \line0[0]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[0]_net_1\);
    
    \line2[34]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[34]_net_1\);
    
    \line4_RNIOG4F1[37]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[5]\, C => \line5[37]_net_1\, D => 
        \line4[37]_net_1\, Y => N_1404);
    
    \raddr_pos_RNI8JPV6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1642, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[19]\, D => N_1418, Y => N_1706);
    
    \line6[6]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[6]_net_1\);
    
    \line1[33]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[33]_net_1\);
    
    \line3[20]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[20]_net_1\);
    
    \line0_RNI2K881[1]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[1]_net_1\, B => \line0[1]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[1]\);
    
    \raddr_pos_RNI1GIC4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_922, 
        D => N_1146, Y => \data_out_31_1_1[3]\);
    
    \line4[31]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[31]_net_1\);
    
    \line2[31]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[31]_net_1\);
    
    \line6[62]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[62]_net_1\);
    
    \line0[14]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[14]_net_1\);
    
    \line6_RNIQQED1[54]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[22]\, C => \line7[54]_net_1\, D => 
        \line6[54]_net_1\, Y => N_1645);
    
    \line2_RNIFNVT[48]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[16]\, C => \line3[48]_net_1\, D => 
        \line2[48]_net_1\, Y => N_1159);
    
    \line0[40]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[40]_net_1\);
    
    \raddr_pos_RNIO99D3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_929, 
        D => N_1153, Y => \data_out_31_1_1[10]\);
    
    \line6_RNIGG8S[25]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[25]_net_1\, B => \line6[25]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[25]\);
    
    \raddr_pos_RNIS8CU6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1635, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[12]\, D => N_1411, Y => N_1699);
    
    \line7[32]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[32]_net_1\);
    
    \line3[58]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[58]_net_1\);
    
    \line0_RNIDOK01[8]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[8]_net_1\, B => \line0[8]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[8]\);
    
    \line5_or[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line5_0_62, B => 
        sha256_system_sb_0_GPIO_9_M2F, Y => \line5_or[0]_net_1\);
    
    \line0[11]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[11]_net_1\);
    
    m22 : CFG4
      generic map(INIT => x"4F0B")

      port map(A => waddr_in_net_0(3), B => waddr_in_net_0(2), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_13_0, Y => 
        N_23_0);
    
    m29 : CFG4
      generic map(INIT => x"1F0E")

      port map(A => waddr_in_net_0(3), B => waddr_in_net_0(2), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_13_0, Y => N_30);
    
    \line5[1]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[1]_net_1\);
    
    \line4_RNIN8TI[7]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line5[7]_net_1\, B => \line4[7]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_22_1_1[7]\);
    
    \line1[29]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[29]_net_1\);
    
    \line2[60]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[60]_net_1\);
    
    \line6[0]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[0]_net_1\);
    
    m34 : CFG4
      generic map(INIT => x"1302")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_30, Y => 
        line0_0_62);
    
    \line2[53]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[53]_net_1\);
    
    \line1[8]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[8]_net_1\);
    
    \line5[8]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[8]_net_1\);
    
    \line6_RNIFCAP[17]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[17]_net_1\, B => \line6[17]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[17]\);
    
    \line0_RNI50371[27]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[27]_net_1\, B => \line0[27]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_7_1_1[27]\);
    
    \line6[23]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[23]_net_1\);
    
    \line6_RNIACAS[31]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[31]_net_1\, B => \line6[31]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[31]\);
    
    \line0[23]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[23]_net_1\);
    
    \line3[16]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[16]_net_1\);
    
    \line1[38]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[38]_net_1\);
    
    \line1[40]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[40]_net_1\);
    
    \line0_RNIC6U82[61]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[29]\, C => \line1[61]_net_1\, D => 
        \line0[61]_net_1\, Y => N_948);
    
    \line4_RNIT6QE2[56]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[24]\, C => \line5[56]_net_1\, D => 
        \line4[56]_net_1\, Y => N_1423);
    
    \line4_RNIT3UB[0]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[0]_net_1\, B => \line5[0]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[0]\);
    
    \line4_RNIV5UB[1]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[1]_net_1\, B => \line5[1]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[1]\);
    
    \line2[23]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[23]_net_1\);
    
    raddr_pos_fast_0_rep2 : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_fast_0_rep2\);
    
    \line2_RNIHQGE1[6]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[6]_net_1\, B => \line2[6]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[6]\);
    
    \line0[39]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[39]_net_1\);
    
    \line6_RNIK0941[34]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[2]\, C => \line7[34]_net_1\, D => 
        \line6[34]_net_1\, Y => N_1625);
    
    \line3[14]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[14]_net_1\);
    
    \line5[15]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[15]_net_1\);
    
    \line2_RNIEUCA1[55]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[23]\, C => \line3[55]_net_1\, D => 
        \line2[55]_net_1\, Y => N_1166);
    
    \line6[32]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[32]_net_1\);
    
    \line4_RNI5MH81[14]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[14]_net_1\, B => \line4[14]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[14]\);
    
    \raddr_pos_RNIT58A7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1627, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[4]\, D => N_1403, Y => N_1691);
    
    \line3[40]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[40]_net_1\);
    
    \line2_RNI38PN[15]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[15]_net_1\, B => \line2[15]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_14_1_1[15]\);
    
    \line5[37]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[37]_net_1\);
    
    \line2_RNI186K[31]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line2[31]_net_1\, B => \line3[31]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_14_1_1[31]\);
    
    \line6[46]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[46]_net_1\);
    
    \line0_RNI8SE81[22]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[22]_net_1\, B => \line0[22]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[22]\);
    
    \line4[53]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[53]_net_1\);
    
    \line7[19]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[19]_net_1\);
    
    \line5[29]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[29]_net_1\);
    
    \line3[11]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[11]_net_1\);
    
    \line4[22]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[22]_net_1\);
    
    m36 : CFG2
      generic map(INIT => x"2")

      port map(A => N_49_mux, B => waddr_in_net_0(0), Y => 
        line8_0_62);
    
    \line6_RNI42AP[12]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[12]_net_1\, B => \line6[12]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[12]\);
    
    \line7[60]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[60]_net_1\);
    
    \line5[52]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[52]_net_1\);
    
    \line2[58]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[58]_net_1\);
    
    \line7[6]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[6]_net_1\);
    
    \line5[5]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[5]_net_1\);
    
    \line7[59]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[59]_net_1\);
    
    \line6[63]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[63]_net_1\);
    
    \line6[28]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[28]_net_1\);
    
    \line6[44]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[44]_net_1\);
    
    \line2[8]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[8]_net_1\);
    
    \raddr_pos_RNIPC244[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_946, 
        D => N_1170, Y => \data_out_31_1_1[27]\);
    
    \line0[28]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[28]_net_1\);
    
    \line6_RNIII8S[26]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[26]_net_1\, B => \line6[26]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[26]\);
    
    \line4_RNIDUH81[18]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[18]_net_1\, B => \line4[18]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[18]\);
    
    \line0_RNIA2S82[56]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[24]\, C => \line1[56]_net_1\, D => 
        \line0[56]_net_1\, Y => N_943);
    
    \line7[33]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[33]_net_1\);
    
    \line5[49]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[49]_net_1\);
    
    \line6[56]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[56]_net_1\);
    
    \line4_RNI9EA52[52]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[20]\, C => \line5[52]_net_1\, D => 
        \line4[52]_net_1\, Y => N_1419);
    
    \line1[10]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[10]_net_1\);
    
    m9_e : CFG4
      generic map(INIT => x"0002")

      port map(A => waddr_in_net_0(4), B => waddr_in_net_0(3), C
         => waddr_in_net_0(2), D => waddr_in_net_0(1), Y => N_49);
    
    \line6[41]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[41]_net_1\);
    
    \line0_RNIFQK01[9]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[9]_net_1\, B => \line0[9]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[9]\);
    
    \line2[28]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[28]_net_1\);
    
    m24 : CFG4
      generic map(INIT => x"2301")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_23_0, Y => 
        line3_0_62);
    
    \line4_RNI3MJ81[22]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[22]_net_1\, B => \line4[22]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[22]\);
    
    \line0[6]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[6]_net_1\);
    
    \line6_RNI32CP[20]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[20]_net_1\, B => \line6[20]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[20]\);
    
    \line5[4]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[4]_net_1\);
    
    \line6_RNILIR61[53]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[21]\, C => \line7[53]_net_1\, D => 
        \line6[53]_net_1\, Y => N_1644);
    
    \line2[1]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[1]_net_1\);
    
    \line6[54]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[54]_net_1\);
    
    \line2_RNI473I[18]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[18]_net_1\, B => \line2[18]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[18]\);
    
    \line2[45]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[45]_net_1\);
    
    \line0_RNI1JGS1[51]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[19]\, 
        C => \line1[51]_net_1\, D => \line0[51]_net_1\, Y => 
        N_938);
    
    \line4_RNII6GB1[28]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[28]_net_1\, B => \line4[28]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[28]\);
    
    \line4[49]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[49]_net_1\);
    
    \line0[61]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[61]_net_1\);
    
    \line4[58]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[58]_net_1\);
    
    \line0_RNIIAS82[58]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[26]\, C => \line1[58]_net_1\, D => 
        \line0[58]_net_1\, Y => N_945);
    
    \line3[25]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[25]_net_1\);
    
    \line2_or[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line2_0_62, B => 
        sha256_system_sb_0_GPIO_9_M2F, Y => \line2_or[0]_net_1\);
    
    \raddr_pos_RNIAPK48[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1654, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[31]\, D => N_1430, Y => N_1718);
    
    \line3[60]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[60]_net_1\);
    
    \raddr_pos_RNIA3944[2]\ : CFG4
      generic map(INIT => x"4567")

      port map(A => \raddr_pos_2\, B => \raddr_pos_3\, C => N_949, 
        D => N_1173, Y => \data_out_31_1_1[30]\);
    
    \line6[51]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[51]_net_1\);
    
    \line4[39]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[39]_net_1\);
    
    \line2[39]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[39]_net_1\);
    
    \line4[60]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[60]_net_1\);
    
    \line0[45]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[45]_net_1\);
    
    \line2_RNILS551[54]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[22]\, C => \line3[54]_net_1\, D => 
        \line2[54]_net_1\, Y => N_1165);
    
    \line6_RNIRMP61[50]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[18]\, C => \line7[50]_net_1\, D => 
        \line6[50]_net_1\, Y => N_1641);
    
    \line4_or[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line4_0_62, B => 
        sha256_system_sb_0_GPIO_9_M2F, Y => \line4_or[0]_net_1\);
    
    \line4_RNIR6SE2[60]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[28]\, C => \line5[60]_net_1\, D => 
        \line4[60]_net_1\, Y => N_1427);
    
    \line4_RNI18UB[2]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[2]_net_1\, B => \line5[2]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[2]\);
    
    \line1[50]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[50]_net_1\);
    
    \line3[30]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[30]_net_1\);
    
    \raddr_pos_RNI03HV6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1637, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[14]\, D => N_1413, Y => N_1701);
    
    \line1[27]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[27]_net_1\);
    
    \line7[38]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[38]_net_1\);
    
    \raddr_pos_RNIFIGV6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1636, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[13]\, D => N_1412, Y => N_1700);
    
    \line0_RNI82U82[60]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[28]\, C => \line1[60]_net_1\, D => 
        \line0[60]_net_1\, Y => N_947);
    
    \line0[50]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[50]_net_1\);
    
    \line0[19]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[19]_net_1\);
    
    \line6[33]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[33]_net_1\);
    
    \line6[12]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[12]_net_1\);
    
    \line3[56]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[56]_net_1\);
    
    \line1[62]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[62]_net_1\);
    
    \line2_RNI253I[17]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[17]_net_1\, B => \line2[17]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[17]\);
    
    data_out_ready : SLE
      port map(D => \data_out_ready_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SHA256_Module_0_data_out_ready\);
    
    \line4[4]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[4]_net_1\);
    
    \line2_RNIF2151[7]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[7]_net_1\, B => \line2[7]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[7]\);
    
    \line2_RNI9J1U[51]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[19]\, C => \line3[51]_net_1\, D => 
        \line2[51]_net_1\, Y => N_1162);
    
    \raddr_pos[3]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_3\);
    
    \line4_RNIGI652[45]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[13]\, C => \line5[45]_net_1\, D => 
        \line4[45]_net_1\, Y => N_1412);
    
    \line2_RNIG2FA1[60]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[28]\, C => \line3[60]_net_1\, D => 
        \line2[60]_net_1\, Y => N_1171);
    
    \line2_RNIDMGE1[4]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[4]_net_1\, B => \line2[4]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[4]\);
    
    m44 : CFG4
      generic map(INIT => x"4C08")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_39, Y => 
        line6_0);
    
    \line4[23]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[23]_net_1\);
    
    \line2_RNIEADT[44]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[12]\, C => \line3[44]_net_1\, D => 
        \line2[44]_net_1\, Y => N_1155);
    
    \line5[53]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[53]_net_1\);
    
    \line0_RNI8Q881[4]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[4]_net_1\, B => \line0[4]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[4]\);
    
    \line6[4]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[4]_net_1\);
    
    \line2_RNIA4LC1[3]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[3]_net_1\, B => \line2[3]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[3]\);
    
    \line7[22]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[22]_net_1\);
    
    \line3[54]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[54]_net_1\);
    
    \line7[42]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[42]_net_1\);
    
    \line6_RNI37DG1[60]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[28]\, C => \line7[60]_net_1\, D => 
        \line6[60]_net_1\, Y => N_1651);
    
    \line0[37]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[37]_net_1\);
    
    \line1[45]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[45]_net_1\);
    
    \line3[51]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[51]_net_1\);
    
    \raddr_pos_RNI6BKB8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1649, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[26]\, D => N_1425, Y => N_1713);
    
    \line5[61]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[61]_net_1\);
    
    \line1[36]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[36]_net_1\);
    
    \line8[0]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line8_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => first_block);
    
    \line2[10]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[10]_net_1\);
    
    \line7_or[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line7_0_62, B => 
        sha256_system_sb_0_GPIO_9_M2F, Y => \line7_or[0]_net_1\);
    
    \raddr_pos_RNIN82C8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1653, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[30]\, D => N_1429, Y => N_1717);
    
    \line2_RNIQADA1[58]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[26]\, C => \line3[58]_net_1\, D => 
        \line2[58]_net_1\, Y => N_1169);
    
    \line2_RNI5CRN[25]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[25]_net_1\, B => \line2[25]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_14_1_1[25]\);
    
    \line0_RNI6EA32[34]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[2]\, 
        C => \line1[34]_net_1\, D => \line0[34]_net_1\, Y => 
        N_921);
    
    \line6_RNI9OAG[4]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[4]_net_1\, B => \line7[4]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[4]\);
    
    \line6_or[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line6_0_62, B => 
        sha256_system_sb_0_GPIO_9_M2F, Y => \line6_or[0]_net_1\);
    
    \line7[3]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[3]_net_1\);
    
    \line2_RNI3BVT[45]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[13]\, C => \line3[45]_net_1\, D => 
        \line2[45]_net_1\, Y => N_1156);
    
    \raddr_pos_RNIH4244[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_945, 
        D => N_1169, Y => \data_out_31_1_1[26]\);
    
    \line6_RNI5RM41[40]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_29_1_1[8]\, 
        C => \line7[40]_net_1\, D => \line6[40]_net_1\, Y => 
        N_1631);
    
    \line2_RNI7QGA1[62]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[30]\, C => \line3[62]_net_1\, D => 
        \line2[62]_net_1\, Y => N_1173);
    
    \line7[17]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[17]_net_1\);
    
    \line6_RNIVO9N[9]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line7[9]_net_1\, B => \line6[9]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_29_1_1[9]\);
    
    \line5[27]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[27]_net_1\);
    
    \line3[45]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[45]_net_1\);
    
    \line6[38]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[38]_net_1\);
    
    \raddr_pos_RNIBUI17[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1633, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[10]\, D => N_1409, Y => N_1697);
    
    \line6_RNI3IAG[1]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[1]_net_1\, B => \line7[1]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[1]\);
    
    \line1[34]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[34]_net_1\);
    
    \line3[19]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[19]_net_1\);
    
    \line7[57]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[57]_net_1\);
    
    \line4_RNIL2UE2[63]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[31]\, C => \line5[63]_net_1\, D => 
        \line4[63]_net_1\, Y => N_1430);
    
    \line2_RNIIEFO1[35]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[3]\, 
        C => \line3[35]_net_1\, D => \line2[35]_net_1\, Y => 
        N_1146);
    
    \line4[28]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[28]_net_1\);
    
    \line1[31]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[31]_net_1\);
    
    \line5[58]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[58]_net_1\);
    
    \line4[10]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[10]_net_1\);
    
    \line4_RNIG4GB1[27]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[27]_net_1\, B => \line4[27]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[27]\);
    
    \line2[56]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[56]_net_1\);
    
    \line5[47]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[47]_net_1\);
    
    \line0_RNIVP271[24]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[24]_net_1\, B => \line0[24]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_7_1_1[24]\);
    
    \line4[3]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[3]_net_1\);
    
    \line2_RNI7UGH[12]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[12]_net_1\, B => \line2[12]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[12]\);
    
    raddr_pos_0_rep1 : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_0_rep1\);
    
    \line6[26]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[26]_net_1\);
    
    \line5_or[32]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line5_0, B => sha256_system_sb_0_GPIO_9_M2F, 
        Y => \line5_or[32]_net_1\);
    
    \line0[26]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[26]_net_1\);
    
    \line1[15]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[15]_net_1\);
    
    \line6[49]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[49]_net_1\);
    
    \line6[13]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[13]_net_1\);
    
    \line1[63]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[63]_net_1\);
    
    \raddr_pos_RNIMQJB8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1648, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[25]\, D => N_1424, Y => N_1712);
    
    \line4_RNIG84F1[35]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[3]\, C => \line5[35]_net_1\, D => 
        \line4[35]_net_1\, Y => N_1402);
    
    \line2[54]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[54]_net_1\);
    
    \line2[26]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[26]_net_1\);
    
    \line6_RNI5VN61[48]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[16]\, C => \line7[48]_net_1\, D => 
        \line6[48]_net_1\, Y => N_1639);
    
    \line2_RNI3ARN[24]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[24]_net_1\, B => \line2[24]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_14_1_1[24]\);
    
    \line4[47]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[47]_net_1\);
    
    \raddr_pos_RNI9S144[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_944, 
        D => N_1168, Y => \data_out_31_1_1[25]\);
    
    \line6[24]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[24]_net_1\);
    
    \line4_RNI2KH81[13]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[13]_net_1\, B => \line4[13]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[13]\);
    
    \line0_RNI2AA32[33]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[1]\, 
        C => \line1[33]_net_1\, D => \line0[33]_net_1\, Y => 
        N_920);
    
    data_available : SLE
      port map(D => N_12_0_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SHA256_Module_0_data_available\);
    
    \line0[24]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[24]_net_1\);
    
    \line4_RNI7EUB[5]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[5]_net_1\, B => \line5[5]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[5]\);
    
    \line2[51]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[51]_net_1\);
    
    \line7[23]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[23]_net_1\);
    
    \raddr_pos_RNIHR1A3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_930, 
        D => N_1154, Y => \data_out_31_1_1[11]\);
    
    \line6[21]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[21]_net_1\);
    
    \line4[37]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[37]_net_1\);
    
    \line2[37]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[37]_net_1\);
    
    \line4[56]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[56]_net_1\);
    
    \line2[24]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[24]_net_1\);
    
    \line0[21]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[21]_net_1\);
    
    \line7[9]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[9]_net_1\);
    
    \line7[43]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[43]_net_1\);
    
    \line0_RNIRAES1[45]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[13]\, 
        C => \line1[45]_net_1\, D => \line0[45]_net_1\, Y => 
        N_932);
    
    \line6_RNI5KAG[2]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[2]_net_1\, B => \line7[2]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[2]\);
    
    \line6[59]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[59]_net_1\);
    
    \line0_RNIJA652[37]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[5]\, 
        C => \line1[37]_net_1\, D => \line0[37]_net_1\, Y => 
        N_924);
    
    \line5[12]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[12]_net_1\);
    
    \line2_RNIR6BQ1[37]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[5]\, 
        C => \line3[37]_net_1\, D => \line2[37]_net_1\, Y => 
        N_1148);
    
    \line2_or[32]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line2_0, B => sha256_system_sb_0_GPIO_9_M2F, 
        Y => \line2_or[32]_net_1\);
    
    \line6_RNIHJBG1[59]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[27]\, C => \line7[59]_net_1\, D => 
        \line6[59]_net_1\, Y => N_1650);
    
    \raddr_pos_RNI367B3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_936, 
        D => N_1160, Y => \data_out_31_1_1[17]\);
    
    \line2[21]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[21]_net_1\);
    
    \line0[17]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[17]_net_1\);
    
    \line2_RNII2DA1[56]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[24]\, C => \line3[56]_net_1\, D => 
        \line2[56]_net_1\, Y => N_1167);
    
    \line1[55]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[55]_net_1\);
    
    \line3[35]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[35]_net_1\);
    
    \line6_RNIC6N61[42]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[10]\, C => \line7[42]_net_1\, D => 
        \line6[42]_net_1\, Y => N_1633);
    
    \line4[54]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[54]_net_1\);
    
    \line0[55]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[55]_net_1\);
    
    \line5[3]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[3]_net_1\);
    
    \line7[36]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[36]_net_1\);
    
    \line6[18]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[18]_net_1\);
    
    raddr_pos_1_rep1 : SLE
      port map(D => sha256_controller_0_read_addr_0(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_1_rep1\);
    
    \line6_RNIPIN61[45]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[13]\, C => \line7[45]_net_1\, D => 
        \line6[45]_net_1\, Y => N_1636);
    
    \line6_RNIEE8S[24]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[24]_net_1\, B => \line6[24]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[24]\);
    
    \line4[51]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[51]_net_1\);
    
    \raddr_pos_RNIR8AG4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_925, 
        D => N_1149, Y => \data_out_31_1_1[6]\);
    
    \line4_RNIJM852[50]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[18]\, C => \line5[50]_net_1\, D => 
        \line4[50]_net_1\, Y => N_1417);
    
    \raddr_pos_fast_fast[0]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_fast_fast[0]_net_1\);
    
    \line5[30]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[30]_net_1\);
    
    \line0_RNIEMA32[36]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[4]\, 
        C => \line1[36]_net_1\, D => \line0[36]_net_1\, Y => 
        N_923);
    
    \line2_RNIJRVT[49]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[17]\, C => \line3[49]_net_1\, D => 
        \line2[49]_net_1\, Y => N_1160);
    
    \line7[34]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[34]_net_1\);
    
    \line7[28]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[28]_net_1\);
    
    \line4_RNI1BQE2[57]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[25]\, C => \line5[57]_net_1\, D => 
        \line4[57]_net_1\, Y => N_1424);
    
    \line6[61]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[61]_net_1\);
    
    \raddr_pos_RNICOBU6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1634, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[11]\, D => N_1410, Y => N_1698);
    
    \line2_RNI5SGH[11]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[11]_net_1\, B => \line2[11]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[11]\);
    
    \raddr_pos[0]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos[0]_net_1\);
    
    \line7[48]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[48]_net_1\);
    
    \line2_RNISU2I[14]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[14]_net_1\, B => \line2[14]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[14]\);
    
    \line3[59]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[59]_net_1\);
    
    \line7[31]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[31]_net_1\);
    
    \line2[15]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[15]_net_1\);
    
    \line4_RNI5CUB[4]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[4]_net_1\, B => \line5[4]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[4]\);
    
    \line2[42]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[42]_net_1\);
    
    \raddr_pos_RNIRGT34[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_927, 
        D => N_1151, Y => \data_out_31_1_1[8]\);
    
    \line4_RNIC44F1[34]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[2]\, C => \line5[34]_net_1\, D => 
        \line4[34]_net_1\, Y => N_1401);
    
    \line2_RNI62DT[42]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[10]\, C => \line3[42]_net_1\, D => 
        \line2[42]_net_1\, Y => N_1153);
    
    \line1_or[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line1_0_62, B => 
        sha256_system_sb_0_GPIO_9_M2F, Y => \line1_or[0]_net_1\);
    
    \line3[22]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[22]_net_1\);
    
    \line0_RNIMCA11[13]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[13]_net_1\, B => \line0[13]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[13]\);
    
    \line5[0]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[0]_net_1\);
    
    \line6_RNITMN61[46]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[14]\, C => \line7[46]_net_1\, D => 
        \line6[46]_net_1\, Y => N_1637);
    
    \line4_RNISU282[47]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[15]\, C => \line5[47]_net_1\, D => 
        \line4[47]_net_1\, Y => N_1414);
    
    \line4_RNIVASE2[61]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[29]\, C => \line5[61]_net_1\, D => 
        \line4[61]_net_1\, Y => N_1428);
    
    \line3[17]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[17]_net_1\);
    
    \line6_RNIS8941[36]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[4]\, C => \line7[36]_net_1\, D => 
        \line6[36]_net_1\, Y => N_1627);
    
    \line4_RNI13752[49]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[17]\, C => \line5[49]_net_1\, D => 
        \line4[49]_net_1\, Y => N_1416);
    
    \line4_RNI4S3F1[32]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[0]\, C => \line5[32]_net_1\, D => 
        \line4[32]_net_1\, Y => N_1399);
    
    \line6[36]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[36]_net_1\);
    
    \line0[42]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[42]_net_1\);
    
    \line2[5]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[5]_net_1\);
    
    \raddr_pos_RNIMRKB8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1650, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[27]\, D => N_1426, Y => N_1714);
    
    \line1[39]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[39]_net_1\);
    
    \line5[13]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[13]_net_1\);
    
    \line6_RNITM9N[8]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line7[8]_net_1\, B => \line6[8]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_29_1_1[8]\);
    
    \line4[26]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[26]_net_1\);
    
    \line4[15]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[15]_net_1\);
    
    m35 : CFG4
      generic map(INIT => x"4C08")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_30, Y => 
        line0_0);
    
    \line4_RNILM652[46]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[14]\, C => \line5[46]_net_1\, D => 
        \line4[46]_net_1\, Y => N_1413);
    
    \line5[56]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[56]_net_1\);
    
    \raddr_pos_RNIL1PK7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1645, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[22]\, D => N_1421, Y => N_1709);
    
    \line6_RNI4H941[38]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[6]\, C => \line7[38]_net_1\, D => 
        \line6[38]_net_1\, Y => N_1629);
    
    \line2_RNI18RN[23]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[23]_net_1\, B => \line2[23]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_14_1_1[23]\);
    
    \line6[47]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[47]_net_1\);
    
    \line6[34]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[34]_net_1\);
    
    \line2[62]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[62]_net_1\);
    
    \line0_RNI72371[28]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[28]_net_1\, B => \line0[28]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_7_1_1[28]\);
    
    \line0_RNI0NA11[18]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[18]_net_1\, B => \line0[18]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[18]\);
    
    m38 : CFG4
      generic map(INIT => x"8F07")

      port map(A => waddr_in_net_0(3), B => waddr_in_net_0(2), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_13_0, Y => N_39);
    
    m1 : CFG2
      generic map(INIT => x"8")

      port map(A => sha256_system_sb_0_GPIO_9_M2F, B => 
        sha256_system_sb_0_GPIO_1_M2F, Y => 
        data_out_ready_0_sqmuxa);
    
    \line1[1]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[1]_net_1\);
    
    \line6[31]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[31]_net_1\);
    
    \line4[24]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[24]_net_1\);
    
    \line5[54]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[54]_net_1\);
    
    \line6_RNIDSAG[6]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[6]_net_1\, B => \line7[6]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[6]\);
    
    \line1[20]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[20]_net_1\);
    
    \line1[42]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[42]_net_1\);
    
    \line4[21]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[21]_net_1\);
    
    \line2[59]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[59]_net_1\);
    
    \raddr_pos_fast[0]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_fast[0]_net_1\);
    
    \line5[51]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[51]_net_1\);
    
    \line6[57]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[57]_net_1\);
    
    \line7[8]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[8]_net_1\);
    
    \raddr_pos_RNIRT6B3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_935, 
        D => N_1159, Y => \data_out_31_1_1[16]\);
    
    \line0[3]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[3]_net_1\);
    
    \line6[29]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[29]_net_1\);
    
    \line0[29]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[29]_net_1\);
    
    \line6_RNIGAN61[43]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[11]\, C => \line7[43]_net_1\, D => 
        \line6[43]_net_1\, Y => N_1634);
    
    \raddr_pos_RNIG3J07[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1632, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[9]\, D => N_1408, Y => N_1696);
    
    \line3[42]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[42]_net_1\);
    
    \line5[18]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[18]_net_1\);
    
    \line4_RNI9GUB[6]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[6]_net_1\, B => \line5[6]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[6]\);
    
    \line2[43]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[43]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line2_RNI7ERN[26]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[26]_net_1\, B => \line2[26]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_14_1_1[26]\);
    
    \line2[29]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[29]_net_1\);
    
    \line6_RNI7MAG[3]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[3]_net_1\, B => \line7[3]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[3]\);
    
    \line0[30]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[30]_net_1\);
    
    \line3[23]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[23]_net_1\);
    
    \line7[62]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[62]_net_1\);
    
    \line1[5]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[5]_net_1\);
    
    \line4_RNI13IF1[41]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_22_1_1[9]\, 
        C => \line5[41]_net_1\, D => \line4[41]_net_1\, Y => 
        N_1408);
    
    \raddr_pos_RNI1K144[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_943, 
        D => N_1167, Y => \data_out_31_1_1[24]\);
    
    \line6[16]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[16]_net_1\);
    
    \line0[9]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[9]_net_1\);
    
    \line6_RNI8AAS[30]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[30]_net_1\, B => \line6[30]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[30]\);
    
    \line0[4]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[4]_net_1\);
    
    \line0[43]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[43]_net_1\);
    
    \line5[2]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[2]_net_1\);
    
    \line4[59]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[59]_net_1\);
    
    raddr_pos_0_rep2 : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_0_rep2\);
    
    \line3_or[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line3_0_62, B => 
        sha256_system_sb_0_GPIO_9_M2F, Y => \line3_or[0]_net_1\);
    
    m25 : CFG4
      generic map(INIT => x"8C04")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_23_0, Y => 
        line3_0);
    
    \line4_RNI8SFB1[23]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[23]_net_1\, B => \line4[23]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[23]\);
    
    \line7[10]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[10]_net_1\);
    
    \line5[20]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[20]_net_1\);
    
    \line6_RNIJGAP[19]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[19]_net_1\, B => \line6[19]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[19]\);
    
    \line1[12]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[12]_net_1\);
    
    \line6_RNIGS841[33]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[1]\, C => \line7[33]_net_1\, D => 
        \line6[33]_net_1\, Y => N_1624);
    
    \line5[35]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[35]_net_1\);
    
    \raddr_pos[1]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos[1]_net_1\);
    
    \line3[57]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[57]_net_1\);
    
    \line2_RNIEAFO1[34]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[2]\, 
        C => \line3[34]_net_1\, D => \line2[34]_net_1\, Y => 
        N_1145);
    
    \line6[3]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[3]_net_1\);
    
    \line4_RNI9OQ41[15]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[15]_net_1\, B => \line5[15]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[15]\);
    
    \line0[5]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[5]_net_1\);
    
    m28 : CFG4
      generic map(INIT => x"4C08")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_23_0, Y => 
        line2_0);
    
    \line7[26]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[26]_net_1\);
    
    \line6[14]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[14]_net_1\);
    
    \line2[63]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[63]_net_1\);
    
    \line2_RNIN2BQ1[36]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[4]\, 
        C => \line3[36]_net_1\, D => \line2[36]_net_1\, Y => 
        N_1147);
    
    \line2_RNI60LC1[1]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[1]_net_1\, B => \line2[1]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[1]\);
    
    \line0[2]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[2]_net_1\);
    
    \line7[50]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[50]_net_1\);
    
    \line4_RNICE652[44]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[12]\, C => \line5[44]_net_1\, D => 
        \line4[44]_net_1\, Y => N_1411);
    
    \line2_RNI62FO1[32]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[0]\, 
        C => \line3[32]_net_1\, D => \line2[32]_net_1\, Y => 
        N_1143);
    
    \line7[46]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[46]_net_1\);
    
    \line7[39]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[39]_net_1\);
    
    \line6[11]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[11]_net_1\);
    
    \line1[61]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[61]_net_1\);
    
    \line5[40]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[40]_net_1\);
    
    \line2[48]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[48]_net_1\);
    
    \line3[62]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[62]_net_1\);
    
    \line7[24]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[24]_net_1\);
    
    \line3[28]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[28]_net_1\);
    
    \line1[43]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[43]_net_1\);
    
    \line2_RNIL6FA1[61]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[29]\, C => \line3[61]_net_1\, D => 
        \line2[61]_net_1\, Y => N_1172);
    
    \line0_RNI1S271[25]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[25]_net_1\, B => \line0[25]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_7_1_1[25]\);
    
    \line7[44]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[44]_net_1\);
    
    \line4[62]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[62]_net_1\);
    
    \line1[37]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[37]_net_1\);
    
    \raddr_pos_RNI3PT34[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_928, 
        D => N_1152, Y => \data_out_31_1_1[9]\);
    
    \line6_RNICO841[32]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[0]\, C => \line7[32]_net_1\, D => 
        \line6[32]_net_1\, Y => N_1623);
    
    \line7[21]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[21]_net_1\);
    
    \line0[48]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[48]_net_1\);
    
    \raddr_pos_RNI78JP3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_941, 
        D => N_1165, Y => \data_out_31_1_1[22]\);
    
    \line1[52]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[52]_net_1\);
    
    \line4[40]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[40]_net_1\);
    
    \line3[32]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[32]_net_1\);
    
    \line0_RNIPL471[30]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[30]_net_1\, B => \line0[30]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_7_1_1[30]\);
    
    \line7[41]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[41]_net_1\);
    
    \line4_RNIAUFB1[24]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[24]_net_1\, B => \line4[24]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[24]\);
    
    \line0[52]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[52]_net_1\);
    
    \line6_RNI9VM41[41]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_29_1_1[9]\, 
        C => \line7[41]_net_1\, D => \line6[41]_net_1\, Y => 
        N_1632);
    
    \line4_or[32]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line4_0, B => sha256_system_sb_0_GPIO_9_M2F, 
        Y => \line4_or[32]_net_1\);
    
    \line2_RNIS63U[52]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[20]\, C => \line3[52]_net_1\, D => 
        \line2[52]_net_1\, Y => N_1163);
    
    \line3[43]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[43]_net_1\);
    
    \line0_RNIBMK01[7]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[7]_net_1\, B => \line0[7]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[7]\);
    
    \line4_RNIE2GB1[26]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[26]_net_1\, B => \line4[26]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[26]\);
    
    raddr_pos_1_rep2 : SLE
      port map(D => sha256_controller_0_read_addr_0(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_1_rep2\);
    
    \line4[30]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[30]_net_1\);
    
    \raddr_pos_RNI7DAB3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_937, 
        D => N_1161, Y => \data_out_31_1_1[18]\);
    
    \line6_RNICC8S[23]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[23]_net_1\, B => \line6[23]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[23]\);
    
    \line2[30]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[30]_net_1\);
    
    \raddr_pos_RNIGKIV6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1640, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[17]\, D => N_1416, Y => N_1704);
    
    \line1[6]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[6]_net_1\);
    
    \line0_RNI4U852[63]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[31]\, C => \line1[63]_net_1\, D => 
        \line0[63]_net_1\, Y => N_950);
    
    \raddr_pos_RNI2I007[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1644, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[21]\, D => N_1420, Y => N_1708);
    
    \line0_RNI3EO01[12]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[12]_net_1\, B => \line0[12]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[12]\);
    
    \line7[63]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[63]_net_1\);
    
    \line4_RNIPATI[8]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line5[8]_net_1\, B => \line4[8]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_22_1_1[8]\);
    
    \line4_RNITU652[48]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[16]\, C => \line5[48]_net_1\, D => 
        \line4[48]_net_1\, Y => N_1415);
    
    \line6[39]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[39]_net_1\);
    
    \line0[10]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[10]_net_1\);
    
    \line4[5]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[5]_net_1\);
    
    \line2_RNI3QGH[10]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[10]_net_1\, B => \line2[10]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[10]\);
    
    \line0_RNIIAC11[20]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[20]_net_1\, B => \line0[20]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[20]\);
    
    \line2[57]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[57]_net_1\);
    
    \line2[0]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[0]_net_1\);
    
    \line1[25]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[25]_net_1\);
    
    \line4[2]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[2]_net_1\);
    
    \line6[27]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[27]_net_1\);
    
    \line4[29]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[29]_net_1\);
    
    \line1[48]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[48]_net_1\);
    
    \line1[13]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[13]_net_1\);
    
    \line2[12]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[12]_net_1\);
    
    \line0[27]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[27]_net_1\);
    
    \line5[59]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[59]_net_1\);
    
    \line0_RNI1CO01[11]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[11]_net_1\, B => \line0[11]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[11]\);
    
    m31 : CFG4
      generic map(INIT => x"2301")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_30, Y => 
        line1_0_62);
    
    \line2_RNI033I[16]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[16]_net_1\, B => \line2[16]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[16]\);
    
    m17 : CFG4
      generic map(INIT => x"8C04")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_15_0, Y => 
        line5_0);
    
    \line2[27]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[27]_net_1\);
    
    \line2_RNIVABQ1[38]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[6]\, 
        C => \line3[38]_net_1\, D => \line2[38]_net_1\, Y => 
        N_1149);
    
    \line3[48]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[48]_net_1\);
    
    \line4_RNIP2QE2[55]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[23]\, C => \line5[55]_net_1\, D => 
        \line4[55]_net_1\, Y => N_1422);
    
    \line6[7]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[7]_net_1\);
    
    \raddr_pos_RNI356B3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_932, 
        D => N_1156, Y => \data_out_31_1_1[13]\);
    
    \line5[16]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[16]_net_1\);
    
    \line4_RNIUFH81[11]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[11]_net_1\, B => \line4[11]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[11]\);
    
    \line3_or[32]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line3_0, B => sha256_system_sb_0_GPIO_9_M2F, 
        Y => \line3_or[32]_net_1\);
    
    \line0[35]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[35]_net_1\);
    
    \line6_RNIHER61[52]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[20]\, C => \line7[52]_net_1\, D => 
        \line6[52]_net_1\, Y => N_1643);
    
    \line0_RNIBRES1[49]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[17]\, 
        C => \line1[49]_net_1\, D => \line0[49]_net_1\, Y => 
        N_936);
    
    \line3[63]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[63]_net_1\);
    
    \line4[57]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[57]_net_1\);
    
    \line0_RNI94371[29]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[29]_net_1\, B => \line0[29]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_7_1_1[29]\);
    
    \line0_RNIOEA11[14]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[14]_net_1\, B => \line0[14]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[14]\);
    
    \line6_RNIJ7L41[39]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_29_1_1[7]\, 
        C => \line7[39]_net_1\, D => \line6[39]_net_1\, Y => 
        N_1630);
    
    \line4[12]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[12]_net_1\);
    
    \line0_or[32]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line0_0, B => sha256_system_sb_0_GPIO_9_M2F, 
        Y => \line0_or[32]_net_1\);
    
    \line4[63]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[63]_net_1\);
    
    \line5[14]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[14]_net_1\);
    
    \raddr_pos_RNIP32A3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_931, 
        D => N_1155, Y => \data_out_31_1_1[12]\);
    
    \line6_RNI4VJ91[47]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[15]\, C => \line7[47]_net_1\, D => 
        \line6[47]_net_1\, Y => N_1638);
    
    \line1[53]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[53]_net_1\);
    
    \line7[15]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[15]_net_1\);
    
    \line6_RNI13BG1[55]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[23]\, C => \line7[55]_net_1\, D => 
        \line6[55]_net_1\, Y => N_1646);
    
    \line4_RNI3AUB[3]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[3]_net_1\, B => \line5[3]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[3]\);
    
    \line3[33]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[33]_net_1\);
    
    \line5[25]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[25]_net_1\);
    
    \line0_or[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => line0_0_62, B => 
        sha256_system_sb_0_GPIO_9_M2F, Y => \line0_or[0]_net_1\);
    
    \line3[10]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[10]_net_1\);
    
    \line0[53]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[53]_net_1\);
    
    \line7[2]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[2]_net_1\);
    
    \line1[18]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[18]_net_1\);
    
    \line5[11]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[11]_net_1\);
    
    \raddr_pos_RNIUM4C7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1629, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[6]\, D => N_1405, Y => N_1693);
    
    \raddr_pos_RNIC5C87[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1626, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[3]\, D => N_1402, Y => N_1690);
    
    \line7[37]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[37]_net_1\);
    
    \line4_RNI0IH81[12]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[12]_net_1\, B => \line4[12]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[12]\);
    
    \line6_RNIDFBG1[58]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[26]\, C => \line7[58]_net_1\, D => 
        \line6[58]_net_1\, Y => N_1649);
    
    \line2_RNIUEDA1[59]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[27]\, C => \line3[59]_net_1\, D => 
        \line2[59]_net_1\, Y => N_1170);
    
    \line7[55]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[55]_net_1\);
    
    \line0_RNIDO3V1[42]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_7_1_1[10]\, C => \line1[42]_net_1\, D => 
        \line0[42]_net_1\, Y => N_929);
    
    \line1[3]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[3]_net_1\);
    
    \line2_RNI9GRN[27]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[27]_net_1\, B => \line2[27]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_14_1_1[27]\);
    
    \line5[45]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[45]_net_1\);
    
    \line6[19]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[19]_net_1\);
    
    \line6[40]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[40]_net_1\);
    
    \line2[46]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[46]_net_1\);
    
    \line0_RNIBC4A1[5]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[5]_net_1\, B => \line0[5]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[5]\);
    
    \raddr_pos[2]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_3_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \raddr_pos_2\);
    
    \line0_RNISIA11[16]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[16]_net_1\, B => \line0[16]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[16]\);
    
    \line3[3]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[3]_net_1\);
    
    \line3[26]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[26]_net_1\);
    
    \line6_RNI93O61[49]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[17]\, C => \line7[49]_net_1\, D => 
        \line6[49]_net_1\, Y => N_1640);
    
    m9 : CFG4
      generic map(INIT => x"08FF")

      port map(A => AHB_slave_dummy_0_write_en, B => N_49, C => 
        sha256_system_sb_0_GPIO_1_M2F, D => 
        sha256_system_sb_0_GPIO_9_M2F, Y => N_49_mux);
    
    \line6_RNI96AP[14]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[14]_net_1\, B => \line6[14]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[14]\);
    
    \line2[13]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[13]_net_1\);
    
    \line7[29]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[29]_net_1\);
    
    \line4[45]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[45]_net_1\);
    
    \line1[58]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[58]_net_1\);
    
    \line0[46]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[46]_net_1\);
    
    \line0[60]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[60]_net_1\);
    
    \line3[38]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[38]_net_1\);
    
    \line2[44]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[44]_net_1\);
    
    \line6_RNI76CP[22]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[22]_net_1\, B => \line6[22]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[22]\);
    
    \line7[49]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line7_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line7[49]_net_1\);
    
    \line0[58]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[58]_net_1\);
    
    \line4_RNIC0GB1[25]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[25]_net_1\, B => \line4[25]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[25]\);
    
    \line0[7]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[7]_net_1\);
    
    \line6[50]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[50]_net_1\);
    
    \line3[24]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[24]_net_1\);
    
    \line6_RNIVQP61[51]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[19]\, C => \line7[51]_net_1\, D => 
        \line6[51]_net_1\, Y => N_1642);
    
    \line4[35]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[35]_net_1\);
    
    \line6[9]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[9]_net_1\);
    
    \line2[41]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[41]_net_1\);
    
    \line2[35]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[35]_net_1\);
    
    \line0_RNI7NES1[48]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[16]\, 
        C => \line1[48]_net_1\, D => \line0[48]_net_1\, Y => 
        N_935);
    
    \line6[37]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[37]_net_1\);
    
    \raddr_pos_RNI0JI07[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1631, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[8]\, D => N_1407, Y => N_1695);
    
    \line0[44]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[44]_net_1\);
    
    \line3[21]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[21]_net_1\);
    
    \line4_RNI804F1[33]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[1]\, C => \line5[33]_net_1\, D => 
        \line4[33]_net_1\, Y => N_1400);
    
    \line5[32]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[32]_net_1\);
    
    \line4[13]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[13]_net_1\);
    
    \line2_RNIVU4K1[40]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_14_1_1[8]\, C => \line3[40]_net_1\, D => 
        \line2[40]_net_1\, Y => N_1151);
    
    \line0[15]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[15]_net_1\);
    
    \line2_RNIA6FO1[33]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[1]\, 
        C => \line3[33]_net_1\, D => \line2[33]_net_1\, Y => 
        N_1144);
    
    \line2_RNIA6DT[43]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[11]\, C => \line3[43]_net_1\, D => 
        \line2[43]_net_1\, Y => N_1154);
    
    \line4[27]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[27]_net_1\);
    
    data_out_ready_1 : CFG4
      generic map(INIT => x"CDCC")

      port map(A => N_3_0, B => data_out_ready_0_sqmuxa, C => 
        AHB_slave_dummy_0_write_en, D => 
        \SHA256_Module_0_data_out_ready\, Y => \data_out_ready_1\);
    
    \line5[6]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[6]_net_1\);
    
    \raddr_pos_RNITJ544[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos_3\, B => \raddr_pos_2\, C => N_947, 
        D => N_1171, Y => \data_out_31_1_1[28]\);
    
    \line2_RNIM6DA1[57]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[25]\, C => \line3[57]_net_1\, D => 
        \line2[57]_net_1\, Y => N_1168);
    
    \line5[57]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[57]_net_1\);
    
    \line0[41]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[41]_net_1\);
    
    \line3[6]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[6]_net_1\);
    
    \line0_RNI0I881[0]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[0]_net_1\, B => \line0[0]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[0]\);
    
    \line6_RNI0U9P[10]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[10]_net_1\, B => \line6[10]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[10]\);
    
    \line2[18]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[18]_net_1\);
    
    \line1[46]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[46]_net_1\);
    
    m41 : CFG4
      generic map(INIT => x"8C04")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_39, Y => 
        line7_0);
    
    m12 : CFG4
      generic map(INIT => x"3733")

      port map(A => sha256_system_sb_0_GPIO_1_M2F, B => 
        sha256_system_sb_0_GPIO_9_M2F, C => waddr_in_net_0(4), D
         => AHB_slave_dummy_0_write_en, Y => N_13_0);
    
    m19 : CFG4
      generic map(INIT => x"1302")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_15_0, Y => 
        line4_0_62);
    
    \line2[61]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[61]_net_1\);
    
    \line5[7]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[7]_net_1\);
    
    \line0_RNIE6S82[57]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[25]\, C => \line1[57]_net_1\, D => 
        \line0[57]_net_1\, Y => N_944);
    
    \line6[8]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line6_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line6[8]_net_1\);
    
    \line2_RNIFOGE1[5]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[5]_net_1\, B => \line2[5]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[5]\);
    
    \line2[9]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line2_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line2[9]_net_1\);
    
    \line0[1]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line0_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line0[1]_net_1\);
    
    \line3[50]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[50]_net_1\);
    
    \line3[46]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[46]_net_1\);
    
    \line5[60]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line5_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line5[60]_net_1\);
    
    \line1[44]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[44]_net_1\);
    
    \line4_RNI4QHB1[30]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[30]_net_1\, B => \line4[30]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[30]\);
    
    \raddr_pos_RNIH1007[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1643, B => \raddr_pos_3\, C => 
        \data_out_31_1_1[20]\, D => N_1419, Y => N_1707);
    
    \line0_RNITEGS1[50]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[18]\, 
        C => \line1[50]_net_1\, D => \line0[50]_net_1\, Y => 
        N_937);
    
    \line4_RNIHMA52[54]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[22]\, C => \line5[54]_net_1\, D => 
        \line4[54]_net_1\, Y => N_1421);
    
    \line1[41]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[41]_net_1\);
    
    \line4[18]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line4_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line4[18]_net_1\);
    
    m20 : CFG4
      generic map(INIT => x"4C08")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(0), C
         => sha256_system_sb_0_GPIO_9_M2F, D => N_15_0, Y => 
        line4_0);
    
    data_available_RNO : CFG4
      generic map(INIT => x"DFCE")

      port map(A => waddr_in_net_0(0), B => 
        \SHA256_Module_0_data_available\, C => 
        sha256_system_sb_0_GPIO_9_M2F, D => N_49_mux, Y => 
        N_12_0_i_0);
    
    \line3[44]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[32]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line3[44]_net_1\);
    
    \line1[4]\ : SLE
      port map(D => AHB_slave_dummy_0_mem_wdata(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line1_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT => 
        GND_net_1, Q => \line1[4]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity SHA256_BLOCK is

    port( SHA256_BLOCK_0_H0_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o            : out   std_logic_vector(31 downto 0);
          AHB_slave_dummy_0_mem_wdata    : in    std_logic_vector(31 downto 0);
          waddr_in_net_0                 : in    std_logic_vector(4 downto 0);
          state_out_net_0                : out   std_logic_vector(0 to 0);
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic;
          SHA256_Module_0_di_req_o       : out   std_logic;
          SHA256_Module_0_do_valid_o     : out   std_logic;
          SHA256_Module_0_error_o        : out   std_logic;
          SHA256_Module_0_data_out_ready : out   std_logic;
          sha256_system_sb_0_GPIO_9_M2F  : in    std_logic;
          SHA256_Module_0_data_available : out   std_logic;
          sha256_system_sb_0_GPIO_1_M2F  : in    std_logic;
          AHB_slave_dummy_0_write_en     : in    std_logic;
          ce_i_i_2_i_0                   : out   std_logic;
          N_88_i_0                       : out   std_logic;
          N_87_i_0                       : out   std_logic
        );

end SHA256_BLOCK;

architecture DEF_ARCH of SHA256_BLOCK is 

  component sha256_controller
    port( sha256_controller_0_read_addr_0 : out   std_logic_vector(3 downto 0);
          sha256_controller_0_bytes_o     : out   std_logic_vector(1 to 1);
          state_out_net_0                 : out   std_logic_vector(0 to 0);
          state_4                         : out   std_logic;
          state_3                         : out   std_logic;
          state_1                         : out   std_logic;
          ce_i_i_2                        : out   std_logic;
          ce_i_i_2_i_0                    : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK    : in    std_logic := 'U';
          sha256_system_sb_0_GPIO_9_M2F   : in    std_logic := 'U';
          sha256_controller_0_end_o       : out   std_logic;
          last_block_0                    : out   std_logic;
          N_88_i_0                        : out   std_logic;
          N_28                            : out   std_logic;
          SHA256_Module_0_di_req_o        : in    std_logic := 'U';
          N_89                            : out   std_logic;
          SHA256_Module_0_do_valid_o      : in    std_logic := 'U';
          last_block                      : in    std_logic := 'U';
          prev_sig                        : in    std_logic := 'U';
          first_block                     : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready  : in    std_logic := 'U';
          prev_sig_0                      : in    std_logic := 'U';
          N_87_i_0                        : out   std_logic
        );
  end component;

  component gv_sha256
    port( sha256_controller_0_bytes_o  : in    std_logic_vector(1 to 1) := (others => 'U');
          raddr_pos                    : in    std_logic_vector(3 downto 2) := (others => 'U');
          SHA256_BLOCK_0_H0_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o          : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o          : out   std_logic_vector(31 downto 0);
          state_2                      : in    std_logic := 'U';
          state_0                      : in    std_logic := 'U';
          state_3                      : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK : in    std_logic := 'U';
          SHA256_Module_0_di_req_o     : out   std_logic;
          SHA256_Module_0_do_valid_o   : out   std_logic;
          sha256_controller_0_end_o    : in    std_logic := 'U';
          last_block_0                 : in    std_logic := 'U';
          ce_i_i_2                     : in    std_logic := 'U';
          N_28                         : in    std_logic := 'U';
          SHA256_Module_0_error_o      : out   std_logic;
          N_1696                       : in    std_logic := 'U';
          N_1400                       : in    std_logic := 'U';
          N_1624                       : in    std_logic := 'U';
          N_920                        : in    std_logic := 'U';
          N_1144                       : in    std_logic := 'U';
          N_1399                       : in    std_logic := 'U';
          N_1623                       : in    std_logic := 'U';
          N_919                        : in    std_logic := 'U';
          N_1143                       : in    std_logic := 'U';
          N_1401                       : in    std_logic := 'U';
          N_1625                       : in    std_logic := 'U';
          N_921                        : in    std_logic := 'U';
          N_1145                       : in    std_logic := 'U';
          ren_pos                      : in    std_logic := 'U';
          N_1694                       : in    std_logic := 'U';
          N_1692                       : in    std_logic := 'U';
          N_1693                       : in    std_logic := 'U';
          N_1691                       : in    std_logic := 'U';
          N_1690                       : in    std_logic := 'U';
          N_89                         : in    std_logic := 'U';
          N_1695                       : in    std_logic := 'U';
          N_1708                       : in    std_logic := 'U';
          N_1709                       : in    std_logic := 'U';
          N_1707                       : in    std_logic := 'U';
          N_1706                       : in    std_logic := 'U';
          N_1705                       : in    std_logic := 'U';
          N_1704                       : in    std_logic := 'U';
          N_1703                       : in    std_logic := 'U';
          N_1700                       : in    std_logic := 'U';
          N_1701                       : in    std_logic := 'U';
          N_1697                       : in    std_logic := 'U';
          N_1699                       : in    std_logic := 'U';
          N_1698                       : in    std_logic := 'U';
          N_1717                       : in    std_logic := 'U';
          N_1712                       : in    std_logic := 'U';
          N_1716                       : in    std_logic := 'U';
          N_1715                       : in    std_logic := 'U';
          N_1711                       : in    std_logic := 'U';
          N_1713                       : in    std_logic := 'U';
          N_1714                       : in    std_logic := 'U';
          N_1718                       : in    std_logic := 'U';
          N_1702                       : in    std_logic := 'U';
          N_1710                       : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component limiter_1cycle_0
    port( prev_sig                     : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK : in    std_logic := 'U';
          first_block                  : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component limiter_1cycle_1
    port( prev_sig                       : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready : in    std_logic := 'U'
        );
  end component;

  component reg_17x32
    port( AHB_slave_dummy_0_mem_wdata     : in    std_logic_vector(31 downto 0) := (others => 'U');
          sha256_controller_0_read_addr_0 : in    std_logic_vector(3 downto 0) := (others => 'U');
          waddr_in_net_0                  : in    std_logic_vector(4 downto 0) := (others => 'U');
          raddr_pos_3                     : out   std_logic;
          raddr_pos_2                     : out   std_logic;
          SHA256_Module_0_data_out_ready  : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK    : in    std_logic := 'U';
          sha256_system_sb_0_GPIO_9_M2F   : in    std_logic := 'U';
          SHA256_Module_0_data_available  : out   std_logic;
          ren_pos                         : out   std_logic;
          last_block                      : out   std_logic;
          first_block                     : out   std_logic;
          N_1717                          : out   std_logic;
          N_1716                          : out   std_logic;
          N_1711                          : out   std_logic;
          N_1710                          : out   std_logic;
          N_1708                          : out   std_logic;
          N_1705                          : out   std_logic;
          N_1704                          : out   std_logic;
          N_1701                          : out   std_logic;
          N_1690                          : out   std_logic;
          N_1691                          : out   std_logic;
          N_1707                          : out   std_logic;
          N_1703                          : out   std_logic;
          N_1715                          : out   std_logic;
          N_1700                          : out   std_logic;
          N_1714                          : out   std_logic;
          N_1697                          : out   std_logic;
          N_1693                          : out   std_logic;
          N_1706                          : out   std_logic;
          N_1696                          : out   std_logic;
          N_1709                          : out   std_logic;
          N_1698                          : out   std_logic;
          N_1699                          : out   std_logic;
          N_1694                          : out   std_logic;
          N_1702                          : out   std_logic;
          N_1712                          : out   std_logic;
          N_1695                          : out   std_logic;
          N_1692                          : out   std_logic;
          N_1718                          : out   std_logic;
          N_1713                          : out   std_logic;
          N_1144                          : out   std_logic;
          N_921                           : out   std_logic;
          N_1401                          : out   std_logic;
          N_1145                          : out   std_logic;
          N_919                           : out   std_logic;
          N_1400                          : out   std_logic;
          N_1623                          : out   std_logic;
          N_920                           : out   std_logic;
          N_1143                          : out   std_logic;
          N_1624                          : out   std_logic;
          N_1625                          : out   std_logic;
          N_1399                          : out   std_logic;
          sha256_system_sb_0_GPIO_1_M2F   : in    std_logic := 'U';
          AHB_slave_dummy_0_write_en      : in    std_logic := 'U'
        );
  end component;

    signal \sha256_controller_0_bytes_o[1]\, \raddr_pos[2]\, 
        \raddr_pos[3]\, \state[3]\, \state[1]\, \state[4]\, 
        \SHA256_Module_0_di_req_o\, \SHA256_Module_0_do_valid_o\, 
        sha256_controller_0_end_o, last_block_0, ce_i_i_2, N_28, 
        N_1696, N_1400, N_1624, N_920, N_1144, N_1399, N_1623, 
        N_919, N_1143, N_1401, N_1625, N_921, N_1145, ren_pos, 
        N_1694, N_1692, N_1693, N_1691, N_1690, N_89, N_1695, 
        N_1708, N_1709, N_1707, N_1706, N_1705, N_1704, N_1703, 
        N_1700, N_1701, N_1697, N_1699, N_1698, N_1717, N_1712, 
        N_1716, N_1715, N_1711, N_1713, N_1714, N_1718, N_1702, 
        N_1710, prev_sig, first_block, prev_sig_0, 
        \SHA256_Module_0_data_out_ready\, 
        \sha256_controller_0_read_addr_0[0]\, 
        \sha256_controller_0_read_addr_0[1]\, 
        \sha256_controller_0_read_addr_0[2]\, 
        \sha256_controller_0_read_addr_0[3]\, last_block, 
        GND_net_1, VCC_net_1 : std_logic;

    for all : sha256_controller
	Use entity work.sha256_controller(DEF_ARCH);
    for all : gv_sha256
	Use entity work.gv_sha256(DEF_ARCH);
    for all : limiter_1cycle_0
	Use entity work.limiter_1cycle_0(DEF_ARCH);
    for all : limiter_1cycle_1
	Use entity work.limiter_1cycle_1(DEF_ARCH);
    for all : reg_17x32
	Use entity work.reg_17x32(DEF_ARCH);
begin 

    SHA256_Module_0_di_req_o <= \SHA256_Module_0_di_req_o\;
    SHA256_Module_0_do_valid_o <= \SHA256_Module_0_do_valid_o\;
    SHA256_Module_0_data_out_ready <= 
        \SHA256_Module_0_data_out_ready\;

    sha256_controller_0 : sha256_controller
      port map(sha256_controller_0_read_addr_0(3) => 
        \sha256_controller_0_read_addr_0[3]\, 
        sha256_controller_0_read_addr_0(2) => 
        \sha256_controller_0_read_addr_0[2]\, 
        sha256_controller_0_read_addr_0(1) => 
        \sha256_controller_0_read_addr_0[1]\, 
        sha256_controller_0_read_addr_0(0) => 
        \sha256_controller_0_read_addr_0[0]\, 
        sha256_controller_0_bytes_o(1) => 
        \sha256_controller_0_bytes_o[1]\, state_out_net_0(0) => 
        state_out_net_0(0), state_4 => \state[4]\, state_3 => 
        \state[3]\, state_1 => \state[1]\, ce_i_i_2 => ce_i_i_2, 
        ce_i_i_2_i_0 => ce_i_i_2_i_0, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, 
        sha256_system_sb_0_GPIO_9_M2F => 
        sha256_system_sb_0_GPIO_9_M2F, sha256_controller_0_end_o
         => sha256_controller_0_end_o, last_block_0 => 
        last_block_0, N_88_i_0 => N_88_i_0, N_28 => N_28, 
        SHA256_Module_0_di_req_o => \SHA256_Module_0_di_req_o\, 
        N_89 => N_89, SHA256_Module_0_do_valid_o => 
        \SHA256_Module_0_do_valid_o\, last_block => last_block, 
        prev_sig => prev_sig, first_block => first_block, 
        SHA256_Module_0_data_out_ready => 
        \SHA256_Module_0_data_out_ready\, prev_sig_0 => 
        prev_sig_0, N_87_i_0 => N_87_i_0);
    
    gv_sha256_0 : gv_sha256
      port map(sha256_controller_0_bytes_o(1) => 
        \sha256_controller_0_bytes_o[1]\, raddr_pos(3) => 
        \raddr_pos[3]\, raddr_pos(2) => \raddr_pos[2]\, 
        SHA256_BLOCK_0_H0_o(31) => SHA256_BLOCK_0_H0_o(31), 
        SHA256_BLOCK_0_H0_o(30) => SHA256_BLOCK_0_H0_o(30), 
        SHA256_BLOCK_0_H0_o(29) => SHA256_BLOCK_0_H0_o(29), 
        SHA256_BLOCK_0_H0_o(28) => SHA256_BLOCK_0_H0_o(28), 
        SHA256_BLOCK_0_H0_o(27) => SHA256_BLOCK_0_H0_o(27), 
        SHA256_BLOCK_0_H0_o(26) => SHA256_BLOCK_0_H0_o(26), 
        SHA256_BLOCK_0_H0_o(25) => SHA256_BLOCK_0_H0_o(25), 
        SHA256_BLOCK_0_H0_o(24) => SHA256_BLOCK_0_H0_o(24), 
        SHA256_BLOCK_0_H0_o(23) => SHA256_BLOCK_0_H0_o(23), 
        SHA256_BLOCK_0_H0_o(22) => SHA256_BLOCK_0_H0_o(22), 
        SHA256_BLOCK_0_H0_o(21) => SHA256_BLOCK_0_H0_o(21), 
        SHA256_BLOCK_0_H0_o(20) => SHA256_BLOCK_0_H0_o(20), 
        SHA256_BLOCK_0_H0_o(19) => SHA256_BLOCK_0_H0_o(19), 
        SHA256_BLOCK_0_H0_o(18) => SHA256_BLOCK_0_H0_o(18), 
        SHA256_BLOCK_0_H0_o(17) => SHA256_BLOCK_0_H0_o(17), 
        SHA256_BLOCK_0_H0_o(16) => SHA256_BLOCK_0_H0_o(16), 
        SHA256_BLOCK_0_H0_o(15) => SHA256_BLOCK_0_H0_o(15), 
        SHA256_BLOCK_0_H0_o(14) => SHA256_BLOCK_0_H0_o(14), 
        SHA256_BLOCK_0_H0_o(13) => SHA256_BLOCK_0_H0_o(13), 
        SHA256_BLOCK_0_H0_o(12) => SHA256_BLOCK_0_H0_o(12), 
        SHA256_BLOCK_0_H0_o(11) => SHA256_BLOCK_0_H0_o(11), 
        SHA256_BLOCK_0_H0_o(10) => SHA256_BLOCK_0_H0_o(10), 
        SHA256_BLOCK_0_H0_o(9) => SHA256_BLOCK_0_H0_o(9), 
        SHA256_BLOCK_0_H0_o(8) => SHA256_BLOCK_0_H0_o(8), 
        SHA256_BLOCK_0_H0_o(7) => SHA256_BLOCK_0_H0_o(7), 
        SHA256_BLOCK_0_H0_o(6) => SHA256_BLOCK_0_H0_o(6), 
        SHA256_BLOCK_0_H0_o(5) => SHA256_BLOCK_0_H0_o(5), 
        SHA256_BLOCK_0_H0_o(4) => SHA256_BLOCK_0_H0_o(4), 
        SHA256_BLOCK_0_H0_o(3) => SHA256_BLOCK_0_H0_o(3), 
        SHA256_BLOCK_0_H0_o(2) => SHA256_BLOCK_0_H0_o(2), 
        SHA256_BLOCK_0_H0_o(1) => SHA256_BLOCK_0_H0_o(1), 
        SHA256_BLOCK_0_H0_o(0) => SHA256_BLOCK_0_H0_o(0), 
        SHA256_BLOCK_0_H1_o(31) => SHA256_BLOCK_0_H1_o(31), 
        SHA256_BLOCK_0_H1_o(30) => SHA256_BLOCK_0_H1_o(30), 
        SHA256_BLOCK_0_H1_o(29) => SHA256_BLOCK_0_H1_o(29), 
        SHA256_BLOCK_0_H1_o(28) => SHA256_BLOCK_0_H1_o(28), 
        SHA256_BLOCK_0_H1_o(27) => SHA256_BLOCK_0_H1_o(27), 
        SHA256_BLOCK_0_H1_o(26) => SHA256_BLOCK_0_H1_o(26), 
        SHA256_BLOCK_0_H1_o(25) => SHA256_BLOCK_0_H1_o(25), 
        SHA256_BLOCK_0_H1_o(24) => SHA256_BLOCK_0_H1_o(24), 
        SHA256_BLOCK_0_H1_o(23) => SHA256_BLOCK_0_H1_o(23), 
        SHA256_BLOCK_0_H1_o(22) => SHA256_BLOCK_0_H1_o(22), 
        SHA256_BLOCK_0_H1_o(21) => SHA256_BLOCK_0_H1_o(21), 
        SHA256_BLOCK_0_H1_o(20) => SHA256_BLOCK_0_H1_o(20), 
        SHA256_BLOCK_0_H1_o(19) => SHA256_BLOCK_0_H1_o(19), 
        SHA256_BLOCK_0_H1_o(18) => SHA256_BLOCK_0_H1_o(18), 
        SHA256_BLOCK_0_H1_o(17) => SHA256_BLOCK_0_H1_o(17), 
        SHA256_BLOCK_0_H1_o(16) => SHA256_BLOCK_0_H1_o(16), 
        SHA256_BLOCK_0_H1_o(15) => SHA256_BLOCK_0_H1_o(15), 
        SHA256_BLOCK_0_H1_o(14) => SHA256_BLOCK_0_H1_o(14), 
        SHA256_BLOCK_0_H1_o(13) => SHA256_BLOCK_0_H1_o(13), 
        SHA256_BLOCK_0_H1_o(12) => SHA256_BLOCK_0_H1_o(12), 
        SHA256_BLOCK_0_H1_o(11) => SHA256_BLOCK_0_H1_o(11), 
        SHA256_BLOCK_0_H1_o(10) => SHA256_BLOCK_0_H1_o(10), 
        SHA256_BLOCK_0_H1_o(9) => SHA256_BLOCK_0_H1_o(9), 
        SHA256_BLOCK_0_H1_o(8) => SHA256_BLOCK_0_H1_o(8), 
        SHA256_BLOCK_0_H1_o(7) => SHA256_BLOCK_0_H1_o(7), 
        SHA256_BLOCK_0_H1_o(6) => SHA256_BLOCK_0_H1_o(6), 
        SHA256_BLOCK_0_H1_o(5) => SHA256_BLOCK_0_H1_o(5), 
        SHA256_BLOCK_0_H1_o(4) => SHA256_BLOCK_0_H1_o(4), 
        SHA256_BLOCK_0_H1_o(3) => SHA256_BLOCK_0_H1_o(3), 
        SHA256_BLOCK_0_H1_o(2) => SHA256_BLOCK_0_H1_o(2), 
        SHA256_BLOCK_0_H1_o(1) => SHA256_BLOCK_0_H1_o(1), 
        SHA256_BLOCK_0_H1_o(0) => SHA256_BLOCK_0_H1_o(0), 
        SHA256_BLOCK_0_H2_o(31) => SHA256_BLOCK_0_H2_o(31), 
        SHA256_BLOCK_0_H2_o(30) => SHA256_BLOCK_0_H2_o(30), 
        SHA256_BLOCK_0_H2_o(29) => SHA256_BLOCK_0_H2_o(29), 
        SHA256_BLOCK_0_H2_o(28) => SHA256_BLOCK_0_H2_o(28), 
        SHA256_BLOCK_0_H2_o(27) => SHA256_BLOCK_0_H2_o(27), 
        SHA256_BLOCK_0_H2_o(26) => SHA256_BLOCK_0_H2_o(26), 
        SHA256_BLOCK_0_H2_o(25) => SHA256_BLOCK_0_H2_o(25), 
        SHA256_BLOCK_0_H2_o(24) => SHA256_BLOCK_0_H2_o(24), 
        SHA256_BLOCK_0_H2_o(23) => SHA256_BLOCK_0_H2_o(23), 
        SHA256_BLOCK_0_H2_o(22) => SHA256_BLOCK_0_H2_o(22), 
        SHA256_BLOCK_0_H2_o(21) => SHA256_BLOCK_0_H2_o(21), 
        SHA256_BLOCK_0_H2_o(20) => SHA256_BLOCK_0_H2_o(20), 
        SHA256_BLOCK_0_H2_o(19) => SHA256_BLOCK_0_H2_o(19), 
        SHA256_BLOCK_0_H2_o(18) => SHA256_BLOCK_0_H2_o(18), 
        SHA256_BLOCK_0_H2_o(17) => SHA256_BLOCK_0_H2_o(17), 
        SHA256_BLOCK_0_H2_o(16) => SHA256_BLOCK_0_H2_o(16), 
        SHA256_BLOCK_0_H2_o(15) => SHA256_BLOCK_0_H2_o(15), 
        SHA256_BLOCK_0_H2_o(14) => SHA256_BLOCK_0_H2_o(14), 
        SHA256_BLOCK_0_H2_o(13) => SHA256_BLOCK_0_H2_o(13), 
        SHA256_BLOCK_0_H2_o(12) => SHA256_BLOCK_0_H2_o(12), 
        SHA256_BLOCK_0_H2_o(11) => SHA256_BLOCK_0_H2_o(11), 
        SHA256_BLOCK_0_H2_o(10) => SHA256_BLOCK_0_H2_o(10), 
        SHA256_BLOCK_0_H2_o(9) => SHA256_BLOCK_0_H2_o(9), 
        SHA256_BLOCK_0_H2_o(8) => SHA256_BLOCK_0_H2_o(8), 
        SHA256_BLOCK_0_H2_o(7) => SHA256_BLOCK_0_H2_o(7), 
        SHA256_BLOCK_0_H2_o(6) => SHA256_BLOCK_0_H2_o(6), 
        SHA256_BLOCK_0_H2_o(5) => SHA256_BLOCK_0_H2_o(5), 
        SHA256_BLOCK_0_H2_o(4) => SHA256_BLOCK_0_H2_o(4), 
        SHA256_BLOCK_0_H2_o(3) => SHA256_BLOCK_0_H2_o(3), 
        SHA256_BLOCK_0_H2_o(2) => SHA256_BLOCK_0_H2_o(2), 
        SHA256_BLOCK_0_H2_o(1) => SHA256_BLOCK_0_H2_o(1), 
        SHA256_BLOCK_0_H2_o(0) => SHA256_BLOCK_0_H2_o(0), 
        SHA256_BLOCK_0_H3_o(31) => SHA256_BLOCK_0_H3_o(31), 
        SHA256_BLOCK_0_H3_o(30) => SHA256_BLOCK_0_H3_o(30), 
        SHA256_BLOCK_0_H3_o(29) => SHA256_BLOCK_0_H3_o(29), 
        SHA256_BLOCK_0_H3_o(28) => SHA256_BLOCK_0_H3_o(28), 
        SHA256_BLOCK_0_H3_o(27) => SHA256_BLOCK_0_H3_o(27), 
        SHA256_BLOCK_0_H3_o(26) => SHA256_BLOCK_0_H3_o(26), 
        SHA256_BLOCK_0_H3_o(25) => SHA256_BLOCK_0_H3_o(25), 
        SHA256_BLOCK_0_H3_o(24) => SHA256_BLOCK_0_H3_o(24), 
        SHA256_BLOCK_0_H3_o(23) => SHA256_BLOCK_0_H3_o(23), 
        SHA256_BLOCK_0_H3_o(22) => SHA256_BLOCK_0_H3_o(22), 
        SHA256_BLOCK_0_H3_o(21) => SHA256_BLOCK_0_H3_o(21), 
        SHA256_BLOCK_0_H3_o(20) => SHA256_BLOCK_0_H3_o(20), 
        SHA256_BLOCK_0_H3_o(19) => SHA256_BLOCK_0_H3_o(19), 
        SHA256_BLOCK_0_H3_o(18) => SHA256_BLOCK_0_H3_o(18), 
        SHA256_BLOCK_0_H3_o(17) => SHA256_BLOCK_0_H3_o(17), 
        SHA256_BLOCK_0_H3_o(16) => SHA256_BLOCK_0_H3_o(16), 
        SHA256_BLOCK_0_H3_o(15) => SHA256_BLOCK_0_H3_o(15), 
        SHA256_BLOCK_0_H3_o(14) => SHA256_BLOCK_0_H3_o(14), 
        SHA256_BLOCK_0_H3_o(13) => SHA256_BLOCK_0_H3_o(13), 
        SHA256_BLOCK_0_H3_o(12) => SHA256_BLOCK_0_H3_o(12), 
        SHA256_BLOCK_0_H3_o(11) => SHA256_BLOCK_0_H3_o(11), 
        SHA256_BLOCK_0_H3_o(10) => SHA256_BLOCK_0_H3_o(10), 
        SHA256_BLOCK_0_H3_o(9) => SHA256_BLOCK_0_H3_o(9), 
        SHA256_BLOCK_0_H3_o(8) => SHA256_BLOCK_0_H3_o(8), 
        SHA256_BLOCK_0_H3_o(7) => SHA256_BLOCK_0_H3_o(7), 
        SHA256_BLOCK_0_H3_o(6) => SHA256_BLOCK_0_H3_o(6), 
        SHA256_BLOCK_0_H3_o(5) => SHA256_BLOCK_0_H3_o(5), 
        SHA256_BLOCK_0_H3_o(4) => SHA256_BLOCK_0_H3_o(4), 
        SHA256_BLOCK_0_H3_o(3) => SHA256_BLOCK_0_H3_o(3), 
        SHA256_BLOCK_0_H3_o(2) => SHA256_BLOCK_0_H3_o(2), 
        SHA256_BLOCK_0_H3_o(1) => SHA256_BLOCK_0_H3_o(1), 
        SHA256_BLOCK_0_H3_o(0) => SHA256_BLOCK_0_H3_o(0), 
        SHA256_BLOCK_0_H4_o(31) => SHA256_BLOCK_0_H4_o(31), 
        SHA256_BLOCK_0_H4_o(30) => SHA256_BLOCK_0_H4_o(30), 
        SHA256_BLOCK_0_H4_o(29) => SHA256_BLOCK_0_H4_o(29), 
        SHA256_BLOCK_0_H4_o(28) => SHA256_BLOCK_0_H4_o(28), 
        SHA256_BLOCK_0_H4_o(27) => SHA256_BLOCK_0_H4_o(27), 
        SHA256_BLOCK_0_H4_o(26) => SHA256_BLOCK_0_H4_o(26), 
        SHA256_BLOCK_0_H4_o(25) => SHA256_BLOCK_0_H4_o(25), 
        SHA256_BLOCK_0_H4_o(24) => SHA256_BLOCK_0_H4_o(24), 
        SHA256_BLOCK_0_H4_o(23) => SHA256_BLOCK_0_H4_o(23), 
        SHA256_BLOCK_0_H4_o(22) => SHA256_BLOCK_0_H4_o(22), 
        SHA256_BLOCK_0_H4_o(21) => SHA256_BLOCK_0_H4_o(21), 
        SHA256_BLOCK_0_H4_o(20) => SHA256_BLOCK_0_H4_o(20), 
        SHA256_BLOCK_0_H4_o(19) => SHA256_BLOCK_0_H4_o(19), 
        SHA256_BLOCK_0_H4_o(18) => SHA256_BLOCK_0_H4_o(18), 
        SHA256_BLOCK_0_H4_o(17) => SHA256_BLOCK_0_H4_o(17), 
        SHA256_BLOCK_0_H4_o(16) => SHA256_BLOCK_0_H4_o(16), 
        SHA256_BLOCK_0_H4_o(15) => SHA256_BLOCK_0_H4_o(15), 
        SHA256_BLOCK_0_H4_o(14) => SHA256_BLOCK_0_H4_o(14), 
        SHA256_BLOCK_0_H4_o(13) => SHA256_BLOCK_0_H4_o(13), 
        SHA256_BLOCK_0_H4_o(12) => SHA256_BLOCK_0_H4_o(12), 
        SHA256_BLOCK_0_H4_o(11) => SHA256_BLOCK_0_H4_o(11), 
        SHA256_BLOCK_0_H4_o(10) => SHA256_BLOCK_0_H4_o(10), 
        SHA256_BLOCK_0_H4_o(9) => SHA256_BLOCK_0_H4_o(9), 
        SHA256_BLOCK_0_H4_o(8) => SHA256_BLOCK_0_H4_o(8), 
        SHA256_BLOCK_0_H4_o(7) => SHA256_BLOCK_0_H4_o(7), 
        SHA256_BLOCK_0_H4_o(6) => SHA256_BLOCK_0_H4_o(6), 
        SHA256_BLOCK_0_H4_o(5) => SHA256_BLOCK_0_H4_o(5), 
        SHA256_BLOCK_0_H4_o(4) => SHA256_BLOCK_0_H4_o(4), 
        SHA256_BLOCK_0_H4_o(3) => SHA256_BLOCK_0_H4_o(3), 
        SHA256_BLOCK_0_H4_o(2) => SHA256_BLOCK_0_H4_o(2), 
        SHA256_BLOCK_0_H4_o(1) => SHA256_BLOCK_0_H4_o(1), 
        SHA256_BLOCK_0_H4_o(0) => SHA256_BLOCK_0_H4_o(0), 
        SHA256_BLOCK_0_H5_o(31) => SHA256_BLOCK_0_H5_o(31), 
        SHA256_BLOCK_0_H5_o(30) => SHA256_BLOCK_0_H5_o(30), 
        SHA256_BLOCK_0_H5_o(29) => SHA256_BLOCK_0_H5_o(29), 
        SHA256_BLOCK_0_H5_o(28) => SHA256_BLOCK_0_H5_o(28), 
        SHA256_BLOCK_0_H5_o(27) => SHA256_BLOCK_0_H5_o(27), 
        SHA256_BLOCK_0_H5_o(26) => SHA256_BLOCK_0_H5_o(26), 
        SHA256_BLOCK_0_H5_o(25) => SHA256_BLOCK_0_H5_o(25), 
        SHA256_BLOCK_0_H5_o(24) => SHA256_BLOCK_0_H5_o(24), 
        SHA256_BLOCK_0_H5_o(23) => SHA256_BLOCK_0_H5_o(23), 
        SHA256_BLOCK_0_H5_o(22) => SHA256_BLOCK_0_H5_o(22), 
        SHA256_BLOCK_0_H5_o(21) => SHA256_BLOCK_0_H5_o(21), 
        SHA256_BLOCK_0_H5_o(20) => SHA256_BLOCK_0_H5_o(20), 
        SHA256_BLOCK_0_H5_o(19) => SHA256_BLOCK_0_H5_o(19), 
        SHA256_BLOCK_0_H5_o(18) => SHA256_BLOCK_0_H5_o(18), 
        SHA256_BLOCK_0_H5_o(17) => SHA256_BLOCK_0_H5_o(17), 
        SHA256_BLOCK_0_H5_o(16) => SHA256_BLOCK_0_H5_o(16), 
        SHA256_BLOCK_0_H5_o(15) => SHA256_BLOCK_0_H5_o(15), 
        SHA256_BLOCK_0_H5_o(14) => SHA256_BLOCK_0_H5_o(14), 
        SHA256_BLOCK_0_H5_o(13) => SHA256_BLOCK_0_H5_o(13), 
        SHA256_BLOCK_0_H5_o(12) => SHA256_BLOCK_0_H5_o(12), 
        SHA256_BLOCK_0_H5_o(11) => SHA256_BLOCK_0_H5_o(11), 
        SHA256_BLOCK_0_H5_o(10) => SHA256_BLOCK_0_H5_o(10), 
        SHA256_BLOCK_0_H5_o(9) => SHA256_BLOCK_0_H5_o(9), 
        SHA256_BLOCK_0_H5_o(8) => SHA256_BLOCK_0_H5_o(8), 
        SHA256_BLOCK_0_H5_o(7) => SHA256_BLOCK_0_H5_o(7), 
        SHA256_BLOCK_0_H5_o(6) => SHA256_BLOCK_0_H5_o(6), 
        SHA256_BLOCK_0_H5_o(5) => SHA256_BLOCK_0_H5_o(5), 
        SHA256_BLOCK_0_H5_o(4) => SHA256_BLOCK_0_H5_o(4), 
        SHA256_BLOCK_0_H5_o(3) => SHA256_BLOCK_0_H5_o(3), 
        SHA256_BLOCK_0_H5_o(2) => SHA256_BLOCK_0_H5_o(2), 
        SHA256_BLOCK_0_H5_o(1) => SHA256_BLOCK_0_H5_o(1), 
        SHA256_BLOCK_0_H5_o(0) => SHA256_BLOCK_0_H5_o(0), 
        SHA256_BLOCK_0_H6_o(31) => SHA256_BLOCK_0_H6_o(31), 
        SHA256_BLOCK_0_H6_o(30) => SHA256_BLOCK_0_H6_o(30), 
        SHA256_BLOCK_0_H6_o(29) => SHA256_BLOCK_0_H6_o(29), 
        SHA256_BLOCK_0_H6_o(28) => SHA256_BLOCK_0_H6_o(28), 
        SHA256_BLOCK_0_H6_o(27) => SHA256_BLOCK_0_H6_o(27), 
        SHA256_BLOCK_0_H6_o(26) => SHA256_BLOCK_0_H6_o(26), 
        SHA256_BLOCK_0_H6_o(25) => SHA256_BLOCK_0_H6_o(25), 
        SHA256_BLOCK_0_H6_o(24) => SHA256_BLOCK_0_H6_o(24), 
        SHA256_BLOCK_0_H6_o(23) => SHA256_BLOCK_0_H6_o(23), 
        SHA256_BLOCK_0_H6_o(22) => SHA256_BLOCK_0_H6_o(22), 
        SHA256_BLOCK_0_H6_o(21) => SHA256_BLOCK_0_H6_o(21), 
        SHA256_BLOCK_0_H6_o(20) => SHA256_BLOCK_0_H6_o(20), 
        SHA256_BLOCK_0_H6_o(19) => SHA256_BLOCK_0_H6_o(19), 
        SHA256_BLOCK_0_H6_o(18) => SHA256_BLOCK_0_H6_o(18), 
        SHA256_BLOCK_0_H6_o(17) => SHA256_BLOCK_0_H6_o(17), 
        SHA256_BLOCK_0_H6_o(16) => SHA256_BLOCK_0_H6_o(16), 
        SHA256_BLOCK_0_H6_o(15) => SHA256_BLOCK_0_H6_o(15), 
        SHA256_BLOCK_0_H6_o(14) => SHA256_BLOCK_0_H6_o(14), 
        SHA256_BLOCK_0_H6_o(13) => SHA256_BLOCK_0_H6_o(13), 
        SHA256_BLOCK_0_H6_o(12) => SHA256_BLOCK_0_H6_o(12), 
        SHA256_BLOCK_0_H6_o(11) => SHA256_BLOCK_0_H6_o(11), 
        SHA256_BLOCK_0_H6_o(10) => SHA256_BLOCK_0_H6_o(10), 
        SHA256_BLOCK_0_H6_o(9) => SHA256_BLOCK_0_H6_o(9), 
        SHA256_BLOCK_0_H6_o(8) => SHA256_BLOCK_0_H6_o(8), 
        SHA256_BLOCK_0_H6_o(7) => SHA256_BLOCK_0_H6_o(7), 
        SHA256_BLOCK_0_H6_o(6) => SHA256_BLOCK_0_H6_o(6), 
        SHA256_BLOCK_0_H6_o(5) => SHA256_BLOCK_0_H6_o(5), 
        SHA256_BLOCK_0_H6_o(4) => SHA256_BLOCK_0_H6_o(4), 
        SHA256_BLOCK_0_H6_o(3) => SHA256_BLOCK_0_H6_o(3), 
        SHA256_BLOCK_0_H6_o(2) => SHA256_BLOCK_0_H6_o(2), 
        SHA256_BLOCK_0_H6_o(1) => SHA256_BLOCK_0_H6_o(1), 
        SHA256_BLOCK_0_H6_o(0) => SHA256_BLOCK_0_H6_o(0), 
        SHA256_BLOCK_0_H7_o(31) => SHA256_BLOCK_0_H7_o(31), 
        SHA256_BLOCK_0_H7_o(30) => SHA256_BLOCK_0_H7_o(30), 
        SHA256_BLOCK_0_H7_o(29) => SHA256_BLOCK_0_H7_o(29), 
        SHA256_BLOCK_0_H7_o(28) => SHA256_BLOCK_0_H7_o(28), 
        SHA256_BLOCK_0_H7_o(27) => SHA256_BLOCK_0_H7_o(27), 
        SHA256_BLOCK_0_H7_o(26) => SHA256_BLOCK_0_H7_o(26), 
        SHA256_BLOCK_0_H7_o(25) => SHA256_BLOCK_0_H7_o(25), 
        SHA256_BLOCK_0_H7_o(24) => SHA256_BLOCK_0_H7_o(24), 
        SHA256_BLOCK_0_H7_o(23) => SHA256_BLOCK_0_H7_o(23), 
        SHA256_BLOCK_0_H7_o(22) => SHA256_BLOCK_0_H7_o(22), 
        SHA256_BLOCK_0_H7_o(21) => SHA256_BLOCK_0_H7_o(21), 
        SHA256_BLOCK_0_H7_o(20) => SHA256_BLOCK_0_H7_o(20), 
        SHA256_BLOCK_0_H7_o(19) => SHA256_BLOCK_0_H7_o(19), 
        SHA256_BLOCK_0_H7_o(18) => SHA256_BLOCK_0_H7_o(18), 
        SHA256_BLOCK_0_H7_o(17) => SHA256_BLOCK_0_H7_o(17), 
        SHA256_BLOCK_0_H7_o(16) => SHA256_BLOCK_0_H7_o(16), 
        SHA256_BLOCK_0_H7_o(15) => SHA256_BLOCK_0_H7_o(15), 
        SHA256_BLOCK_0_H7_o(14) => SHA256_BLOCK_0_H7_o(14), 
        SHA256_BLOCK_0_H7_o(13) => SHA256_BLOCK_0_H7_o(13), 
        SHA256_BLOCK_0_H7_o(12) => SHA256_BLOCK_0_H7_o(12), 
        SHA256_BLOCK_0_H7_o(11) => SHA256_BLOCK_0_H7_o(11), 
        SHA256_BLOCK_0_H7_o(10) => SHA256_BLOCK_0_H7_o(10), 
        SHA256_BLOCK_0_H7_o(9) => SHA256_BLOCK_0_H7_o(9), 
        SHA256_BLOCK_0_H7_o(8) => SHA256_BLOCK_0_H7_o(8), 
        SHA256_BLOCK_0_H7_o(7) => SHA256_BLOCK_0_H7_o(7), 
        SHA256_BLOCK_0_H7_o(6) => SHA256_BLOCK_0_H7_o(6), 
        SHA256_BLOCK_0_H7_o(5) => SHA256_BLOCK_0_H7_o(5), 
        SHA256_BLOCK_0_H7_o(4) => SHA256_BLOCK_0_H7_o(4), 
        SHA256_BLOCK_0_H7_o(3) => SHA256_BLOCK_0_H7_o(3), 
        SHA256_BLOCK_0_H7_o(2) => SHA256_BLOCK_0_H7_o(2), 
        SHA256_BLOCK_0_H7_o(1) => SHA256_BLOCK_0_H7_o(1), 
        SHA256_BLOCK_0_H7_o(0) => SHA256_BLOCK_0_H7_o(0), state_2
         => \state[3]\, state_0 => \state[1]\, state_3 => 
        \state[4]\, sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, SHA256_Module_0_di_req_o
         => \SHA256_Module_0_di_req_o\, 
        SHA256_Module_0_do_valid_o => 
        \SHA256_Module_0_do_valid_o\, sha256_controller_0_end_o
         => sha256_controller_0_end_o, last_block_0 => 
        last_block_0, ce_i_i_2 => ce_i_i_2, N_28 => N_28, 
        SHA256_Module_0_error_o => SHA256_Module_0_error_o, 
        N_1696 => N_1696, N_1400 => N_1400, N_1624 => N_1624, 
        N_920 => N_920, N_1144 => N_1144, N_1399 => N_1399, 
        N_1623 => N_1623, N_919 => N_919, N_1143 => N_1143, 
        N_1401 => N_1401, N_1625 => N_1625, N_921 => N_921, 
        N_1145 => N_1145, ren_pos => ren_pos, N_1694 => N_1694, 
        N_1692 => N_1692, N_1693 => N_1693, N_1691 => N_1691, 
        N_1690 => N_1690, N_89 => N_89, N_1695 => N_1695, N_1708
         => N_1708, N_1709 => N_1709, N_1707 => N_1707, N_1706
         => N_1706, N_1705 => N_1705, N_1704 => N_1704, N_1703
         => N_1703, N_1700 => N_1700, N_1701 => N_1701, N_1697
         => N_1697, N_1699 => N_1699, N_1698 => N_1698, N_1717
         => N_1717, N_1712 => N_1712, N_1716 => N_1716, N_1715
         => N_1715, N_1711 => N_1711, N_1713 => N_1713, N_1714
         => N_1714, N_1718 => N_1718, N_1702 => N_1702, N_1710
         => N_1710);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    limiter_1cycle_first : limiter_1cycle_0
      port map(prev_sig => prev_sig, sha256_system_sb_0_FIC_0_CLK
         => sha256_system_sb_0_FIC_0_CLK, first_block => 
        first_block);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    limiter_1cycle_ready : limiter_1cycle_1
      port map(prev_sig => prev_sig_0, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, 
        SHA256_Module_0_data_out_ready => 
        \SHA256_Module_0_data_out_ready\);
    
    reg_17x32_0 : reg_17x32
      port map(AHB_slave_dummy_0_mem_wdata(31) => 
        AHB_slave_dummy_0_mem_wdata(31), 
        AHB_slave_dummy_0_mem_wdata(30) => 
        AHB_slave_dummy_0_mem_wdata(30), 
        AHB_slave_dummy_0_mem_wdata(29) => 
        AHB_slave_dummy_0_mem_wdata(29), 
        AHB_slave_dummy_0_mem_wdata(28) => 
        AHB_slave_dummy_0_mem_wdata(28), 
        AHB_slave_dummy_0_mem_wdata(27) => 
        AHB_slave_dummy_0_mem_wdata(27), 
        AHB_slave_dummy_0_mem_wdata(26) => 
        AHB_slave_dummy_0_mem_wdata(26), 
        AHB_slave_dummy_0_mem_wdata(25) => 
        AHB_slave_dummy_0_mem_wdata(25), 
        AHB_slave_dummy_0_mem_wdata(24) => 
        AHB_slave_dummy_0_mem_wdata(24), 
        AHB_slave_dummy_0_mem_wdata(23) => 
        AHB_slave_dummy_0_mem_wdata(23), 
        AHB_slave_dummy_0_mem_wdata(22) => 
        AHB_slave_dummy_0_mem_wdata(22), 
        AHB_slave_dummy_0_mem_wdata(21) => 
        AHB_slave_dummy_0_mem_wdata(21), 
        AHB_slave_dummy_0_mem_wdata(20) => 
        AHB_slave_dummy_0_mem_wdata(20), 
        AHB_slave_dummy_0_mem_wdata(19) => 
        AHB_slave_dummy_0_mem_wdata(19), 
        AHB_slave_dummy_0_mem_wdata(18) => 
        AHB_slave_dummy_0_mem_wdata(18), 
        AHB_slave_dummy_0_mem_wdata(17) => 
        AHB_slave_dummy_0_mem_wdata(17), 
        AHB_slave_dummy_0_mem_wdata(16) => 
        AHB_slave_dummy_0_mem_wdata(16), 
        AHB_slave_dummy_0_mem_wdata(15) => 
        AHB_slave_dummy_0_mem_wdata(15), 
        AHB_slave_dummy_0_mem_wdata(14) => 
        AHB_slave_dummy_0_mem_wdata(14), 
        AHB_slave_dummy_0_mem_wdata(13) => 
        AHB_slave_dummy_0_mem_wdata(13), 
        AHB_slave_dummy_0_mem_wdata(12) => 
        AHB_slave_dummy_0_mem_wdata(12), 
        AHB_slave_dummy_0_mem_wdata(11) => 
        AHB_slave_dummy_0_mem_wdata(11), 
        AHB_slave_dummy_0_mem_wdata(10) => 
        AHB_slave_dummy_0_mem_wdata(10), 
        AHB_slave_dummy_0_mem_wdata(9) => 
        AHB_slave_dummy_0_mem_wdata(9), 
        AHB_slave_dummy_0_mem_wdata(8) => 
        AHB_slave_dummy_0_mem_wdata(8), 
        AHB_slave_dummy_0_mem_wdata(7) => 
        AHB_slave_dummy_0_mem_wdata(7), 
        AHB_slave_dummy_0_mem_wdata(6) => 
        AHB_slave_dummy_0_mem_wdata(6), 
        AHB_slave_dummy_0_mem_wdata(5) => 
        AHB_slave_dummy_0_mem_wdata(5), 
        AHB_slave_dummy_0_mem_wdata(4) => 
        AHB_slave_dummy_0_mem_wdata(4), 
        AHB_slave_dummy_0_mem_wdata(3) => 
        AHB_slave_dummy_0_mem_wdata(3), 
        AHB_slave_dummy_0_mem_wdata(2) => 
        AHB_slave_dummy_0_mem_wdata(2), 
        AHB_slave_dummy_0_mem_wdata(1) => 
        AHB_slave_dummy_0_mem_wdata(1), 
        AHB_slave_dummy_0_mem_wdata(0) => 
        AHB_slave_dummy_0_mem_wdata(0), 
        sha256_controller_0_read_addr_0(3) => 
        \sha256_controller_0_read_addr_0[3]\, 
        sha256_controller_0_read_addr_0(2) => 
        \sha256_controller_0_read_addr_0[2]\, 
        sha256_controller_0_read_addr_0(1) => 
        \sha256_controller_0_read_addr_0[1]\, 
        sha256_controller_0_read_addr_0(0) => 
        \sha256_controller_0_read_addr_0[0]\, waddr_in_net_0(4)
         => waddr_in_net_0(4), waddr_in_net_0(3) => 
        waddr_in_net_0(3), waddr_in_net_0(2) => waddr_in_net_0(2), 
        waddr_in_net_0(1) => waddr_in_net_0(1), waddr_in_net_0(0)
         => waddr_in_net_0(0), raddr_pos_3 => \raddr_pos[3]\, 
        raddr_pos_2 => \raddr_pos[2]\, 
        SHA256_Module_0_data_out_ready => 
        \SHA256_Module_0_data_out_ready\, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, 
        sha256_system_sb_0_GPIO_9_M2F => 
        sha256_system_sb_0_GPIO_9_M2F, 
        SHA256_Module_0_data_available => 
        SHA256_Module_0_data_available, ren_pos => ren_pos, 
        last_block => last_block, first_block => first_block, 
        N_1717 => N_1717, N_1716 => N_1716, N_1711 => N_1711, 
        N_1710 => N_1710, N_1708 => N_1708, N_1705 => N_1705, 
        N_1704 => N_1704, N_1701 => N_1701, N_1690 => N_1690, 
        N_1691 => N_1691, N_1707 => N_1707, N_1703 => N_1703, 
        N_1715 => N_1715, N_1700 => N_1700, N_1714 => N_1714, 
        N_1697 => N_1697, N_1693 => N_1693, N_1706 => N_1706, 
        N_1696 => N_1696, N_1709 => N_1709, N_1698 => N_1698, 
        N_1699 => N_1699, N_1694 => N_1694, N_1702 => N_1702, 
        N_1712 => N_1712, N_1695 => N_1695, N_1692 => N_1692, 
        N_1718 => N_1718, N_1713 => N_1713, N_1144 => N_1144, 
        N_921 => N_921, N_1401 => N_1401, N_1145 => N_1145, N_919
         => N_919, N_1400 => N_1400, N_1623 => N_1623, N_920 => 
        N_920, N_1143 => N_1143, N_1624 => N_1624, N_1625 => 
        N_1625, N_1399 => N_1399, sha256_system_sb_0_GPIO_1_M2F
         => sha256_system_sb_0_GPIO_1_M2F, 
        AHB_slave_dummy_0_write_en => AHB_slave_dummy_0_write_en);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_1 is

    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o            : in    std_logic_vector(31 downto 0);
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic;
          wen_or                         : in    std_logic;
          SHA256_Module_0_data_out_ready : in    std_logic
        );

end reg_1x32_1;

architecture DEF_ARCH of reg_1x32_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity mux_9_1 is

    port( result_addr_net_0 : in    std_logic_vector(3 downto 0);
          line_19           : in    std_logic;
          line_22           : in    std_logic;
          line_12           : in    std_logic;
          line_8            : in    std_logic;
          line_17           : in    std_logic;
          line_21           : in    std_logic;
          line_5_d0         : in    std_logic;
          line_9            : in    std_logic;
          line_13           : in    std_logic;
          line_4_d0         : in    std_logic;
          line_6_d0         : in    std_logic;
          line_18           : in    std_logic;
          line_24           : in    std_logic;
          line_29           : in    std_logic;
          line_30           : in    std_logic;
          line_27           : in    std_logic;
          line_25           : in    std_logic;
          line_16           : in    std_logic;
          line_15           : in    std_logic;
          line_1_d0         : in    std_logic;
          line_23           : in    std_logic;
          line_3_d0         : in    std_logic;
          line_14           : in    std_logic;
          line_26           : in    std_logic;
          line_2_d0         : in    std_logic;
          line_0_d0         : in    std_logic;
          line_0_19         : in    std_logic;
          line_0_22         : in    std_logic;
          line_0_12         : in    std_logic;
          line_0_8          : in    std_logic;
          line_0_17         : in    std_logic;
          line_0_21         : in    std_logic;
          line_0_5          : in    std_logic;
          line_0_9          : in    std_logic;
          line_0_13         : in    std_logic;
          line_0_4          : in    std_logic;
          line_0_6          : in    std_logic;
          line_0_18         : in    std_logic;
          line_0_24         : in    std_logic;
          line_0_29         : in    std_logic;
          line_0_30         : in    std_logic;
          line_0_27         : in    std_logic;
          line_0_25         : in    std_logic;
          line_0_16         : in    std_logic;
          line_0_15         : in    std_logic;
          line_0_1          : in    std_logic;
          line_0_23         : in    std_logic;
          line_0_3          : in    std_logic;
          line_0_14         : in    std_logic;
          line_0_26         : in    std_logic;
          line_0_2          : in    std_logic;
          line_0_0          : in    std_logic;
          line_1_19         : in    std_logic;
          line_1_22         : in    std_logic;
          line_1_12         : in    std_logic;
          line_1_8          : in    std_logic;
          line_1_17         : in    std_logic;
          line_1_21         : in    std_logic;
          line_1_5          : in    std_logic;
          line_1_9          : in    std_logic;
          line_1_13         : in    std_logic;
          line_1_4          : in    std_logic;
          line_1_6          : in    std_logic;
          line_1_18         : in    std_logic;
          line_1_24         : in    std_logic;
          line_1_29         : in    std_logic;
          line_1_30         : in    std_logic;
          line_1_27         : in    std_logic;
          line_1_25         : in    std_logic;
          line_1_16         : in    std_logic;
          line_1_15         : in    std_logic;
          line_1_1          : in    std_logic;
          line_1_23         : in    std_logic;
          line_1_3          : in    std_logic;
          line_1_14         : in    std_logic;
          line_1_26         : in    std_logic;
          line_1_2          : in    std_logic;
          line_1_0          : in    std_logic;
          line_2_19         : in    std_logic;
          line_2_22         : in    std_logic;
          line_2_12         : in    std_logic;
          line_2_8          : in    std_logic;
          line_2_17         : in    std_logic;
          line_2_21         : in    std_logic;
          line_2_5          : in    std_logic;
          line_2_9          : in    std_logic;
          line_2_13         : in    std_logic;
          line_2_4          : in    std_logic;
          line_2_6          : in    std_logic;
          line_2_18         : in    std_logic;
          line_2_24         : in    std_logic;
          line_2_29         : in    std_logic;
          line_2_30         : in    std_logic;
          line_2_27         : in    std_logic;
          line_2_25         : in    std_logic;
          line_2_16         : in    std_logic;
          line_2_15         : in    std_logic;
          line_2_1          : in    std_logic;
          line_2_23         : in    std_logic;
          line_2_3          : in    std_logic;
          line_2_14         : in    std_logic;
          line_2_26         : in    std_logic;
          line_2_2          : in    std_logic;
          line_2_0          : in    std_logic;
          line_3_22         : in    std_logic;
          line_3_12         : in    std_logic;
          line_3_4          : in    std_logic;
          line_3_6          : in    std_logic;
          line_3_29         : in    std_logic;
          line_3_24         : in    std_logic;
          line_3_30         : in    std_logic;
          line_3_27         : in    std_logic;
          line_3_25         : in    std_logic;
          line_3_16         : in    std_logic;
          line_3_15         : in    std_logic;
          line_3_1          : in    std_logic;
          line_3_18         : in    std_logic;
          line_3_13         : in    std_logic;
          line_3_9          : in    std_logic;
          line_3_5          : in    std_logic;
          line_3_23         : in    std_logic;
          line_3_21         : in    std_logic;
          line_3_17         : in    std_logic;
          line_3_3          : in    std_logic;
          line_3_14         : in    std_logic;
          line_3_26         : in    std_logic;
          line_3_2          : in    std_logic;
          line_3_0          : in    std_logic;
          line_3_8          : in    std_logic;
          line_3_19         : in    std_logic;
          line_4_22         : in    std_logic;
          line_4_12         : in    std_logic;
          line_4_4          : in    std_logic;
          line_4_6          : in    std_logic;
          line_4_29         : in    std_logic;
          line_4_24         : in    std_logic;
          line_4_30         : in    std_logic;
          line_4_27         : in    std_logic;
          line_4_25         : in    std_logic;
          line_4_16         : in    std_logic;
          line_4_15         : in    std_logic;
          line_4_1          : in    std_logic;
          line_4_18         : in    std_logic;
          line_4_13         : in    std_logic;
          line_4_9          : in    std_logic;
          line_4_5          : in    std_logic;
          line_4_23         : in    std_logic;
          line_4_21         : in    std_logic;
          line_4_17         : in    std_logic;
          line_4_3          : in    std_logic;
          line_4_14         : in    std_logic;
          line_4_26         : in    std_logic;
          line_4_2          : in    std_logic;
          line_4_0          : in    std_logic;
          line_4_8          : in    std_logic;
          line_4_19         : in    std_logic;
          line_5_22         : in    std_logic;
          line_5_12         : in    std_logic;
          line_5_4          : in    std_logic;
          line_5_6          : in    std_logic;
          line_5_29         : in    std_logic;
          line_5_24         : in    std_logic;
          line_5_30         : in    std_logic;
          line_5_27         : in    std_logic;
          line_5_25         : in    std_logic;
          line_5_16         : in    std_logic;
          line_5_15         : in    std_logic;
          line_5_1          : in    std_logic;
          line_5_18         : in    std_logic;
          line_5_13         : in    std_logic;
          line_5_9          : in    std_logic;
          line_5_5          : in    std_logic;
          line_5_23         : in    std_logic;
          line_5_21         : in    std_logic;
          line_5_17         : in    std_logic;
          line_5_3          : in    std_logic;
          line_5_14         : in    std_logic;
          line_5_26         : in    std_logic;
          line_5_2          : in    std_logic;
          line_5_0          : in    std_logic;
          line_5_8          : in    std_logic;
          line_5_19         : in    std_logic;
          line_6_22         : in    std_logic;
          line_6_12         : in    std_logic;
          line_6_4          : in    std_logic;
          line_6_6          : in    std_logic;
          line_6_29         : in    std_logic;
          line_6_24         : in    std_logic;
          line_6_30         : in    std_logic;
          line_6_27         : in    std_logic;
          line_6_25         : in    std_logic;
          line_6_16         : in    std_logic;
          line_6_15         : in    std_logic;
          line_6_1          : in    std_logic;
          line_6_18         : in    std_logic;
          line_6_13         : in    std_logic;
          line_6_9          : in    std_logic;
          line_6_5          : in    std_logic;
          line_6_23         : in    std_logic;
          line_6_21         : in    std_logic;
          line_6_17         : in    std_logic;
          line_6_3          : in    std_logic;
          line_6_14         : in    std_logic;
          line_6_26         : in    std_logic;
          line_6_2          : in    std_logic;
          line_6_0          : in    std_logic;
          line_6_8          : in    std_logic;
          line_6_19         : in    std_logic;
          line_7_19         : in    std_logic;
          line_7_8          : in    std_logic;
          line_7_1          : in    std_logic;
          line_7_2          : in    std_logic;
          line_7_0          : in    std_logic;
          N_568             : out   std_logic;
          N_579             : out   std_logic;
          N_580             : out   std_logic;
          N_581             : out   std_logic;
          N_583             : out   std_logic;
          N_588             : out   std_logic;
          N_589             : out   std_logic;
          N_590             : out   std_logic;
          N_591             : out   std_logic;
          N_592             : out   std_logic;
          N_595             : out   std_logic;
          N_594             : out   std_logic;
          N_586             : out   std_logic;
          N_582             : out   std_logic;
          N_578             : out   std_logic;
          N_574             : out   std_logic;
          N_571             : out   std_logic;
          N_570             : out   std_logic;
          N_569             : out   std_logic;
          N_96              : out   std_logic;
          N_81              : out   std_logic;
          N_74              : out   std_logic;
          N_75              : out   std_logic;
          N_499             : out   std_logic;
          N_501             : out   std_logic;
          N_525             : out   std_logic;
          N_513             : out   std_logic;
          N_502             : out   std_logic;
          N_522             : out   std_logic;
          N_500             : out   std_logic;
          N_514             : out   std_logic;
          N_515             : out   std_logic;
          N_524             : out   std_logic;
          N_526             : out   std_logic;
          N_529             : out   std_logic;
          N_528             : out   std_logic;
          N_523             : out   std_logic;
          N_517             : out   std_logic;
          N_505             : out   std_logic;
          N_503             : out   std_logic;
          N_512             : out   std_logic;
          N_508             : out   std_logic;
          N_504             : out   std_logic;
          N_520             : out   std_logic;
          N_516             : out   std_logic;
          ren_pos           : in    std_logic;
          N_228             : out   std_logic;
          N_7               : out   std_logic;
          N_566             : out   std_logic;
          N_567             : out   std_logic;
          N_565             : out   std_logic
        );

end mux_9_1;

architecture DEF_ARCH of mux_9_1 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \data_out_5_bm[3]_net_1\, \data_out_5_am[3]_net_1\, 
        \data_out_5_bm[14]_net_1\, \data_out_5_am[14]_net_1\, 
        \data_out_5_bm[15]_net_1\, \data_out_5_am[15]_net_1\, 
        \data_out_5_bm[16]_net_1\, \data_out_5_am[16]_net_1\, 
        \data_out_5_bm[18]_net_1\, \data_out_5_am[18]_net_1\, 
        \data_out_5_bm[23]_net_1\, \data_out_5_am[23]_net_1\, 
        \data_out_5_bm[24]_net_1\, \data_out_5_am[24]_net_1\, 
        \data_out_5_bm[25]_net_1\, \data_out_5_am[25]_net_1\, 
        \data_out_5_bm[26]_net_1\, \data_out_5_am[26]_net_1\, 
        \data_out_5_bm[27]_net_1\, \data_out_5_am[27]_net_1\, 
        \data_out_5_bm[30]_net_1\, \data_out_5_am[30]_net_1\, 
        \data_out_5_bm[29]_net_1\, \data_out_5_am[29]_net_1\, 
        \data_out_5_bm[21]_net_1\, \data_out_5_am[21]_net_1\, 
        \data_out_5_bm[17]_net_1\, \data_out_5_am[17]_net_1\, 
        \data_out_5_bm[13]_net_1\, \data_out_5_am[13]_net_1\, 
        \data_out_5_bm[9]_net_1\, \data_out_5_am[9]_net_1\, 
        \data_out_5_bm[6]_net_1\, \data_out_5_am[6]_net_1\, 
        \data_out_5_bm[5]_net_1\, \data_out_5_am[5]_net_1\, 
        \data_out_5_bm[4]_net_1\, \data_out_5_am[4]_net_1\, 
        \data_out_6_i_m2_1_1[19]\, N_255, 
        \data_out_i_m2_4_1_1[22]\, N_83, 
        \data_out_i_m2_4_1_1[12]\, N_68, \data_out_6_i_m2_1_1[8]\, 
        N_211, \data_out_i_m2_ns_1_1_1[22]_net_1\, 
        \data_out_i_m2_ns_1[22]_net_1\, 
        \data_out_i_m2_ns_1_1_1[12]_net_1\, 
        \data_out_i_m2_ns_1[12]_net_1\, 
        \data_out_4_i_m2_bm[19]_net_1\, 
        \data_out_4_i_m2_am[19]_net_1\, 
        \data_out_4_i_m2_bm[8]_net_1\, 
        \data_out_4_i_m2_am[8]_net_1\, \data_out_5_bm[0]_net_1\, 
        \data_out_5_am[0]_net_1\, N_531, \data_out_4_bm[0]_net_1\, 
        \data_out_4_am[0]_net_1\, \data_out_5_bm[2]_net_1\, 
        \data_out_5_am[2]_net_1\, N_533, \data_out_4_bm[2]_net_1\, 
        \data_out_4_am[2]_net_1\, \data_out_4_bm[26]_net_1\, 
        \data_out_4_am[26]_net_1\, \data_out_4_bm[14]_net_1\, 
        \data_out_4_am[14]_net_1\, \data_out_4_bm[3]_net_1\, 
        \data_out_4_am[3]_net_1\, \data_out_4_bm[23]_net_1\, 
        \data_out_4_am[23]_net_1\, \data_out_4_bm[1]_net_1\, 
        \data_out_4_am[1]_net_1\, \data_out_4_bm[15]_net_1\, 
        \data_out_4_am[15]_net_1\, \data_out_4_bm[16]_net_1\, 
        \data_out_4_am[16]_net_1\, \data_out_4_bm[25]_net_1\, 
        \data_out_4_am[25]_net_1\, \data_out_4_bm[27]_net_1\, 
        \data_out_4_am[27]_net_1\, \data_out_4_bm[30]_net_1\, 
        \data_out_4_am[30]_net_1\, \data_out_5_bm[1]_net_1\, 
        \data_out_5_am[1]_net_1\, N_532, 
        \data_out_4_bm[29]_net_1\, \data_out_4_am[29]_net_1\, 
        \data_out_4_bm[24]_net_1\, \data_out_4_am[24]_net_1\, 
        \data_out_4_bm[18]_net_1\, \data_out_4_am[18]_net_1\, 
        \data_out_4_bm[6]_net_1\, \data_out_4_am[6]_net_1\, 
        \data_out_4_bm[4]_net_1\, \data_out_4_am[4]_net_1\, 
        \data_out_4_bm[13]_net_1\, \data_out_4_am[13]_net_1\, 
        \data_out_4_bm[9]_net_1\, \data_out_4_am[9]_net_1\, 
        \data_out_4_bm[5]_net_1\, \data_out_4_am[5]_net_1\, 
        \data_out_4_bm[21]_net_1\, \data_out_4_am[21]_net_1\, 
        \data_out_4_bm[17]_net_1\, \data_out_4_am[17]_net_1\, 
        GND_net_1, VCC_net_1 : std_logic;

begin 


    \data_out_5_bm[2]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_2, B => line_4_2, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[2]_net_1\);
    
    \data_out_4_am[24]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_24, B => line_2_24, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[24]_net_1\);
    
    \data_out_6_i_RNO[19]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => result_addr_net_0(1), B => 
        \data_out_6_i_m2_1_1[19]\, C => line_19, D => line_0_19, 
        Y => N_255);
    
    \data_out_6[29]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[29]_net_1\, D
         => \data_out_5_am[29]_net_1\, Y => N_594);
    
    \data_out_6[9]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[9]_net_1\, D
         => \data_out_5_am[9]_net_1\, Y => N_574);
    
    \data_out_5_am[0]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_0, B => line_6_0, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[0]_net_1\);
    
    \data_out_4_bm[15]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_15, B => line_4_15, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[15]_net_1\);
    
    \data_out_6[3]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[3]_net_1\, D
         => \data_out_5_am[3]_net_1\, Y => N_568);
    
    \data_out_5_ns[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_5_bm[0]_net_1\, C => \data_out_5_am[0]_net_1\, 
        Y => N_531);
    
    \data_out_i_m2_ns_RNO_0[12]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_12, B => line_2_12, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \data_out_i_m2_4_1_1[12]\);
    
    \data_out_6[4]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[4]_net_1\, D
         => \data_out_5_am[4]_net_1\, Y => N_569);
    
    \data_out_4_ns[16]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[16]_net_1\, C => \data_out_4_am[16]_net_1\, 
        Y => N_515);
    
    \data_out_5_am[2]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_2, B => line_6_2, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[2]_net_1\);
    
    \data_out_4_ns[5]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[5]_net_1\, C => \data_out_4_am[5]_net_1\, 
        Y => N_504);
    
    \data_out_6[6]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[6]_net_1\, D
         => \data_out_5_am[6]_net_1\, Y => N_571);
    
    \data_out_4_bm[5]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_d0, B => line_0_5, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[5]_net_1\);
    
    \data_out_4_bm[25]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_25, B => line_4_25, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[25]_net_1\);
    
    \data_out_4_bm[9]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_9, B => line_0_9, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[9]_net_1\);
    
    \data_out_4_am[30]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_30, B => line_6_30, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[30]_net_1\);
    
    \data_out_5_am[13]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_13, B => line_6_13, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[13]_net_1\);
    
    \data_out_4_ns[26]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[26]_net_1\, C => \data_out_4_am[26]_net_1\, 
        Y => N_525);
    
    \data_out_5_bm[16]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_16, B => line_0_16, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[16]_net_1\);
    
    \data_out_4_bm[14]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_14, B => line_0_14, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[14]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \data_out_4_bm[0]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_0_d0, B => line_0_0, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[0]_net_1\);
    
    \data_out_5_am[23]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_23, B => line_2_23, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[23]_net_1\);
    
    \data_out_5_bm[18]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_18, B => line_4_18, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[18]_net_1\);
    
    \data_out_4_ns[6]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[6]_net_1\, C => \data_out_4_am[6]_net_1\, 
        Y => N_505);
    
    \data_out_5_bm[26]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_26, B => line_4_26, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[26]_net_1\);
    
    \data_out_6_i_RNO_0[19]\ : CFG4
      generic map(INIT => x"350F")

      port map(A => line_1_19, B => line_2_19, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \data_out_6_i_m2_1_1[19]\);
    
    \data_out_5_ns[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_5_bm[1]_net_1\, C => \data_out_5_am[1]_net_1\, 
        Y => N_532);
    
    \data_out_4_bm[24]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_24, B => line_0_24, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[24]_net_1\);
    
    \data_out_4_ns[3]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[3]_net_1\, C => \data_out_4_am[3]_net_1\, 
        Y => N_502);
    
    \data_out_5_am[15]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_15, B => line_2_15, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[15]_net_1\);
    
    \data_out_4_bm[2]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_2_d0, B => line_0_2, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[2]_net_1\);
    
    \data_out_6_i_RNO[8]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => result_addr_net_0(1), B => 
        \data_out_6_i_m2_1_1[8]\, C => line_8, D => line_0_8, Y
         => N_211);
    
    \data_out_4_i_m2_bm[19]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_19, B => line_4_19, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_i_m2_bm[19]_net_1\);
    
    \data_out_4_am[1]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_1, B => line_6_1, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[1]_net_1\);
    
    \data_out_4_i_m2_am[8]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_8, B => line_6_8, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_i_m2_am[8]_net_1\);
    
    \data_out_5_bm[13]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_13, B => line_4_13, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[13]_net_1\);
    
    \data_out_4_am[17]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_17, B => line_2_17, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[17]_net_1\);
    
    \data_out_5_am[25]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_25, B => line_2_25, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[25]_net_1\);
    
    \data_out_6[18]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[18]_net_1\, D
         => \data_out_5_am[18]_net_1\, Y => N_583);
    
    \data_out_4_i_m2_ns[8]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_i_m2_bm[8]_net_1\, C => 
        \data_out_4_i_m2_am[8]_net_1\, Y => N_75);
    
    \data_out_i_m2_ns_1_1_1[12]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_12, B => line_6_12, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \data_out_i_m2_ns_1_1_1[12]_net_1\);
    
    \data_out_4_ns[13]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[13]_net_1\, C => \data_out_4_am[13]_net_1\, 
        Y => N_512);
    
    \data_out_4_ns[18]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[18]_net_1\, C => \data_out_4_am[18]_net_1\, 
        Y => N_517);
    
    \data_out_5_bm[1]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_d0, B => line_0_1, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[1]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \data_out_6[21]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[21]_net_1\, D
         => \data_out_5_am[21]_net_1\, Y => N_586);
    
    \data_out_4_ns[9]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[9]_net_1\, C => \data_out_4_am[9]_net_1\, 
        Y => N_508);
    
    \data_out_4_am[15]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_15, B => line_6_15, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[15]_net_1\);
    
    \data_out_4_bm[30]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_30, B => line_4_30, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[30]_net_1\);
    
    \data_out_5_bm[21]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_21, B => line_4_21, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[21]_net_1\);
    
    \data_out_6[30]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[30]_net_1\, D
         => \data_out_5_am[30]_net_1\, Y => N_595);
    
    \data_out_6[23]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[23]_net_1\, D
         => \data_out_5_am[23]_net_1\, Y => N_588);
    
    \data_out_5_bm[23]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_23, B => line_0_23, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[23]_net_1\);
    
    \data_out_4_ns[4]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[4]_net_1\, C => \data_out_4_am[4]_net_1\, 
        Y => N_503);
    
    \data_out_4_bm[16]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_16, B => line_4_16, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[16]_net_1\);
    
    \data_out_4_am[27]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_27, B => line_6_27, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[27]_net_1\);
    
    \data_out_5_am[17]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_17, B => line_6_17, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[17]_net_1\);
    
    \data_out_4_ns[23]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[23]_net_1\, C => \data_out_4_am[23]_net_1\, 
        Y => N_522);
    
    \data_out_4_bm[18]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_18, B => line_0_18, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[18]_net_1\);
    
    \data_out_i_m2_ns_RNO[12]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => result_addr_net_0(1), B => 
        \data_out_i_m2_4_1_1[12]\, C => line_12, D => line_0_12, 
        Y => N_68);
    
    \data_out_4_bm[29]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_29, B => line_0_29, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[29]_net_1\);
    
    \data_out_4_am[3]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_3, B => line_2_3, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[3]_net_1\);
    
    \data_out_i_m2_ns_RNO_0[22]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_22, B => line_2_22, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \data_out_i_m2_4_1_1[22]\);
    
    \data_out_4_am[25]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_25, B => line_6_25, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[25]_net_1\);
    
    \data_out_5_bm[15]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_15, B => line_0_15, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[15]_net_1\);
    
    \data_out_4_ns[29]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[29]_net_1\, C => \data_out_4_am[29]_net_1\, 
        Y => N_528);
    
    \data_out_4_ns[2]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[2]_net_1\, C => \data_out_4_am[2]_net_1\, 
        Y => N_501);
    
    \data_out_4_ns[14]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[14]_net_1\, C => \data_out_4_am[14]_net_1\, 
        Y => N_513);
    
    \data_out_5_bm[3]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_3, B => line_4_3, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[3]_net_1\);
    
    \data_out_5_am[1]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_1, B => line_2_1, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[1]_net_1\);
    
    \data_out_4_bm[26]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_26, B => line_0_26, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[26]_net_1\);
    
    \data_out_5_am[27]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_27, B => line_2_27, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[27]_net_1\);
    
    \data_out_5_bm[25]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_25, B => line_0_25, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[25]_net_1\);
    
    \data_out_4_ns[24]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[24]_net_1\, C => \data_out_4_am[24]_net_1\, 
        Y => N_523);
    
    \data_out_4_am[4]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_4, B => line_2_4, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[4]_net_1\);
    
    \data_out_6[13]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[13]_net_1\, D
         => \data_out_5_am[13]_net_1\, Y => N_578);
    
    \data_out_4_bm[17]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_17, B => line_0_17, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[17]_net_1\);
    
    \data_out_4_am[21]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_21, B => line_2_21, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[21]_net_1\);
    
    \data_out_5_bm[4]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_4, B => line_4_4, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[4]_net_1\);
    
    \data_out_5_am[3]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_3, B => line_6_3, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[3]_net_1\);
    
    \data_out_4_am[18]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_18, B => line_2_18, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[18]_net_1\);
    
    \data_out_6[26]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[26]_net_1\, D
         => \data_out_5_am[26]_net_1\, Y => N_591);
    
    \data_out_4_bm[21]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_21, B => line_0_21, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[21]_net_1\);
    
    \data_out_5_am[21]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_21, B => line_6_21, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[21]_net_1\);
    
    \data_out_4_bm[27]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_27, B => line_4_27, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[27]_net_1\);
    
    \data_out_4_am[6]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_6, B => line_2_6, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[6]_net_1\);
    
    \data_out_6[25]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[25]_net_1\, D
         => \data_out_5_am[25]_net_1\, Y => N_590);
    
    \data_out_4_bm[1]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_1, B => line_4_1, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[1]_net_1\);
    
    \data_out_5_am[29]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_29, B => line_6_29, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[29]_net_1\);
    
    \data_out_6_i[8]\ : CFG4
      generic map(INIT => x"27FF")

      port map(A => result_addr_net_0(3), B => line_7_8, C => 
        N_211, D => ren_pos, Y => N_7);
    
    \data_out_6[5]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[5]_net_1\, D
         => \data_out_5_am[5]_net_1\, Y => N_570);
    
    \data_out_4_am[16]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_16, B => line_6_16, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[16]_net_1\);
    
    \data_out_5_bm[6]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_6, B => line_4_6, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[6]_net_1\);
    
    \data_out_5_am[14]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_14, B => line_6_14, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[14]_net_1\);
    
    \data_out_4_ns[15]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[15]_net_1\, C => \data_out_4_am[15]_net_1\, 
        Y => N_514);
    
    \data_out_5_am[4]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_4, B => line_6_4, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[4]_net_1\);
    
    \data_out_5_bm[17]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_17, B => line_4_17, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[17]_net_1\);
    
    \data_out_4_am[13]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_13, B => line_2_13, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[13]_net_1\);
    
    \data_out_6[1]\ : CFG4
      generic map(INIT => x"D850")

      port map(A => result_addr_net_0(3), B => line_7_1, C => 
        N_532, D => ren_pos, Y => N_566);
    
    \data_out_5_bm[29]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_29, B => line_4_29, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[29]_net_1\);
    
    \data_out_4_ns[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[0]_net_1\, C => \data_out_4_am[0]_net_1\, 
        Y => N_499);
    
    \data_out_6[16]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[16]_net_1\, D
         => \data_out_5_am[16]_net_1\, Y => N_581);
    
    \data_out_5_bm[14]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_14, B => line_4_14, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[14]_net_1\);
    
    \data_out_4_ns[25]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[25]_net_1\, C => \data_out_4_am[25]_net_1\, 
        Y => N_524);
    
    \data_out_4_am[26]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_26, B => line_2_26, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[26]_net_1\);
    
    \data_out_5_am[24]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_24, B => line_6_24, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[24]_net_1\);
    
    \data_out_4_bm[3]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_d0, B => line_0_3, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[3]_net_1\);
    
    \data_out_4_am[29]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_29, B => line_2_29, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[29]_net_1\);
    
    \data_out_4_i_m2_bm[8]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_8, B => line_4_8, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_i_m2_bm[8]_net_1\);
    
    \data_out_6[15]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[15]_net_1\, D
         => \data_out_5_am[15]_net_1\, Y => N_580);
    
    \data_out_6[27]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[27]_net_1\, D
         => \data_out_5_am[27]_net_1\, Y => N_592);
    
    \data_out_5_bm[27]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_27, B => line_0_27, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[27]_net_1\);
    
    \data_out_4_am[23]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_23, B => line_6_23, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[23]_net_1\);
    
    \data_out_5_am[6]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_6, B => line_6_6, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[6]_net_1\);
    
    \data_out_i_m2_ns_1[22]\ : CFG4
      generic map(INIT => x"46CE")

      port map(A => result_addr_net_0(1), B => 
        \data_out_i_m2_ns_1_1_1[22]_net_1\, C => line_3_22, D => 
        line_4_22, Y => \data_out_i_m2_ns_1[22]_net_1\);
    
    \data_out_5_bm[24]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_24, B => line_4_24, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[24]_net_1\);
    
    \data_out_6_i[19]\ : CFG4
      generic map(INIT => x"27FF")

      port map(A => result_addr_net_0(3), B => line_7_19, C => 
        N_255, D => ren_pos, Y => N_228);
    
    \data_out_6[24]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[24]_net_1\, D
         => \data_out_5_am[24]_net_1\, Y => N_589);
    
    \data_out_5_am[16]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_16, B => line_2_16, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[16]_net_1\);
    
    \data_out_4_i_m2_ns[19]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_i_m2_bm[19]_net_1\, C => 
        \data_out_4_i_m2_am[19]_net_1\, Y => N_74);
    
    \data_out_4_ns[21]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[21]_net_1\, C => \data_out_4_am[21]_net_1\, 
        Y => N_520);
    
    \data_out_4_am[5]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_5, B => line_2_5, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[5]_net_1\);
    
    \data_out_4_bm[4]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_4_d0, B => line_0_4, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[4]_net_1\);
    
    \data_out_4_am[9]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_9, B => line_2_9, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[9]_net_1\);
    
    \data_out_i_m2_ns_1[12]\ : CFG4
      generic map(INIT => x"46CE")

      port map(A => result_addr_net_0(1), B => 
        \data_out_i_m2_ns_1_1_1[12]_net_1\, C => line_3_12, D => 
        line_4_12, Y => \data_out_i_m2_ns_1[12]_net_1\);
    
    \data_out_5_ns[2]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_5_bm[2]_net_1\, C => \data_out_5_am[2]_net_1\, 
        Y => N_533);
    
    \data_out_4_ns[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[1]_net_1\, C => \data_out_4_am[1]_net_1\, 
        Y => N_500);
    
    \data_out_6[0]\ : CFG4
      generic map(INIT => x"D850")

      port map(A => result_addr_net_0(3), B => line_7_0, C => 
        N_531, D => ren_pos, Y => N_565);
    
    \data_out_5_am[26]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_26, B => line_6_26, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[26]_net_1\);
    
    \data_out_5_bm[5]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_5, B => line_4_5, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[5]_net_1\);
    
    \data_out_6[17]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[17]_net_1\, D
         => \data_out_5_am[17]_net_1\, Y => N_582);
    
    \data_out_4_i_m2_am[19]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_19, B => line_6_19, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_i_m2_am[19]_net_1\);
    
    \data_out_5_bm[9]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_9, B => line_4_9, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[9]_net_1\);
    
    \data_out_5_am[18]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_18, B => line_6_18, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[18]_net_1\);
    
    \data_out_6_i_RNO_0[8]\ : CFG4
      generic map(INIT => x"350F")

      port map(A => line_1_8, B => line_2_8, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \data_out_6_i_m2_1_1[8]\);
    
    \data_out_4_ns[30]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[30]_net_1\, C => \data_out_4_am[30]_net_1\, 
        Y => N_529);
    
    \data_out_i_m2_ns_1_1_1[22]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_22, B => line_6_22, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \data_out_i_m2_ns_1_1_1[22]_net_1\);
    
    \data_out_4_bm[13]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_13, B => line_0_13, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[13]_net_1\);
    
    \data_out_4_am[0]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_0, B => line_2_0, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[0]_net_1\);
    
    \data_out_6[14]\ : CFG4
      generic map(INIT => x"5140")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(1), C => \data_out_5_bm[14]_net_1\, D
         => \data_out_5_am[14]_net_1\, Y => N_579);
    
    \data_out_4_bm[6]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_6_d0, B => line_0_6, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[6]_net_1\);
    
    \data_out_4_ns[17]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[17]_net_1\, C => \data_out_4_am[17]_net_1\, 
        Y => N_516);
    
    \data_out_i_m2_ns_RNO[22]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => result_addr_net_0(1), B => 
        \data_out_i_m2_4_1_1[22]\, C => line_22, D => line_0_22, 
        Y => N_83);
    
    \data_out_i_m2_ns[22]\ : CFG4
      generic map(INIT => x"1D0C")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(0), C => \data_out_i_m2_ns_1[22]_net_1\, 
        D => N_83, Y => N_96);
    
    \data_out_5_am[30]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_30, B => line_2_30, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[30]_net_1\);
    
    \data_out_6[2]\ : CFG4
      generic map(INIT => x"D850")

      port map(A => result_addr_net_0(3), B => line_7_2, C => 
        N_533, D => ren_pos, Y => N_567);
    
    \data_out_5_bm[30]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_30, B => line_0_30, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[30]_net_1\);
    
    \data_out_5_bm[0]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_0, B => line_4_0, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[0]_net_1\);
    
    \data_out_4_am[14]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_14, B => line_2_14, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[14]_net_1\);
    
    \data_out_4_am[2]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_2, B => line_2_2, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[2]_net_1\);
    
    \data_out_4_bm[23]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_23, B => line_4_23, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[23]_net_1\);
    
    \data_out_4_ns[27]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[27]_net_1\, C => \data_out_4_am[27]_net_1\, 
        Y => N_526);
    
    \data_out_5_am[5]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_5, B => line_6_5, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[5]_net_1\);
    
    \data_out_i_m2_ns[12]\ : CFG4
      generic map(INIT => x"1D0C")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(0), C => \data_out_i_m2_ns_1[12]_net_1\, 
        D => N_68, Y => N_81);
    
    \data_out_5_am[9]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_9, B => line_6_9, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[9]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32 is

    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H0_o            : in    std_logic_vector(31 downto 0);
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic;
          wen_or                         : out   std_logic;
          SHA256_Module_0_data_out_ready : in    std_logic;
          ren_pos                        : out   std_logic;
          AHB_slave_dummy_0_read_en      : in    std_logic;
          SHA256_Module_0_do_valid_o     : in    std_logic;
          prev_sig                       : in    std_logic;
          limiter_1cycle_0_sig_1cycle    : out   std_logic
        );

end reg_1x32;

architecture DEF_ARCH of reg_1x32 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \wen_or\, GND_net_1, ren_pos_0, 
        \limiter_1cycle_0_sig_1cycle\ : std_logic;

begin 

    wen_or <= \wen_or\;
    limiter_1cycle_0_sig_1cycle <= \limiter_1cycle_0_sig_1cycle\;

    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(17));
    
    wen_or_0 : CFG2
      generic map(INIT => x"B")

      port map(A => \limiter_1cycle_0_sig_1cycle\, B => 
        SHA256_Module_0_data_out_ready, Y => \wen_or\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(18));
    
    \ren_pos\ : SLE
      port map(D => ren_pos_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ren_pos);
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(29));
    
    wen_or_0_a2 : CFG2
      generic map(INIT => x"2")

      port map(A => SHA256_Module_0_do_valid_o, B => prev_sig, Y
         => \limiter_1cycle_0_sig_1cycle\);
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(7));
    
    ren_pos_r : CFG2
      generic map(INIT => x"8")

      port map(A => SHA256_Module_0_data_out_ready, B => 
        AHB_slave_dummy_0_read_en, Y => ren_pos_0);
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \wen_or\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_7 is

    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o            : in    std_logic_vector(31 downto 0);
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic;
          wen_or                         : in    std_logic;
          SHA256_Module_0_data_out_ready : in    std_logic
        );

end reg_1x32_7;

architecture DEF_ARCH of reg_1x32_7 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_6 is

    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o            : in    std_logic_vector(31 downto 0);
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic;
          wen_or                         : in    std_logic;
          SHA256_Module_0_data_out_ready : in    std_logic
        );

end reg_1x32_6;

architecture DEF_ARCH of reg_1x32_6 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_5 is

    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o            : in    std_logic_vector(31 downto 0);
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic;
          wen_or                         : in    std_logic;
          SHA256_Module_0_data_out_ready : in    std_logic
        );

end reg_1x32_5;

architecture DEF_ARCH of reg_1x32_5 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_2 is

    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o            : in    std_logic_vector(31 downto 0);
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic;
          wen_or                         : in    std_logic;
          SHA256_Module_0_data_out_ready : in    std_logic
        );

end reg_1x32_2;

architecture DEF_ARCH of reg_1x32_2 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_0 is

    port( line_2                                    : out   std_logic;
          line_1                                    : out   std_logic;
          line_0                                    : out   std_logic;
          line_28                                   : out   std_logic;
          line_20                                   : out   std_logic;
          line_19                                   : out   std_logic;
          line_11                                   : out   std_logic;
          line_10                                   : out   std_logic;
          line_8                                    : out   std_logic;
          line_7                                    : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK              : in    std_logic;
          SHA256_Module_0_error_o                   : in    std_logic;
          wen_or                                    : in    std_logic;
          SHA256_Module_0_data_out_ready            : in    std_logic;
          SHA256_Module_0_di_req_o                  : in    std_logic;
          SHA256_Module_0_do_valid_o                : in    std_logic;
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic;
          limiter_1cycle_0_sig_1cycle               : in    std_logic
        );

end reg_1x32_0;

architecture DEF_ARCH of reg_1x32_0 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1, \line_28\, line_5, \line_20\, 
        line_4, \line_19\, line_3, \line_11\, line_2_0, \line_10\, 
        line_1_0, \line_8\, line_0_0, \line_7\, line, 
        \SHA256_Module_0_data_available_lastbank_8\, 
        \data_available\ : std_logic;

begin 

    line_28 <= \line_28\;
    line_20 <= \line_20\;
    line_19 <= \line_19\;
    line_11 <= \line_11\;
    line_10 <= \line_10\;
    line_8 <= \line_8\;
    line_7 <= \line_7\;
    SHA256_Module_0_data_available_lastbank_8 <= 
        \SHA256_Module_0_data_available_lastbank_8\;

    \line_r[28]\ : CFG3
      generic map(INIT => x"20")

      port map(A => SHA256_Module_0_data_out_ready, B => 
        limiter_1cycle_0_sig_1cycle, C => \line_28\, Y => line_5);
    
    data_available : SLE
      port map(D => \data_available\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_Module_0_data_available_lastbank_8\);
    
    \line_r[19]\ : CFG3
      generic map(INIT => x"20")

      port map(A => SHA256_Module_0_data_out_ready, B => 
        limiter_1cycle_0_sig_1cycle, C => \line_19\, Y => line_3);
    
    \line[28]\ : SLE
      port map(D => line_5, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \line_28\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[1]\ : SLE
      port map(D => SHA256_Module_0_di_req_o, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line_1);
    
    \line_r[11]\ : CFG3
      generic map(INIT => x"20")

      port map(A => SHA256_Module_0_data_out_ready, B => 
        limiter_1cycle_0_sig_1cycle, C => \line_11\, Y => 
        line_2_0);
    
    \line[7]\ : SLE
      port map(D => line, CLK => sha256_system_sb_0_FIC_0_CLK, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \line_7\);
    
    \line[19]\ : SLE
      port map(D => line_3, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \line_19\);
    
    \line[20]\ : SLE
      port map(D => line_4, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \line_20\);
    
    \line_r[20]\ : CFG3
      generic map(INIT => x"20")

      port map(A => SHA256_Module_0_data_out_ready, B => 
        limiter_1cycle_0_sig_1cycle, C => \line_20\, Y => line_4);
    
    \line[0]\ : SLE
      port map(D => SHA256_Module_0_do_valid_o, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line_r[8]\ : CFG3
      generic map(INIT => x"20")

      port map(A => SHA256_Module_0_data_out_ready, B => 
        limiter_1cycle_0_sig_1cycle, C => \line_8\, Y => line_0_0);
    
    \line[2]\ : SLE
      port map(D => SHA256_Module_0_error_o, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line_2);
    
    \line_r[10]\ : CFG3
      generic map(INIT => x"20")

      port map(A => SHA256_Module_0_data_out_ready, B => 
        limiter_1cycle_0_sig_1cycle, C => \line_10\, Y => 
        line_1_0);
    
    \line[11]\ : SLE
      port map(D => line_2_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \line_11\);
    
    \line[8]\ : SLE
      port map(D => line_0_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \line_8\);
    
    \line[10]\ : SLE
      port map(D => line_1_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \line_10\);
    
    data_available_r : CFG3
      generic map(INIT => x"A8")

      port map(A => SHA256_Module_0_data_out_ready, B => 
        limiter_1cycle_0_sig_1cycle, C => 
        \SHA256_Module_0_data_available_lastbank_8\, Y => 
        \data_available\);
    
    \line_r[7]\ : CFG3
      generic map(INIT => x"20")

      port map(A => SHA256_Module_0_data_out_ready, B => 
        limiter_1cycle_0_sig_1cycle, C => \line_7\, Y => line);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_3 is

    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o            : in    std_logic_vector(31 downto 0);
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic;
          wen_or                         : in    std_logic;
          SHA256_Module_0_data_out_ready : in    std_logic
        );

end reg_1x32_3;

architecture DEF_ARCH of reg_1x32_3 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_4 is

    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o            : in    std_logic_vector(31 downto 0);
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic;
          wen_or                         : in    std_logic;
          SHA256_Module_0_data_out_ready : in    std_logic
        );

end reg_1x32_4;

architecture DEF_ARCH of reg_1x32_4 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(12), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(23), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(10), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(26), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(31), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(15), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(19), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(14), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(5), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(22), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(20), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(17), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(18), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(4), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(25), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(30), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(29), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(11), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(24), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(9), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(13), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(27), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(16), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(8), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(28), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(7), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(21), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(6), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => wen_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        SHA256_Module_0_data_out_ready, SD => GND_net_1, LAT => 
        GND_net_1, Q => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg9_1x32 is

    port( result_addr_net_0                         : in    std_logic_vector(3 downto 0);
          SHA256_BLOCK_0_H0_o                       : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o                       : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o                       : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o                       : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o                       : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o                       : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o                       : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o                       : in    std_logic_vector(31 downto 0);
          line_7_d0                                 : out   std_logic;
          line_10                                   : out   std_logic;
          line_11                                   : out   std_logic;
          line_20                                   : out   std_logic;
          line_28                                   : out   std_logic;
          line_31                                   : out   std_logic;
          line_0_7                                  : out   std_logic;
          line_0_10                                 : out   std_logic;
          line_0_11                                 : out   std_logic;
          line_0_20                                 : out   std_logic;
          line_0_28                                 : out   std_logic;
          line_0_31                                 : out   std_logic;
          line_1_7                                  : out   std_logic;
          line_1_10                                 : out   std_logic;
          line_1_11                                 : out   std_logic;
          line_1_20                                 : out   std_logic;
          line_1_28                                 : out   std_logic;
          line_1_31                                 : out   std_logic;
          line_2_7                                  : out   std_logic;
          line_2_10                                 : out   std_logic;
          line_2_11                                 : out   std_logic;
          line_2_20                                 : out   std_logic;
          line_2_28                                 : out   std_logic;
          line_2_31                                 : out   std_logic;
          line_3_7                                  : out   std_logic;
          line_3_10                                 : out   std_logic;
          line_3_11                                 : out   std_logic;
          line_3_20                                 : out   std_logic;
          line_3_28                                 : out   std_logic;
          line_3_31                                 : out   std_logic;
          line_4_7                                  : out   std_logic;
          line_4_10                                 : out   std_logic;
          line_4_11                                 : out   std_logic;
          line_4_20                                 : out   std_logic;
          line_4_28                                 : out   std_logic;
          line_4_31                                 : out   std_logic;
          line_5_7                                  : out   std_logic;
          line_5_10                                 : out   std_logic;
          line_5_11                                 : out   std_logic;
          line_5_20                                 : out   std_logic;
          line_5_28                                 : out   std_logic;
          line_5_31                                 : out   std_logic;
          line_6_7                                  : out   std_logic;
          line_6_10                                 : out   std_logic;
          line_6_11                                 : out   std_logic;
          line_6_20                                 : out   std_logic;
          line_6_28                                 : out   std_logic;
          line_6_31                                 : out   std_logic;
          line_7_28                                 : out   std_logic;
          line_7_20                                 : out   std_logic;
          line_7_11                                 : out   std_logic;
          line_7_10                                 : out   std_logic;
          line_7_7                                  : out   std_logic;
          N_568                                     : out   std_logic;
          N_579                                     : out   std_logic;
          N_580                                     : out   std_logic;
          N_581                                     : out   std_logic;
          N_583                                     : out   std_logic;
          N_588                                     : out   std_logic;
          N_589                                     : out   std_logic;
          N_590                                     : out   std_logic;
          N_591                                     : out   std_logic;
          N_592                                     : out   std_logic;
          N_595                                     : out   std_logic;
          N_594                                     : out   std_logic;
          N_586                                     : out   std_logic;
          N_582                                     : out   std_logic;
          N_578                                     : out   std_logic;
          N_574                                     : out   std_logic;
          N_571                                     : out   std_logic;
          N_570                                     : out   std_logic;
          N_569                                     : out   std_logic;
          N_96                                      : out   std_logic;
          N_81                                      : out   std_logic;
          N_74                                      : out   std_logic;
          N_75                                      : out   std_logic;
          N_499                                     : out   std_logic;
          N_501                                     : out   std_logic;
          N_525                                     : out   std_logic;
          N_513                                     : out   std_logic;
          N_502                                     : out   std_logic;
          N_522                                     : out   std_logic;
          N_500                                     : out   std_logic;
          N_514                                     : out   std_logic;
          N_515                                     : out   std_logic;
          N_524                                     : out   std_logic;
          N_526                                     : out   std_logic;
          N_529                                     : out   std_logic;
          N_528                                     : out   std_logic;
          N_523                                     : out   std_logic;
          N_517                                     : out   std_logic;
          N_505                                     : out   std_logic;
          N_503                                     : out   std_logic;
          N_512                                     : out   std_logic;
          N_508                                     : out   std_logic;
          N_504                                     : out   std_logic;
          N_520                                     : out   std_logic;
          N_516                                     : out   std_logic;
          ren_pos                                   : out   std_logic;
          N_228                                     : out   std_logic;
          N_7                                       : out   std_logic;
          N_566                                     : out   std_logic;
          N_567                                     : out   std_logic;
          N_565                                     : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK              : in    std_logic;
          SHA256_Module_0_data_out_ready            : in    std_logic;
          AHB_slave_dummy_0_read_en                 : in    std_logic;
          SHA256_Module_0_do_valid_o                : in    std_logic;
          prev_sig                                  : in    std_logic;
          SHA256_Module_0_error_o                   : in    std_logic;
          SHA256_Module_0_di_req_o                  : in    std_logic;
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic
        );

end reg9_1x32;

architecture DEF_ARCH of reg9_1x32 is 

  component reg_1x32_1
    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o            : in    std_logic_vector(31 downto 0) := (others => 'U');
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          wen_or                         : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready : in    std_logic := 'U'
        );
  end component;

  component mux_9_1
    port( result_addr_net_0 : in    std_logic_vector(3 downto 0) := (others => 'U');
          line_19           : in    std_logic := 'U';
          line_22           : in    std_logic := 'U';
          line_12           : in    std_logic := 'U';
          line_8            : in    std_logic := 'U';
          line_17           : in    std_logic := 'U';
          line_21           : in    std_logic := 'U';
          line_5_d0         : in    std_logic := 'U';
          line_9            : in    std_logic := 'U';
          line_13           : in    std_logic := 'U';
          line_4_d0         : in    std_logic := 'U';
          line_6_d0         : in    std_logic := 'U';
          line_18           : in    std_logic := 'U';
          line_24           : in    std_logic := 'U';
          line_29           : in    std_logic := 'U';
          line_30           : in    std_logic := 'U';
          line_27           : in    std_logic := 'U';
          line_25           : in    std_logic := 'U';
          line_16           : in    std_logic := 'U';
          line_15           : in    std_logic := 'U';
          line_1_d0         : in    std_logic := 'U';
          line_23           : in    std_logic := 'U';
          line_3_d0         : in    std_logic := 'U';
          line_14           : in    std_logic := 'U';
          line_26           : in    std_logic := 'U';
          line_2_d0         : in    std_logic := 'U';
          line_0_d0         : in    std_logic := 'U';
          line_0_19         : in    std_logic := 'U';
          line_0_22         : in    std_logic := 'U';
          line_0_12         : in    std_logic := 'U';
          line_0_8          : in    std_logic := 'U';
          line_0_17         : in    std_logic := 'U';
          line_0_21         : in    std_logic := 'U';
          line_0_5          : in    std_logic := 'U';
          line_0_9          : in    std_logic := 'U';
          line_0_13         : in    std_logic := 'U';
          line_0_4          : in    std_logic := 'U';
          line_0_6          : in    std_logic := 'U';
          line_0_18         : in    std_logic := 'U';
          line_0_24         : in    std_logic := 'U';
          line_0_29         : in    std_logic := 'U';
          line_0_30         : in    std_logic := 'U';
          line_0_27         : in    std_logic := 'U';
          line_0_25         : in    std_logic := 'U';
          line_0_16         : in    std_logic := 'U';
          line_0_15         : in    std_logic := 'U';
          line_0_1          : in    std_logic := 'U';
          line_0_23         : in    std_logic := 'U';
          line_0_3          : in    std_logic := 'U';
          line_0_14         : in    std_logic := 'U';
          line_0_26         : in    std_logic := 'U';
          line_0_2          : in    std_logic := 'U';
          line_0_0          : in    std_logic := 'U';
          line_1_19         : in    std_logic := 'U';
          line_1_22         : in    std_logic := 'U';
          line_1_12         : in    std_logic := 'U';
          line_1_8          : in    std_logic := 'U';
          line_1_17         : in    std_logic := 'U';
          line_1_21         : in    std_logic := 'U';
          line_1_5          : in    std_logic := 'U';
          line_1_9          : in    std_logic := 'U';
          line_1_13         : in    std_logic := 'U';
          line_1_4          : in    std_logic := 'U';
          line_1_6          : in    std_logic := 'U';
          line_1_18         : in    std_logic := 'U';
          line_1_24         : in    std_logic := 'U';
          line_1_29         : in    std_logic := 'U';
          line_1_30         : in    std_logic := 'U';
          line_1_27         : in    std_logic := 'U';
          line_1_25         : in    std_logic := 'U';
          line_1_16         : in    std_logic := 'U';
          line_1_15         : in    std_logic := 'U';
          line_1_1          : in    std_logic := 'U';
          line_1_23         : in    std_logic := 'U';
          line_1_3          : in    std_logic := 'U';
          line_1_14         : in    std_logic := 'U';
          line_1_26         : in    std_logic := 'U';
          line_1_2          : in    std_logic := 'U';
          line_1_0          : in    std_logic := 'U';
          line_2_19         : in    std_logic := 'U';
          line_2_22         : in    std_logic := 'U';
          line_2_12         : in    std_logic := 'U';
          line_2_8          : in    std_logic := 'U';
          line_2_17         : in    std_logic := 'U';
          line_2_21         : in    std_logic := 'U';
          line_2_5          : in    std_logic := 'U';
          line_2_9          : in    std_logic := 'U';
          line_2_13         : in    std_logic := 'U';
          line_2_4          : in    std_logic := 'U';
          line_2_6          : in    std_logic := 'U';
          line_2_18         : in    std_logic := 'U';
          line_2_24         : in    std_logic := 'U';
          line_2_29         : in    std_logic := 'U';
          line_2_30         : in    std_logic := 'U';
          line_2_27         : in    std_logic := 'U';
          line_2_25         : in    std_logic := 'U';
          line_2_16         : in    std_logic := 'U';
          line_2_15         : in    std_logic := 'U';
          line_2_1          : in    std_logic := 'U';
          line_2_23         : in    std_logic := 'U';
          line_2_3          : in    std_logic := 'U';
          line_2_14         : in    std_logic := 'U';
          line_2_26         : in    std_logic := 'U';
          line_2_2          : in    std_logic := 'U';
          line_2_0          : in    std_logic := 'U';
          line_3_22         : in    std_logic := 'U';
          line_3_12         : in    std_logic := 'U';
          line_3_4          : in    std_logic := 'U';
          line_3_6          : in    std_logic := 'U';
          line_3_29         : in    std_logic := 'U';
          line_3_24         : in    std_logic := 'U';
          line_3_30         : in    std_logic := 'U';
          line_3_27         : in    std_logic := 'U';
          line_3_25         : in    std_logic := 'U';
          line_3_16         : in    std_logic := 'U';
          line_3_15         : in    std_logic := 'U';
          line_3_1          : in    std_logic := 'U';
          line_3_18         : in    std_logic := 'U';
          line_3_13         : in    std_logic := 'U';
          line_3_9          : in    std_logic := 'U';
          line_3_5          : in    std_logic := 'U';
          line_3_23         : in    std_logic := 'U';
          line_3_21         : in    std_logic := 'U';
          line_3_17         : in    std_logic := 'U';
          line_3_3          : in    std_logic := 'U';
          line_3_14         : in    std_logic := 'U';
          line_3_26         : in    std_logic := 'U';
          line_3_2          : in    std_logic := 'U';
          line_3_0          : in    std_logic := 'U';
          line_3_8          : in    std_logic := 'U';
          line_3_19         : in    std_logic := 'U';
          line_4_22         : in    std_logic := 'U';
          line_4_12         : in    std_logic := 'U';
          line_4_4          : in    std_logic := 'U';
          line_4_6          : in    std_logic := 'U';
          line_4_29         : in    std_logic := 'U';
          line_4_24         : in    std_logic := 'U';
          line_4_30         : in    std_logic := 'U';
          line_4_27         : in    std_logic := 'U';
          line_4_25         : in    std_logic := 'U';
          line_4_16         : in    std_logic := 'U';
          line_4_15         : in    std_logic := 'U';
          line_4_1          : in    std_logic := 'U';
          line_4_18         : in    std_logic := 'U';
          line_4_13         : in    std_logic := 'U';
          line_4_9          : in    std_logic := 'U';
          line_4_5          : in    std_logic := 'U';
          line_4_23         : in    std_logic := 'U';
          line_4_21         : in    std_logic := 'U';
          line_4_17         : in    std_logic := 'U';
          line_4_3          : in    std_logic := 'U';
          line_4_14         : in    std_logic := 'U';
          line_4_26         : in    std_logic := 'U';
          line_4_2          : in    std_logic := 'U';
          line_4_0          : in    std_logic := 'U';
          line_4_8          : in    std_logic := 'U';
          line_4_19         : in    std_logic := 'U';
          line_5_22         : in    std_logic := 'U';
          line_5_12         : in    std_logic := 'U';
          line_5_4          : in    std_logic := 'U';
          line_5_6          : in    std_logic := 'U';
          line_5_29         : in    std_logic := 'U';
          line_5_24         : in    std_logic := 'U';
          line_5_30         : in    std_logic := 'U';
          line_5_27         : in    std_logic := 'U';
          line_5_25         : in    std_logic := 'U';
          line_5_16         : in    std_logic := 'U';
          line_5_15         : in    std_logic := 'U';
          line_5_1          : in    std_logic := 'U';
          line_5_18         : in    std_logic := 'U';
          line_5_13         : in    std_logic := 'U';
          line_5_9          : in    std_logic := 'U';
          line_5_5          : in    std_logic := 'U';
          line_5_23         : in    std_logic := 'U';
          line_5_21         : in    std_logic := 'U';
          line_5_17         : in    std_logic := 'U';
          line_5_3          : in    std_logic := 'U';
          line_5_14         : in    std_logic := 'U';
          line_5_26         : in    std_logic := 'U';
          line_5_2          : in    std_logic := 'U';
          line_5_0          : in    std_logic := 'U';
          line_5_8          : in    std_logic := 'U';
          line_5_19         : in    std_logic := 'U';
          line_6_22         : in    std_logic := 'U';
          line_6_12         : in    std_logic := 'U';
          line_6_4          : in    std_logic := 'U';
          line_6_6          : in    std_logic := 'U';
          line_6_29         : in    std_logic := 'U';
          line_6_24         : in    std_logic := 'U';
          line_6_30         : in    std_logic := 'U';
          line_6_27         : in    std_logic := 'U';
          line_6_25         : in    std_logic := 'U';
          line_6_16         : in    std_logic := 'U';
          line_6_15         : in    std_logic := 'U';
          line_6_1          : in    std_logic := 'U';
          line_6_18         : in    std_logic := 'U';
          line_6_13         : in    std_logic := 'U';
          line_6_9          : in    std_logic := 'U';
          line_6_5          : in    std_logic := 'U';
          line_6_23         : in    std_logic := 'U';
          line_6_21         : in    std_logic := 'U';
          line_6_17         : in    std_logic := 'U';
          line_6_3          : in    std_logic := 'U';
          line_6_14         : in    std_logic := 'U';
          line_6_26         : in    std_logic := 'U';
          line_6_2          : in    std_logic := 'U';
          line_6_0          : in    std_logic := 'U';
          line_6_8          : in    std_logic := 'U';
          line_6_19         : in    std_logic := 'U';
          line_7_19         : in    std_logic := 'U';
          line_7_8          : in    std_logic := 'U';
          line_7_1          : in    std_logic := 'U';
          line_7_2          : in    std_logic := 'U';
          line_7_0          : in    std_logic := 'U';
          N_568             : out   std_logic;
          N_579             : out   std_logic;
          N_580             : out   std_logic;
          N_581             : out   std_logic;
          N_583             : out   std_logic;
          N_588             : out   std_logic;
          N_589             : out   std_logic;
          N_590             : out   std_logic;
          N_591             : out   std_logic;
          N_592             : out   std_logic;
          N_595             : out   std_logic;
          N_594             : out   std_logic;
          N_586             : out   std_logic;
          N_582             : out   std_logic;
          N_578             : out   std_logic;
          N_574             : out   std_logic;
          N_571             : out   std_logic;
          N_570             : out   std_logic;
          N_569             : out   std_logic;
          N_96              : out   std_logic;
          N_81              : out   std_logic;
          N_74              : out   std_logic;
          N_75              : out   std_logic;
          N_499             : out   std_logic;
          N_501             : out   std_logic;
          N_525             : out   std_logic;
          N_513             : out   std_logic;
          N_502             : out   std_logic;
          N_522             : out   std_logic;
          N_500             : out   std_logic;
          N_514             : out   std_logic;
          N_515             : out   std_logic;
          N_524             : out   std_logic;
          N_526             : out   std_logic;
          N_529             : out   std_logic;
          N_528             : out   std_logic;
          N_523             : out   std_logic;
          N_517             : out   std_logic;
          N_505             : out   std_logic;
          N_503             : out   std_logic;
          N_512             : out   std_logic;
          N_508             : out   std_logic;
          N_504             : out   std_logic;
          N_520             : out   std_logic;
          N_516             : out   std_logic;
          ren_pos           : in    std_logic := 'U';
          N_228             : out   std_logic;
          N_7               : out   std_logic;
          N_566             : out   std_logic;
          N_567             : out   std_logic;
          N_565             : out   std_logic
        );
  end component;

  component reg_1x32
    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H0_o            : in    std_logic_vector(31 downto 0) := (others => 'U');
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          wen_or                         : out   std_logic;
          SHA256_Module_0_data_out_ready : in    std_logic := 'U';
          ren_pos                        : out   std_logic;
          AHB_slave_dummy_0_read_en      : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o     : in    std_logic := 'U';
          prev_sig                       : in    std_logic := 'U';
          limiter_1cycle_0_sig_1cycle    : out   std_logic
        );
  end component;

  component reg_1x32_7
    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o            : in    std_logic_vector(31 downto 0) := (others => 'U');
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          wen_or                         : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_6
    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o            : in    std_logic_vector(31 downto 0) := (others => 'U');
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          wen_or                         : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component reg_1x32_5
    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o            : in    std_logic_vector(31 downto 0) := (others => 'U');
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          wen_or                         : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_2
    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o            : in    std_logic_vector(31 downto 0) := (others => 'U');
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          wen_or                         : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_0
    port( line_2                                    : out   std_logic;
          line_1                                    : out   std_logic;
          line_0                                    : out   std_logic;
          line_28                                   : out   std_logic;
          line_20                                   : out   std_logic;
          line_19                                   : out   std_logic;
          line_11                                   : out   std_logic;
          line_10                                   : out   std_logic;
          line_8                                    : out   std_logic;
          line_7                                    : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK              : in    std_logic := 'U';
          SHA256_Module_0_error_o                   : in    std_logic := 'U';
          wen_or                                    : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready            : in    std_logic := 'U';
          SHA256_Module_0_di_req_o                  : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o                : in    std_logic := 'U';
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic;
          limiter_1cycle_0_sig_1cycle               : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_3
    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o            : in    std_logic_vector(31 downto 0) := (others => 'U');
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          wen_or                         : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_4
    port( line                           : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o            : in    std_logic_vector(31 downto 0) := (others => 'U');
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          wen_or                         : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready : in    std_logic := 'U'
        );
  end component;

    signal \line[19]\, \line[22]\, \line[12]\, \line[8]\, 
        \line[17]\, \line[21]\, \line[5]\, \line[9]\, \line[13]\, 
        \line[4]\, \line[6]\, \line[18]\, \line[24]\, \line[29]\, 
        \line[30]\, \line[27]\, \line[25]\, \line[16]\, 
        \line[15]\, \line[1]\, \line[23]\, \line[3]\, \line[14]\, 
        \line[26]\, \line[2]\, \line[0]\, \line_0[19]\, 
        \line_0[22]\, \line_0[12]\, \line_0[8]\, \line_0[17]\, 
        \line_0[21]\, \line_0[5]\, \line_0[9]\, \line_0[13]\, 
        \line_0[4]\, \line_0[6]\, \line_0[18]\, \line_0[24]\, 
        \line_0[29]\, \line_0[30]\, \line_0[27]\, \line_0[25]\, 
        \line_0[16]\, \line_0[15]\, \line_0[1]\, \line_0[23]\, 
        \line_0[3]\, \line_0[14]\, \line_0[26]\, \line_0[2]\, 
        \line_0[0]\, \line_1[19]\, \line_1[22]\, \line_1[12]\, 
        \line_1[8]\, \line_1[17]\, \line_1[21]\, \line_1[5]\, 
        \line_1[9]\, \line_1[13]\, \line_1[4]\, \line_1[6]\, 
        \line_1[18]\, \line_1[24]\, \line_1[29]\, \line_1[30]\, 
        \line_1[27]\, \line_1[25]\, \line_1[16]\, \line_1[15]\, 
        \line_1[1]\, \line_1[23]\, \line_1[3]\, \line_1[14]\, 
        \line_1[26]\, \line_1[2]\, \line_1[0]\, \line_2[19]\, 
        \line_2[22]\, \line_2[12]\, \line_2[8]\, \line_2[17]\, 
        \line_2[21]\, \line_2[5]\, \line_2[9]\, \line_2[13]\, 
        \line_2[4]\, \line_2[6]\, \line_2[18]\, \line_2[24]\, 
        \line_2[29]\, \line_2[30]\, \line_2[27]\, \line_2[25]\, 
        \line_2[16]\, \line_2[15]\, \line_2[1]\, \line_2[23]\, 
        \line_2[3]\, \line_2[14]\, \line_2[26]\, \line_2[2]\, 
        \line_2[0]\, \line_3[22]\, \line_3[12]\, \line_3[4]\, 
        \line_3[6]\, \line_3[29]\, \line_3[24]\, \line_3[30]\, 
        \line_3[27]\, \line_3[25]\, \line_3[16]\, \line_3[15]\, 
        \line_3[1]\, \line_3[18]\, \line_3[13]\, \line_3[9]\, 
        \line_3[5]\, \line_3[23]\, \line_3[21]\, \line_3[17]\, 
        \line_3[3]\, \line_3[14]\, \line_3[26]\, \line_3[2]\, 
        \line_3[0]\, \line_3[8]\, \line_3[19]\, \line_4[22]\, 
        \line_4[12]\, \line_4[4]\, \line_4[6]\, \line_4[29]\, 
        \line_4[24]\, \line_4[30]\, \line_4[27]\, \line_4[25]\, 
        \line_4[16]\, \line_4[15]\, \line_4[1]\, \line_4[18]\, 
        \line_4[13]\, \line_4[9]\, \line_4[5]\, \line_4[23]\, 
        \line_4[21]\, \line_4[17]\, \line_4[3]\, \line_4[14]\, 
        \line_4[26]\, \line_4[2]\, \line_4[0]\, \line_4[8]\, 
        \line_4[19]\, \line_5[22]\, \line_5[12]\, \line_5[4]\, 
        \line_5[6]\, \line_5[29]\, \line_5[24]\, \line_5[30]\, 
        \line_5[27]\, \line_5[25]\, \line_5[16]\, \line_5[15]\, 
        \line_5[1]\, \line_5[18]\, \line_5[13]\, \line_5[9]\, 
        \line_5[5]\, \line_5[23]\, \line_5[21]\, \line_5[17]\, 
        \line_5[3]\, \line_5[14]\, \line_5[26]\, \line_5[2]\, 
        \line_5[0]\, \line_5[8]\, \line_5[19]\, \line_6[22]\, 
        \line_6[12]\, \line_6[4]\, \line_6[6]\, \line_6[29]\, 
        \line_6[24]\, \line_6[30]\, \line_6[27]\, \line_6[25]\, 
        \line_6[16]\, \line_6[15]\, \line_6[1]\, \line_6[18]\, 
        \line_6[13]\, \line_6[9]\, \line_6[5]\, \line_6[23]\, 
        \line_6[21]\, \line_6[17]\, \line_6[3]\, \line_6[14]\, 
        \line_6[26]\, \line_6[2]\, \line_6[0]\, \line_6[8]\, 
        \line_6[19]\, \line_7[19]\, \line_7[8]\, \line_7[1]\, 
        \line_7[2]\, \line_7[0]\, \ren_pos\, wen_or, 
        limiter_1cycle_0_sig_1cycle, GND_net_1, VCC_net_1
         : std_logic;

    for all : reg_1x32_1
	Use entity work.reg_1x32_1(DEF_ARCH);
    for all : mux_9_1
	Use entity work.mux_9_1(DEF_ARCH);
    for all : reg_1x32
	Use entity work.reg_1x32(DEF_ARCH);
    for all : reg_1x32_7
	Use entity work.reg_1x32_7(DEF_ARCH);
    for all : reg_1x32_6
	Use entity work.reg_1x32_6(DEF_ARCH);
    for all : reg_1x32_5
	Use entity work.reg_1x32_5(DEF_ARCH);
    for all : reg_1x32_2
	Use entity work.reg_1x32_2(DEF_ARCH);
    for all : reg_1x32_0
	Use entity work.reg_1x32_0(DEF_ARCH);
    for all : reg_1x32_3
	Use entity work.reg_1x32_3(DEF_ARCH);
    for all : reg_1x32_4
	Use entity work.reg_1x32_4(DEF_ARCH);
begin 

    ren_pos <= \ren_pos\;

    \reg_1x32_1\ : reg_1x32_1
      port map(line(31) => line_0_31, line(30) => \line_5[30]\, 
        line(29) => \line_1[29]\, line(28) => line_0_28, line(27)
         => \line_5[27]\, line(26) => \line_1[26]\, line(25) => 
        \line_5[25]\, line(24) => \line_1[24]\, line(23) => 
        \line_5[23]\, line(22) => \line_5[22]\, line(21) => 
        \line_1[21]\, line(20) => line_0_20, line(19) => 
        \line_5[19]\, line(18) => \line_1[18]\, line(17) => 
        \line_1[17]\, line(16) => \line_5[16]\, line(15) => 
        \line_5[15]\, line(14) => \line_1[14]\, line(13) => 
        \line_1[13]\, line(12) => \line_5[12]\, line(11) => 
        line_0_11, line(10) => line_0_10, line(9) => \line_1[9]\, 
        line(8) => \line_5[8]\, line(7) => line_0_7, line(6) => 
        \line_1[6]\, line(5) => \line_1[5]\, line(4) => 
        \line_1[4]\, line(3) => \line_1[3]\, line(2) => 
        \line_1[2]\, line(1) => \line_5[1]\, line(0) => 
        \line_1[0]\, SHA256_BLOCK_0_H1_o(31) => 
        SHA256_BLOCK_0_H1_o(31), SHA256_BLOCK_0_H1_o(30) => 
        SHA256_BLOCK_0_H1_o(30), SHA256_BLOCK_0_H1_o(29) => 
        SHA256_BLOCK_0_H1_o(29), SHA256_BLOCK_0_H1_o(28) => 
        SHA256_BLOCK_0_H1_o(28), SHA256_BLOCK_0_H1_o(27) => 
        SHA256_BLOCK_0_H1_o(27), SHA256_BLOCK_0_H1_o(26) => 
        SHA256_BLOCK_0_H1_o(26), SHA256_BLOCK_0_H1_o(25) => 
        SHA256_BLOCK_0_H1_o(25), SHA256_BLOCK_0_H1_o(24) => 
        SHA256_BLOCK_0_H1_o(24), SHA256_BLOCK_0_H1_o(23) => 
        SHA256_BLOCK_0_H1_o(23), SHA256_BLOCK_0_H1_o(22) => 
        SHA256_BLOCK_0_H1_o(22), SHA256_BLOCK_0_H1_o(21) => 
        SHA256_BLOCK_0_H1_o(21), SHA256_BLOCK_0_H1_o(20) => 
        SHA256_BLOCK_0_H1_o(20), SHA256_BLOCK_0_H1_o(19) => 
        SHA256_BLOCK_0_H1_o(19), SHA256_BLOCK_0_H1_o(18) => 
        SHA256_BLOCK_0_H1_o(18), SHA256_BLOCK_0_H1_o(17) => 
        SHA256_BLOCK_0_H1_o(17), SHA256_BLOCK_0_H1_o(16) => 
        SHA256_BLOCK_0_H1_o(16), SHA256_BLOCK_0_H1_o(15) => 
        SHA256_BLOCK_0_H1_o(15), SHA256_BLOCK_0_H1_o(14) => 
        SHA256_BLOCK_0_H1_o(14), SHA256_BLOCK_0_H1_o(13) => 
        SHA256_BLOCK_0_H1_o(13), SHA256_BLOCK_0_H1_o(12) => 
        SHA256_BLOCK_0_H1_o(12), SHA256_BLOCK_0_H1_o(11) => 
        SHA256_BLOCK_0_H1_o(11), SHA256_BLOCK_0_H1_o(10) => 
        SHA256_BLOCK_0_H1_o(10), SHA256_BLOCK_0_H1_o(9) => 
        SHA256_BLOCK_0_H1_o(9), SHA256_BLOCK_0_H1_o(8) => 
        SHA256_BLOCK_0_H1_o(8), SHA256_BLOCK_0_H1_o(7) => 
        SHA256_BLOCK_0_H1_o(7), SHA256_BLOCK_0_H1_o(6) => 
        SHA256_BLOCK_0_H1_o(6), SHA256_BLOCK_0_H1_o(5) => 
        SHA256_BLOCK_0_H1_o(5), SHA256_BLOCK_0_H1_o(4) => 
        SHA256_BLOCK_0_H1_o(4), SHA256_BLOCK_0_H1_o(3) => 
        SHA256_BLOCK_0_H1_o(3), SHA256_BLOCK_0_H1_o(2) => 
        SHA256_BLOCK_0_H1_o(2), SHA256_BLOCK_0_H1_o(1) => 
        SHA256_BLOCK_0_H1_o(1), SHA256_BLOCK_0_H1_o(0) => 
        SHA256_BLOCK_0_H1_o(0), sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, wen_or => wen_or, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready);
    
    mux_9_1_0 : mux_9_1
      port map(result_addr_net_0(3) => result_addr_net_0(3), 
        result_addr_net_0(2) => result_addr_net_0(2), 
        result_addr_net_0(1) => result_addr_net_0(1), 
        result_addr_net_0(0) => result_addr_net_0(0), line_19 => 
        \line[19]\, line_22 => \line[22]\, line_12 => \line[12]\, 
        line_8 => \line[8]\, line_17 => \line[17]\, line_21 => 
        \line[21]\, line_5_d0 => \line[5]\, line_9 => \line[9]\, 
        line_13 => \line[13]\, line_4_d0 => \line[4]\, line_6_d0
         => \line[6]\, line_18 => \line[18]\, line_24 => 
        \line[24]\, line_29 => \line[29]\, line_30 => \line[30]\, 
        line_27 => \line[27]\, line_25 => \line[25]\, line_16 => 
        \line[16]\, line_15 => \line[15]\, line_1_d0 => \line[1]\, 
        line_23 => \line[23]\, line_3_d0 => \line[3]\, line_14
         => \line[14]\, line_26 => \line[26]\, line_2_d0 => 
        \line[2]\, line_0_d0 => \line[0]\, line_0_19 => 
        \line_0[19]\, line_0_22 => \line_0[22]\, line_0_12 => 
        \line_0[12]\, line_0_8 => \line_0[8]\, line_0_17 => 
        \line_0[17]\, line_0_21 => \line_0[21]\, line_0_5 => 
        \line_0[5]\, line_0_9 => \line_0[9]\, line_0_13 => 
        \line_0[13]\, line_0_4 => \line_0[4]\, line_0_6 => 
        \line_0[6]\, line_0_18 => \line_0[18]\, line_0_24 => 
        \line_0[24]\, line_0_29 => \line_0[29]\, line_0_30 => 
        \line_0[30]\, line_0_27 => \line_0[27]\, line_0_25 => 
        \line_0[25]\, line_0_16 => \line_0[16]\, line_0_15 => 
        \line_0[15]\, line_0_1 => \line_0[1]\, line_0_23 => 
        \line_0[23]\, line_0_3 => \line_0[3]\, line_0_14 => 
        \line_0[14]\, line_0_26 => \line_0[26]\, line_0_2 => 
        \line_0[2]\, line_0_0 => \line_0[0]\, line_1_19 => 
        \line_1[19]\, line_1_22 => \line_1[22]\, line_1_12 => 
        \line_1[12]\, line_1_8 => \line_1[8]\, line_1_17 => 
        \line_1[17]\, line_1_21 => \line_1[21]\, line_1_5 => 
        \line_1[5]\, line_1_9 => \line_1[9]\, line_1_13 => 
        \line_1[13]\, line_1_4 => \line_1[4]\, line_1_6 => 
        \line_1[6]\, line_1_18 => \line_1[18]\, line_1_24 => 
        \line_1[24]\, line_1_29 => \line_1[29]\, line_1_30 => 
        \line_1[30]\, line_1_27 => \line_1[27]\, line_1_25 => 
        \line_1[25]\, line_1_16 => \line_1[16]\, line_1_15 => 
        \line_1[15]\, line_1_1 => \line_1[1]\, line_1_23 => 
        \line_1[23]\, line_1_3 => \line_1[3]\, line_1_14 => 
        \line_1[14]\, line_1_26 => \line_1[26]\, line_1_2 => 
        \line_1[2]\, line_1_0 => \line_1[0]\, line_2_19 => 
        \line_2[19]\, line_2_22 => \line_2[22]\, line_2_12 => 
        \line_2[12]\, line_2_8 => \line_2[8]\, line_2_17 => 
        \line_2[17]\, line_2_21 => \line_2[21]\, line_2_5 => 
        \line_2[5]\, line_2_9 => \line_2[9]\, line_2_13 => 
        \line_2[13]\, line_2_4 => \line_2[4]\, line_2_6 => 
        \line_2[6]\, line_2_18 => \line_2[18]\, line_2_24 => 
        \line_2[24]\, line_2_29 => \line_2[29]\, line_2_30 => 
        \line_2[30]\, line_2_27 => \line_2[27]\, line_2_25 => 
        \line_2[25]\, line_2_16 => \line_2[16]\, line_2_15 => 
        \line_2[15]\, line_2_1 => \line_2[1]\, line_2_23 => 
        \line_2[23]\, line_2_3 => \line_2[3]\, line_2_14 => 
        \line_2[14]\, line_2_26 => \line_2[26]\, line_2_2 => 
        \line_2[2]\, line_2_0 => \line_2[0]\, line_3_22 => 
        \line_3[22]\, line_3_12 => \line_3[12]\, line_3_4 => 
        \line_3[4]\, line_3_6 => \line_3[6]\, line_3_29 => 
        \line_3[29]\, line_3_24 => \line_3[24]\, line_3_30 => 
        \line_3[30]\, line_3_27 => \line_3[27]\, line_3_25 => 
        \line_3[25]\, line_3_16 => \line_3[16]\, line_3_15 => 
        \line_3[15]\, line_3_1 => \line_3[1]\, line_3_18 => 
        \line_3[18]\, line_3_13 => \line_3[13]\, line_3_9 => 
        \line_3[9]\, line_3_5 => \line_3[5]\, line_3_23 => 
        \line_3[23]\, line_3_21 => \line_3[21]\, line_3_17 => 
        \line_3[17]\, line_3_3 => \line_3[3]\, line_3_14 => 
        \line_3[14]\, line_3_26 => \line_3[26]\, line_3_2 => 
        \line_3[2]\, line_3_0 => \line_3[0]\, line_3_8 => 
        \line_3[8]\, line_3_19 => \line_3[19]\, line_4_22 => 
        \line_4[22]\, line_4_12 => \line_4[12]\, line_4_4 => 
        \line_4[4]\, line_4_6 => \line_4[6]\, line_4_29 => 
        \line_4[29]\, line_4_24 => \line_4[24]\, line_4_30 => 
        \line_4[30]\, line_4_27 => \line_4[27]\, line_4_25 => 
        \line_4[25]\, line_4_16 => \line_4[16]\, line_4_15 => 
        \line_4[15]\, line_4_1 => \line_4[1]\, line_4_18 => 
        \line_4[18]\, line_4_13 => \line_4[13]\, line_4_9 => 
        \line_4[9]\, line_4_5 => \line_4[5]\, line_4_23 => 
        \line_4[23]\, line_4_21 => \line_4[21]\, line_4_17 => 
        \line_4[17]\, line_4_3 => \line_4[3]\, line_4_14 => 
        \line_4[14]\, line_4_26 => \line_4[26]\, line_4_2 => 
        \line_4[2]\, line_4_0 => \line_4[0]\, line_4_8 => 
        \line_4[8]\, line_4_19 => \line_4[19]\, line_5_22 => 
        \line_5[22]\, line_5_12 => \line_5[12]\, line_5_4 => 
        \line_5[4]\, line_5_6 => \line_5[6]\, line_5_29 => 
        \line_5[29]\, line_5_24 => \line_5[24]\, line_5_30 => 
        \line_5[30]\, line_5_27 => \line_5[27]\, line_5_25 => 
        \line_5[25]\, line_5_16 => \line_5[16]\, line_5_15 => 
        \line_5[15]\, line_5_1 => \line_5[1]\, line_5_18 => 
        \line_5[18]\, line_5_13 => \line_5[13]\, line_5_9 => 
        \line_5[9]\, line_5_5 => \line_5[5]\, line_5_23 => 
        \line_5[23]\, line_5_21 => \line_5[21]\, line_5_17 => 
        \line_5[17]\, line_5_3 => \line_5[3]\, line_5_14 => 
        \line_5[14]\, line_5_26 => \line_5[26]\, line_5_2 => 
        \line_5[2]\, line_5_0 => \line_5[0]\, line_5_8 => 
        \line_5[8]\, line_5_19 => \line_5[19]\, line_6_22 => 
        \line_6[22]\, line_6_12 => \line_6[12]\, line_6_4 => 
        \line_6[4]\, line_6_6 => \line_6[6]\, line_6_29 => 
        \line_6[29]\, line_6_24 => \line_6[24]\, line_6_30 => 
        \line_6[30]\, line_6_27 => \line_6[27]\, line_6_25 => 
        \line_6[25]\, line_6_16 => \line_6[16]\, line_6_15 => 
        \line_6[15]\, line_6_1 => \line_6[1]\, line_6_18 => 
        \line_6[18]\, line_6_13 => \line_6[13]\, line_6_9 => 
        \line_6[9]\, line_6_5 => \line_6[5]\, line_6_23 => 
        \line_6[23]\, line_6_21 => \line_6[21]\, line_6_17 => 
        \line_6[17]\, line_6_3 => \line_6[3]\, line_6_14 => 
        \line_6[14]\, line_6_26 => \line_6[26]\, line_6_2 => 
        \line_6[2]\, line_6_0 => \line_6[0]\, line_6_8 => 
        \line_6[8]\, line_6_19 => \line_6[19]\, line_7_19 => 
        \line_7[19]\, line_7_8 => \line_7[8]\, line_7_1 => 
        \line_7[1]\, line_7_2 => \line_7[2]\, line_7_0 => 
        \line_7[0]\, N_568 => N_568, N_579 => N_579, N_580 => 
        N_580, N_581 => N_581, N_583 => N_583, N_588 => N_588, 
        N_589 => N_589, N_590 => N_590, N_591 => N_591, N_592 => 
        N_592, N_595 => N_595, N_594 => N_594, N_586 => N_586, 
        N_582 => N_582, N_578 => N_578, N_574 => N_574, N_571 => 
        N_571, N_570 => N_570, N_569 => N_569, N_96 => N_96, N_81
         => N_81, N_74 => N_74, N_75 => N_75, N_499 => N_499, 
        N_501 => N_501, N_525 => N_525, N_513 => N_513, N_502 => 
        N_502, N_522 => N_522, N_500 => N_500, N_514 => N_514, 
        N_515 => N_515, N_524 => N_524, N_526 => N_526, N_529 => 
        N_529, N_528 => N_528, N_523 => N_523, N_517 => N_517, 
        N_505 => N_505, N_503 => N_503, N_512 => N_512, N_508 => 
        N_508, N_504 => N_504, N_520 => N_520, N_516 => N_516, 
        ren_pos => \ren_pos\, N_228 => N_228, N_7 => N_7, N_566
         => N_566, N_567 => N_567, N_565 => N_565);
    
    \reg_1x32_0\ : reg_1x32
      port map(line(31) => line_31, line(30) => \line_1[30]\, 
        line(29) => \line_5[29]\, line(28) => line_28, line(27)
         => \line_1[27]\, line(26) => \line_5[26]\, line(25) => 
        \line_1[25]\, line(24) => \line_5[24]\, line(23) => 
        \line_1[23]\, line(22) => \line_1[22]\, line(21) => 
        \line_5[21]\, line(20) => line_20, line(19) => 
        \line_0[19]\, line(18) => \line_5[18]\, line(17) => 
        \line_5[17]\, line(16) => \line_1[16]\, line(15) => 
        \line_1[15]\, line(14) => \line_5[14]\, line(13) => 
        \line_5[13]\, line(12) => \line_1[12]\, line(11) => 
        line_11, line(10) => line_10, line(9) => \line_5[9]\, 
        line(8) => \line_0[8]\, line(7) => line_7_d0, line(6) => 
        \line_5[6]\, line(5) => \line_5[5]\, line(4) => 
        \line_5[4]\, line(3) => \line_5[3]\, line(2) => 
        \line_5[2]\, line(1) => \line_1[1]\, line(0) => 
        \line_5[0]\, SHA256_BLOCK_0_H0_o(31) => 
        SHA256_BLOCK_0_H0_o(31), SHA256_BLOCK_0_H0_o(30) => 
        SHA256_BLOCK_0_H0_o(30), SHA256_BLOCK_0_H0_o(29) => 
        SHA256_BLOCK_0_H0_o(29), SHA256_BLOCK_0_H0_o(28) => 
        SHA256_BLOCK_0_H0_o(28), SHA256_BLOCK_0_H0_o(27) => 
        SHA256_BLOCK_0_H0_o(27), SHA256_BLOCK_0_H0_o(26) => 
        SHA256_BLOCK_0_H0_o(26), SHA256_BLOCK_0_H0_o(25) => 
        SHA256_BLOCK_0_H0_o(25), SHA256_BLOCK_0_H0_o(24) => 
        SHA256_BLOCK_0_H0_o(24), SHA256_BLOCK_0_H0_o(23) => 
        SHA256_BLOCK_0_H0_o(23), SHA256_BLOCK_0_H0_o(22) => 
        SHA256_BLOCK_0_H0_o(22), SHA256_BLOCK_0_H0_o(21) => 
        SHA256_BLOCK_0_H0_o(21), SHA256_BLOCK_0_H0_o(20) => 
        SHA256_BLOCK_0_H0_o(20), SHA256_BLOCK_0_H0_o(19) => 
        SHA256_BLOCK_0_H0_o(19), SHA256_BLOCK_0_H0_o(18) => 
        SHA256_BLOCK_0_H0_o(18), SHA256_BLOCK_0_H0_o(17) => 
        SHA256_BLOCK_0_H0_o(17), SHA256_BLOCK_0_H0_o(16) => 
        SHA256_BLOCK_0_H0_o(16), SHA256_BLOCK_0_H0_o(15) => 
        SHA256_BLOCK_0_H0_o(15), SHA256_BLOCK_0_H0_o(14) => 
        SHA256_BLOCK_0_H0_o(14), SHA256_BLOCK_0_H0_o(13) => 
        SHA256_BLOCK_0_H0_o(13), SHA256_BLOCK_0_H0_o(12) => 
        SHA256_BLOCK_0_H0_o(12), SHA256_BLOCK_0_H0_o(11) => 
        SHA256_BLOCK_0_H0_o(11), SHA256_BLOCK_0_H0_o(10) => 
        SHA256_BLOCK_0_H0_o(10), SHA256_BLOCK_0_H0_o(9) => 
        SHA256_BLOCK_0_H0_o(9), SHA256_BLOCK_0_H0_o(8) => 
        SHA256_BLOCK_0_H0_o(8), SHA256_BLOCK_0_H0_o(7) => 
        SHA256_BLOCK_0_H0_o(7), SHA256_BLOCK_0_H0_o(6) => 
        SHA256_BLOCK_0_H0_o(6), SHA256_BLOCK_0_H0_o(5) => 
        SHA256_BLOCK_0_H0_o(5), SHA256_BLOCK_0_H0_o(4) => 
        SHA256_BLOCK_0_H0_o(4), SHA256_BLOCK_0_H0_o(3) => 
        SHA256_BLOCK_0_H0_o(3), SHA256_BLOCK_0_H0_o(2) => 
        SHA256_BLOCK_0_H0_o(2), SHA256_BLOCK_0_H0_o(1) => 
        SHA256_BLOCK_0_H0_o(1), SHA256_BLOCK_0_H0_o(0) => 
        SHA256_BLOCK_0_H0_o(0), sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, wen_or => wen_or, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready, ren_pos => \ren_pos\, 
        AHB_slave_dummy_0_read_en => AHB_slave_dummy_0_read_en, 
        SHA256_Module_0_do_valid_o => SHA256_Module_0_do_valid_o, 
        prev_sig => prev_sig, limiter_1cycle_0_sig_1cycle => 
        limiter_1cycle_0_sig_1cycle);
    
    \reg_1x32_7\ : reg_1x32_7
      port map(line(31) => line_6_31, line(30) => \line_4[30]\, 
        line(29) => \line_0[29]\, line(28) => line_6_28, line(27)
         => \line_4[27]\, line(26) => \line_0[26]\, line(25) => 
        \line_4[25]\, line(24) => \line_0[24]\, line(23) => 
        \line_4[23]\, line(22) => \line_3[22]\, line(21) => 
        \line_0[21]\, line(20) => line_6_20, line(19) => 
        \line_4[19]\, line(18) => \line_0[18]\, line(17) => 
        \line_0[17]\, line(16) => \line_4[16]\, line(15) => 
        \line_4[15]\, line(14) => \line_0[14]\, line(13) => 
        \line_0[13]\, line(12) => \line_3[12]\, line(11) => 
        line_6_11, line(10) => line_6_10, line(9) => \line_0[9]\, 
        line(8) => \line_4[8]\, line(7) => line_6_7, line(6) => 
        \line_0[6]\, line(5) => \line_0[5]\, line(4) => 
        \line_0[4]\, line(3) => \line_0[3]\, line(2) => 
        \line_0[2]\, line(1) => \line_4[1]\, line(0) => 
        \line_0[0]\, SHA256_BLOCK_0_H7_o(31) => 
        SHA256_BLOCK_0_H7_o(31), SHA256_BLOCK_0_H7_o(30) => 
        SHA256_BLOCK_0_H7_o(30), SHA256_BLOCK_0_H7_o(29) => 
        SHA256_BLOCK_0_H7_o(29), SHA256_BLOCK_0_H7_o(28) => 
        SHA256_BLOCK_0_H7_o(28), SHA256_BLOCK_0_H7_o(27) => 
        SHA256_BLOCK_0_H7_o(27), SHA256_BLOCK_0_H7_o(26) => 
        SHA256_BLOCK_0_H7_o(26), SHA256_BLOCK_0_H7_o(25) => 
        SHA256_BLOCK_0_H7_o(25), SHA256_BLOCK_0_H7_o(24) => 
        SHA256_BLOCK_0_H7_o(24), SHA256_BLOCK_0_H7_o(23) => 
        SHA256_BLOCK_0_H7_o(23), SHA256_BLOCK_0_H7_o(22) => 
        SHA256_BLOCK_0_H7_o(22), SHA256_BLOCK_0_H7_o(21) => 
        SHA256_BLOCK_0_H7_o(21), SHA256_BLOCK_0_H7_o(20) => 
        SHA256_BLOCK_0_H7_o(20), SHA256_BLOCK_0_H7_o(19) => 
        SHA256_BLOCK_0_H7_o(19), SHA256_BLOCK_0_H7_o(18) => 
        SHA256_BLOCK_0_H7_o(18), SHA256_BLOCK_0_H7_o(17) => 
        SHA256_BLOCK_0_H7_o(17), SHA256_BLOCK_0_H7_o(16) => 
        SHA256_BLOCK_0_H7_o(16), SHA256_BLOCK_0_H7_o(15) => 
        SHA256_BLOCK_0_H7_o(15), SHA256_BLOCK_0_H7_o(14) => 
        SHA256_BLOCK_0_H7_o(14), SHA256_BLOCK_0_H7_o(13) => 
        SHA256_BLOCK_0_H7_o(13), SHA256_BLOCK_0_H7_o(12) => 
        SHA256_BLOCK_0_H7_o(12), SHA256_BLOCK_0_H7_o(11) => 
        SHA256_BLOCK_0_H7_o(11), SHA256_BLOCK_0_H7_o(10) => 
        SHA256_BLOCK_0_H7_o(10), SHA256_BLOCK_0_H7_o(9) => 
        SHA256_BLOCK_0_H7_o(9), SHA256_BLOCK_0_H7_o(8) => 
        SHA256_BLOCK_0_H7_o(8), SHA256_BLOCK_0_H7_o(7) => 
        SHA256_BLOCK_0_H7_o(7), SHA256_BLOCK_0_H7_o(6) => 
        SHA256_BLOCK_0_H7_o(6), SHA256_BLOCK_0_H7_o(5) => 
        SHA256_BLOCK_0_H7_o(5), SHA256_BLOCK_0_H7_o(4) => 
        SHA256_BLOCK_0_H7_o(4), SHA256_BLOCK_0_H7_o(3) => 
        SHA256_BLOCK_0_H7_o(3), SHA256_BLOCK_0_H7_o(2) => 
        SHA256_BLOCK_0_H7_o(2), SHA256_BLOCK_0_H7_o(1) => 
        SHA256_BLOCK_0_H7_o(1), SHA256_BLOCK_0_H7_o(0) => 
        SHA256_BLOCK_0_H7_o(0), sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, wen_or => wen_or, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready);
    
    \reg_1x32_6\ : reg_1x32_6
      port map(line(31) => line_5_31, line(30) => \line_0[30]\, 
        line(29) => \line_4[29]\, line(28) => line_5_28, line(27)
         => \line_0[27]\, line(26) => \line_4[26]\, line(25) => 
        \line_0[25]\, line(24) => \line_4[24]\, line(23) => 
        \line_0[23]\, line(22) => \line[22]\, line(21) => 
        \line_4[21]\, line(20) => line_5_20, line(19) => 
        \line_2[19]\, line(18) => \line_4[18]\, line(17) => 
        \line_4[17]\, line(16) => \line_0[16]\, line(15) => 
        \line_0[15]\, line(14) => \line_4[14]\, line(13) => 
        \line_4[13]\, line(12) => \line[12]\, line(11) => 
        line_5_11, line(10) => line_5_10, line(9) => \line_4[9]\, 
        line(8) => \line_2[8]\, line(7) => line_5_7, line(6) => 
        \line_4[6]\, line(5) => \line_4[5]\, line(4) => 
        \line_4[4]\, line(3) => \line_4[3]\, line(2) => 
        \line_4[2]\, line(1) => \line_0[1]\, line(0) => 
        \line_4[0]\, SHA256_BLOCK_0_H6_o(31) => 
        SHA256_BLOCK_0_H6_o(31), SHA256_BLOCK_0_H6_o(30) => 
        SHA256_BLOCK_0_H6_o(30), SHA256_BLOCK_0_H6_o(29) => 
        SHA256_BLOCK_0_H6_o(29), SHA256_BLOCK_0_H6_o(28) => 
        SHA256_BLOCK_0_H6_o(28), SHA256_BLOCK_0_H6_o(27) => 
        SHA256_BLOCK_0_H6_o(27), SHA256_BLOCK_0_H6_o(26) => 
        SHA256_BLOCK_0_H6_o(26), SHA256_BLOCK_0_H6_o(25) => 
        SHA256_BLOCK_0_H6_o(25), SHA256_BLOCK_0_H6_o(24) => 
        SHA256_BLOCK_0_H6_o(24), SHA256_BLOCK_0_H6_o(23) => 
        SHA256_BLOCK_0_H6_o(23), SHA256_BLOCK_0_H6_o(22) => 
        SHA256_BLOCK_0_H6_o(22), SHA256_BLOCK_0_H6_o(21) => 
        SHA256_BLOCK_0_H6_o(21), SHA256_BLOCK_0_H6_o(20) => 
        SHA256_BLOCK_0_H6_o(20), SHA256_BLOCK_0_H6_o(19) => 
        SHA256_BLOCK_0_H6_o(19), SHA256_BLOCK_0_H6_o(18) => 
        SHA256_BLOCK_0_H6_o(18), SHA256_BLOCK_0_H6_o(17) => 
        SHA256_BLOCK_0_H6_o(17), SHA256_BLOCK_0_H6_o(16) => 
        SHA256_BLOCK_0_H6_o(16), SHA256_BLOCK_0_H6_o(15) => 
        SHA256_BLOCK_0_H6_o(15), SHA256_BLOCK_0_H6_o(14) => 
        SHA256_BLOCK_0_H6_o(14), SHA256_BLOCK_0_H6_o(13) => 
        SHA256_BLOCK_0_H6_o(13), SHA256_BLOCK_0_H6_o(12) => 
        SHA256_BLOCK_0_H6_o(12), SHA256_BLOCK_0_H6_o(11) => 
        SHA256_BLOCK_0_H6_o(11), SHA256_BLOCK_0_H6_o(10) => 
        SHA256_BLOCK_0_H6_o(10), SHA256_BLOCK_0_H6_o(9) => 
        SHA256_BLOCK_0_H6_o(9), SHA256_BLOCK_0_H6_o(8) => 
        SHA256_BLOCK_0_H6_o(8), SHA256_BLOCK_0_H6_o(7) => 
        SHA256_BLOCK_0_H6_o(7), SHA256_BLOCK_0_H6_o(6) => 
        SHA256_BLOCK_0_H6_o(6), SHA256_BLOCK_0_H6_o(5) => 
        SHA256_BLOCK_0_H6_o(5), SHA256_BLOCK_0_H6_o(4) => 
        SHA256_BLOCK_0_H6_o(4), SHA256_BLOCK_0_H6_o(3) => 
        SHA256_BLOCK_0_H6_o(3), SHA256_BLOCK_0_H6_o(2) => 
        SHA256_BLOCK_0_H6_o(2), SHA256_BLOCK_0_H6_o(1) => 
        SHA256_BLOCK_0_H6_o(1), SHA256_BLOCK_0_H6_o(0) => 
        SHA256_BLOCK_0_H6_o(0), sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, wen_or => wen_or, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \reg_1x32_5\ : reg_1x32_5
      port map(line(31) => line_4_31, line(30) => \line_6[30]\, 
        line(29) => \line_2[29]\, line(28) => line_4_28, line(27)
         => \line_6[27]\, line(26) => \line_2[26]\, line(25) => 
        \line_6[25]\, line(24) => \line_2[24]\, line(23) => 
        \line_6[23]\, line(22) => \line_6[22]\, line(21) => 
        \line_2[21]\, line(20) => line_4_20, line(19) => 
        \line_6[19]\, line(18) => \line_2[18]\, line(17) => 
        \line_2[17]\, line(16) => \line_6[16]\, line(15) => 
        \line_6[15]\, line(14) => \line_2[14]\, line(13) => 
        \line_2[13]\, line(12) => \line_6[12]\, line(11) => 
        line_4_11, line(10) => line_4_10, line(9) => \line_2[9]\, 
        line(8) => \line_6[8]\, line(7) => line_4_7, line(6) => 
        \line_2[6]\, line(5) => \line_2[5]\, line(4) => 
        \line_2[4]\, line(3) => \line_2[3]\, line(2) => 
        \line_2[2]\, line(1) => \line_6[1]\, line(0) => 
        \line_2[0]\, SHA256_BLOCK_0_H5_o(31) => 
        SHA256_BLOCK_0_H5_o(31), SHA256_BLOCK_0_H5_o(30) => 
        SHA256_BLOCK_0_H5_o(30), SHA256_BLOCK_0_H5_o(29) => 
        SHA256_BLOCK_0_H5_o(29), SHA256_BLOCK_0_H5_o(28) => 
        SHA256_BLOCK_0_H5_o(28), SHA256_BLOCK_0_H5_o(27) => 
        SHA256_BLOCK_0_H5_o(27), SHA256_BLOCK_0_H5_o(26) => 
        SHA256_BLOCK_0_H5_o(26), SHA256_BLOCK_0_H5_o(25) => 
        SHA256_BLOCK_0_H5_o(25), SHA256_BLOCK_0_H5_o(24) => 
        SHA256_BLOCK_0_H5_o(24), SHA256_BLOCK_0_H5_o(23) => 
        SHA256_BLOCK_0_H5_o(23), SHA256_BLOCK_0_H5_o(22) => 
        SHA256_BLOCK_0_H5_o(22), SHA256_BLOCK_0_H5_o(21) => 
        SHA256_BLOCK_0_H5_o(21), SHA256_BLOCK_0_H5_o(20) => 
        SHA256_BLOCK_0_H5_o(20), SHA256_BLOCK_0_H5_o(19) => 
        SHA256_BLOCK_0_H5_o(19), SHA256_BLOCK_0_H5_o(18) => 
        SHA256_BLOCK_0_H5_o(18), SHA256_BLOCK_0_H5_o(17) => 
        SHA256_BLOCK_0_H5_o(17), SHA256_BLOCK_0_H5_o(16) => 
        SHA256_BLOCK_0_H5_o(16), SHA256_BLOCK_0_H5_o(15) => 
        SHA256_BLOCK_0_H5_o(15), SHA256_BLOCK_0_H5_o(14) => 
        SHA256_BLOCK_0_H5_o(14), SHA256_BLOCK_0_H5_o(13) => 
        SHA256_BLOCK_0_H5_o(13), SHA256_BLOCK_0_H5_o(12) => 
        SHA256_BLOCK_0_H5_o(12), SHA256_BLOCK_0_H5_o(11) => 
        SHA256_BLOCK_0_H5_o(11), SHA256_BLOCK_0_H5_o(10) => 
        SHA256_BLOCK_0_H5_o(10), SHA256_BLOCK_0_H5_o(9) => 
        SHA256_BLOCK_0_H5_o(9), SHA256_BLOCK_0_H5_o(8) => 
        SHA256_BLOCK_0_H5_o(8), SHA256_BLOCK_0_H5_o(7) => 
        SHA256_BLOCK_0_H5_o(7), SHA256_BLOCK_0_H5_o(6) => 
        SHA256_BLOCK_0_H5_o(6), SHA256_BLOCK_0_H5_o(5) => 
        SHA256_BLOCK_0_H5_o(5), SHA256_BLOCK_0_H5_o(4) => 
        SHA256_BLOCK_0_H5_o(4), SHA256_BLOCK_0_H5_o(3) => 
        SHA256_BLOCK_0_H5_o(3), SHA256_BLOCK_0_H5_o(2) => 
        SHA256_BLOCK_0_H5_o(2), SHA256_BLOCK_0_H5_o(1) => 
        SHA256_BLOCK_0_H5_o(1), SHA256_BLOCK_0_H5_o(0) => 
        SHA256_BLOCK_0_H5_o(0), sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, wen_or => wen_or, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready);
    
    \reg_1x32_2\ : reg_1x32_2
      port map(line(31) => line_1_31, line(30) => \line[30]\, 
        line(29) => \line_3[29]\, line(28) => line_1_28, line(27)
         => \line[27]\, line(26) => \line_3[26]\, line(25) => 
        \line[25]\, line(24) => \line_3[24]\, line(23) => 
        \line[23]\, line(22) => \line_0[22]\, line(21) => 
        \line_3[21]\, line(20) => line_1_20, line(19) => 
        \line_1[19]\, line(18) => \line_3[18]\, line(17) => 
        \line_3[17]\, line(16) => \line[16]\, line(15) => 
        \line[15]\, line(14) => \line_3[14]\, line(13) => 
        \line_3[13]\, line(12) => \line_0[12]\, line(11) => 
        line_1_11, line(10) => line_1_10, line(9) => \line_3[9]\, 
        line(8) => \line_1[8]\, line(7) => line_1_7, line(6) => 
        \line_3[6]\, line(5) => \line_3[5]\, line(4) => 
        \line_3[4]\, line(3) => \line_3[3]\, line(2) => 
        \line_3[2]\, line(1) => \line[1]\, line(0) => \line_3[0]\, 
        SHA256_BLOCK_0_H2_o(31) => SHA256_BLOCK_0_H2_o(31), 
        SHA256_BLOCK_0_H2_o(30) => SHA256_BLOCK_0_H2_o(30), 
        SHA256_BLOCK_0_H2_o(29) => SHA256_BLOCK_0_H2_o(29), 
        SHA256_BLOCK_0_H2_o(28) => SHA256_BLOCK_0_H2_o(28), 
        SHA256_BLOCK_0_H2_o(27) => SHA256_BLOCK_0_H2_o(27), 
        SHA256_BLOCK_0_H2_o(26) => SHA256_BLOCK_0_H2_o(26), 
        SHA256_BLOCK_0_H2_o(25) => SHA256_BLOCK_0_H2_o(25), 
        SHA256_BLOCK_0_H2_o(24) => SHA256_BLOCK_0_H2_o(24), 
        SHA256_BLOCK_0_H2_o(23) => SHA256_BLOCK_0_H2_o(23), 
        SHA256_BLOCK_0_H2_o(22) => SHA256_BLOCK_0_H2_o(22), 
        SHA256_BLOCK_0_H2_o(21) => SHA256_BLOCK_0_H2_o(21), 
        SHA256_BLOCK_0_H2_o(20) => SHA256_BLOCK_0_H2_o(20), 
        SHA256_BLOCK_0_H2_o(19) => SHA256_BLOCK_0_H2_o(19), 
        SHA256_BLOCK_0_H2_o(18) => SHA256_BLOCK_0_H2_o(18), 
        SHA256_BLOCK_0_H2_o(17) => SHA256_BLOCK_0_H2_o(17), 
        SHA256_BLOCK_0_H2_o(16) => SHA256_BLOCK_0_H2_o(16), 
        SHA256_BLOCK_0_H2_o(15) => SHA256_BLOCK_0_H2_o(15), 
        SHA256_BLOCK_0_H2_o(14) => SHA256_BLOCK_0_H2_o(14), 
        SHA256_BLOCK_0_H2_o(13) => SHA256_BLOCK_0_H2_o(13), 
        SHA256_BLOCK_0_H2_o(12) => SHA256_BLOCK_0_H2_o(12), 
        SHA256_BLOCK_0_H2_o(11) => SHA256_BLOCK_0_H2_o(11), 
        SHA256_BLOCK_0_H2_o(10) => SHA256_BLOCK_0_H2_o(10), 
        SHA256_BLOCK_0_H2_o(9) => SHA256_BLOCK_0_H2_o(9), 
        SHA256_BLOCK_0_H2_o(8) => SHA256_BLOCK_0_H2_o(8), 
        SHA256_BLOCK_0_H2_o(7) => SHA256_BLOCK_0_H2_o(7), 
        SHA256_BLOCK_0_H2_o(6) => SHA256_BLOCK_0_H2_o(6), 
        SHA256_BLOCK_0_H2_o(5) => SHA256_BLOCK_0_H2_o(5), 
        SHA256_BLOCK_0_H2_o(4) => SHA256_BLOCK_0_H2_o(4), 
        SHA256_BLOCK_0_H2_o(3) => SHA256_BLOCK_0_H2_o(3), 
        SHA256_BLOCK_0_H2_o(2) => SHA256_BLOCK_0_H2_o(2), 
        SHA256_BLOCK_0_H2_o(1) => SHA256_BLOCK_0_H2_o(1), 
        SHA256_BLOCK_0_H2_o(0) => SHA256_BLOCK_0_H2_o(0), 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, wen_or => wen_or, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready);
    
    reg_1x32_8 : reg_1x32_0
      port map(line_2 => \line_7[2]\, line_1 => \line_7[1]\, 
        line_0 => \line_7[0]\, line_28 => line_7_28, line_20 => 
        line_7_20, line_19 => \line_7[19]\, line_11 => line_7_11, 
        line_10 => line_7_10, line_8 => \line_7[8]\, line_7 => 
        line_7_7, sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, SHA256_Module_0_error_o => 
        SHA256_Module_0_error_o, wen_or => wen_or, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready, SHA256_Module_0_di_req_o
         => SHA256_Module_0_di_req_o, SHA256_Module_0_do_valid_o
         => SHA256_Module_0_do_valid_o, 
        SHA256_Module_0_data_available_lastbank_8 => 
        SHA256_Module_0_data_available_lastbank_8, 
        limiter_1cycle_0_sig_1cycle => 
        limiter_1cycle_0_sig_1cycle);
    
    \reg_1x32_3\ : reg_1x32_3
      port map(line(31) => line_2_31, line(30) => \line_3[30]\, 
        line(29) => \line[29]\, line(28) => line_2_28, line(27)
         => \line_3[27]\, line(26) => \line[26]\, line(25) => 
        \line_3[25]\, line(24) => \line[24]\, line(23) => 
        \line_3[23]\, line(22) => \line_4[22]\, line(21) => 
        \line[21]\, line(20) => line_2_20, line(19) => 
        \line_3[19]\, line(18) => \line[18]\, line(17) => 
        \line[17]\, line(16) => \line_3[16]\, line(15) => 
        \line_3[15]\, line(14) => \line[14]\, line(13) => 
        \line[13]\, line(12) => \line_4[12]\, line(11) => 
        line_2_11, line(10) => line_2_10, line(9) => \line[9]\, 
        line(8) => \line_3[8]\, line(7) => line_2_7, line(6) => 
        \line[6]\, line(5) => \line[5]\, line(4) => \line[4]\, 
        line(3) => \line[3]\, line(2) => \line[2]\, line(1) => 
        \line_3[1]\, line(0) => \line[0]\, 
        SHA256_BLOCK_0_H3_o(31) => SHA256_BLOCK_0_H3_o(31), 
        SHA256_BLOCK_0_H3_o(30) => SHA256_BLOCK_0_H3_o(30), 
        SHA256_BLOCK_0_H3_o(29) => SHA256_BLOCK_0_H3_o(29), 
        SHA256_BLOCK_0_H3_o(28) => SHA256_BLOCK_0_H3_o(28), 
        SHA256_BLOCK_0_H3_o(27) => SHA256_BLOCK_0_H3_o(27), 
        SHA256_BLOCK_0_H3_o(26) => SHA256_BLOCK_0_H3_o(26), 
        SHA256_BLOCK_0_H3_o(25) => SHA256_BLOCK_0_H3_o(25), 
        SHA256_BLOCK_0_H3_o(24) => SHA256_BLOCK_0_H3_o(24), 
        SHA256_BLOCK_0_H3_o(23) => SHA256_BLOCK_0_H3_o(23), 
        SHA256_BLOCK_0_H3_o(22) => SHA256_BLOCK_0_H3_o(22), 
        SHA256_BLOCK_0_H3_o(21) => SHA256_BLOCK_0_H3_o(21), 
        SHA256_BLOCK_0_H3_o(20) => SHA256_BLOCK_0_H3_o(20), 
        SHA256_BLOCK_0_H3_o(19) => SHA256_BLOCK_0_H3_o(19), 
        SHA256_BLOCK_0_H3_o(18) => SHA256_BLOCK_0_H3_o(18), 
        SHA256_BLOCK_0_H3_o(17) => SHA256_BLOCK_0_H3_o(17), 
        SHA256_BLOCK_0_H3_o(16) => SHA256_BLOCK_0_H3_o(16), 
        SHA256_BLOCK_0_H3_o(15) => SHA256_BLOCK_0_H3_o(15), 
        SHA256_BLOCK_0_H3_o(14) => SHA256_BLOCK_0_H3_o(14), 
        SHA256_BLOCK_0_H3_o(13) => SHA256_BLOCK_0_H3_o(13), 
        SHA256_BLOCK_0_H3_o(12) => SHA256_BLOCK_0_H3_o(12), 
        SHA256_BLOCK_0_H3_o(11) => SHA256_BLOCK_0_H3_o(11), 
        SHA256_BLOCK_0_H3_o(10) => SHA256_BLOCK_0_H3_o(10), 
        SHA256_BLOCK_0_H3_o(9) => SHA256_BLOCK_0_H3_o(9), 
        SHA256_BLOCK_0_H3_o(8) => SHA256_BLOCK_0_H3_o(8), 
        SHA256_BLOCK_0_H3_o(7) => SHA256_BLOCK_0_H3_o(7), 
        SHA256_BLOCK_0_H3_o(6) => SHA256_BLOCK_0_H3_o(6), 
        SHA256_BLOCK_0_H3_o(5) => SHA256_BLOCK_0_H3_o(5), 
        SHA256_BLOCK_0_H3_o(4) => SHA256_BLOCK_0_H3_o(4), 
        SHA256_BLOCK_0_H3_o(3) => SHA256_BLOCK_0_H3_o(3), 
        SHA256_BLOCK_0_H3_o(2) => SHA256_BLOCK_0_H3_o(2), 
        SHA256_BLOCK_0_H3_o(1) => SHA256_BLOCK_0_H3_o(1), 
        SHA256_BLOCK_0_H3_o(0) => SHA256_BLOCK_0_H3_o(0), 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, wen_or => wen_or, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready);
    
    \reg_1x32_4\ : reg_1x32_4
      port map(line(31) => line_3_31, line(30) => \line_2[30]\, 
        line(29) => \line_6[29]\, line(28) => line_3_28, line(27)
         => \line_2[27]\, line(26) => \line_6[26]\, line(25) => 
        \line_2[25]\, line(24) => \line_6[24]\, line(23) => 
        \line_2[23]\, line(22) => \line_2[22]\, line(21) => 
        \line_6[21]\, line(20) => line_3_20, line(19) => 
        \line[19]\, line(18) => \line_6[18]\, line(17) => 
        \line_6[17]\, line(16) => \line_2[16]\, line(15) => 
        \line_2[15]\, line(14) => \line_6[14]\, line(13) => 
        \line_6[13]\, line(12) => \line_2[12]\, line(11) => 
        line_3_11, line(10) => line_3_10, line(9) => \line_6[9]\, 
        line(8) => \line[8]\, line(7) => line_3_7, line(6) => 
        \line_6[6]\, line(5) => \line_6[5]\, line(4) => 
        \line_6[4]\, line(3) => \line_6[3]\, line(2) => 
        \line_6[2]\, line(1) => \line_2[1]\, line(0) => 
        \line_6[0]\, SHA256_BLOCK_0_H4_o(31) => 
        SHA256_BLOCK_0_H4_o(31), SHA256_BLOCK_0_H4_o(30) => 
        SHA256_BLOCK_0_H4_o(30), SHA256_BLOCK_0_H4_o(29) => 
        SHA256_BLOCK_0_H4_o(29), SHA256_BLOCK_0_H4_o(28) => 
        SHA256_BLOCK_0_H4_o(28), SHA256_BLOCK_0_H4_o(27) => 
        SHA256_BLOCK_0_H4_o(27), SHA256_BLOCK_0_H4_o(26) => 
        SHA256_BLOCK_0_H4_o(26), SHA256_BLOCK_0_H4_o(25) => 
        SHA256_BLOCK_0_H4_o(25), SHA256_BLOCK_0_H4_o(24) => 
        SHA256_BLOCK_0_H4_o(24), SHA256_BLOCK_0_H4_o(23) => 
        SHA256_BLOCK_0_H4_o(23), SHA256_BLOCK_0_H4_o(22) => 
        SHA256_BLOCK_0_H4_o(22), SHA256_BLOCK_0_H4_o(21) => 
        SHA256_BLOCK_0_H4_o(21), SHA256_BLOCK_0_H4_o(20) => 
        SHA256_BLOCK_0_H4_o(20), SHA256_BLOCK_0_H4_o(19) => 
        SHA256_BLOCK_0_H4_o(19), SHA256_BLOCK_0_H4_o(18) => 
        SHA256_BLOCK_0_H4_o(18), SHA256_BLOCK_0_H4_o(17) => 
        SHA256_BLOCK_0_H4_o(17), SHA256_BLOCK_0_H4_o(16) => 
        SHA256_BLOCK_0_H4_o(16), SHA256_BLOCK_0_H4_o(15) => 
        SHA256_BLOCK_0_H4_o(15), SHA256_BLOCK_0_H4_o(14) => 
        SHA256_BLOCK_0_H4_o(14), SHA256_BLOCK_0_H4_o(13) => 
        SHA256_BLOCK_0_H4_o(13), SHA256_BLOCK_0_H4_o(12) => 
        SHA256_BLOCK_0_H4_o(12), SHA256_BLOCK_0_H4_o(11) => 
        SHA256_BLOCK_0_H4_o(11), SHA256_BLOCK_0_H4_o(10) => 
        SHA256_BLOCK_0_H4_o(10), SHA256_BLOCK_0_H4_o(9) => 
        SHA256_BLOCK_0_H4_o(9), SHA256_BLOCK_0_H4_o(8) => 
        SHA256_BLOCK_0_H4_o(8), SHA256_BLOCK_0_H4_o(7) => 
        SHA256_BLOCK_0_H4_o(7), SHA256_BLOCK_0_H4_o(6) => 
        SHA256_BLOCK_0_H4_o(6), SHA256_BLOCK_0_H4_o(5) => 
        SHA256_BLOCK_0_H4_o(5), SHA256_BLOCK_0_H4_o(4) => 
        SHA256_BLOCK_0_H4_o(4), SHA256_BLOCK_0_H4_o(3) => 
        SHA256_BLOCK_0_H4_o(3), SHA256_BLOCK_0_H4_o(2) => 
        SHA256_BLOCK_0_H4_o(2), SHA256_BLOCK_0_H4_o(1) => 
        SHA256_BLOCK_0_H4_o(1), SHA256_BLOCK_0_H4_o(0) => 
        SHA256_BLOCK_0_H4_o(0), sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, wen_or => wen_or, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity limiter_1cycle is

    port( prev_sig                     : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK : in    std_logic;
          SHA256_Module_0_do_valid_o   : in    std_logic
        );

end limiter_1cycle;

architecture DEF_ARCH of limiter_1cycle is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \prev_sig\ : SLE
      port map(D => SHA256_Module_0_do_valid_o, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => prev_sig);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity SHA256_Module is

    port( result_addr_net_0                         : in    std_logic_vector(3 downto 0);
          AHB_slave_dummy_0_mem_wdata               : in    std_logic_vector(31 downto 0);
          waddr_in_net_0                            : in    std_logic_vector(4 downto 0);
          state_out_net_0                           : out   std_logic_vector(0 to 0);
          line_0_d0                                 : out   std_logic;
          line_3_d0                                 : out   std_logic;
          line_4_d0                                 : out   std_logic;
          line_13                                   : out   std_logic;
          line_21                                   : out   std_logic;
          line_24                                   : out   std_logic;
          line_0_0                                  : out   std_logic;
          line_0_3                                  : out   std_logic;
          line_0_4                                  : out   std_logic;
          line_0_13                                 : out   std_logic;
          line_0_21                                 : out   std_logic;
          line_0_24                                 : out   std_logic;
          line_1_0                                  : out   std_logic;
          line_1_3                                  : out   std_logic;
          line_1_4                                  : out   std_logic;
          line_1_13                                 : out   std_logic;
          line_1_21                                 : out   std_logic;
          line_1_24                                 : out   std_logic;
          line_2_0                                  : out   std_logic;
          line_2_3                                  : out   std_logic;
          line_2_4                                  : out   std_logic;
          line_2_13                                 : out   std_logic;
          line_2_21                                 : out   std_logic;
          line_2_24                                 : out   std_logic;
          line_3_0                                  : out   std_logic;
          line_3_3                                  : out   std_logic;
          line_3_4                                  : out   std_logic;
          line_3_13                                 : out   std_logic;
          line_3_21                                 : out   std_logic;
          line_3_24                                 : out   std_logic;
          line_4_0                                  : out   std_logic;
          line_4_3                                  : out   std_logic;
          line_4_4                                  : out   std_logic;
          line_4_13                                 : out   std_logic;
          line_4_21                                 : out   std_logic;
          line_4_24                                 : out   std_logic;
          line_5_0                                  : out   std_logic;
          line_5_3                                  : out   std_logic;
          line_5_4                                  : out   std_logic;
          line_5_13                                 : out   std_logic;
          line_5_21                                 : out   std_logic;
          line_5_24                                 : out   std_logic;
          line_6_0                                  : out   std_logic;
          line_6_3                                  : out   std_logic;
          line_6_4                                  : out   std_logic;
          line_6_13                                 : out   std_logic;
          line_6_21                                 : out   std_logic;
          line_6_24                                 : out   std_logic;
          line_7_21                                 : out   std_logic;
          line_7_13                                 : out   std_logic;
          line_7_4                                  : out   std_logic;
          line_7_3                                  : out   std_logic;
          line_7_0                                  : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK              : in    std_logic;
          SHA256_Module_0_do_valid_o                : out   std_logic;
          N_568                                     : out   std_logic;
          N_579                                     : out   std_logic;
          N_580                                     : out   std_logic;
          N_581                                     : out   std_logic;
          N_583                                     : out   std_logic;
          N_588                                     : out   std_logic;
          N_589                                     : out   std_logic;
          N_590                                     : out   std_logic;
          N_591                                     : out   std_logic;
          N_592                                     : out   std_logic;
          N_595                                     : out   std_logic;
          N_594                                     : out   std_logic;
          N_586                                     : out   std_logic;
          N_582                                     : out   std_logic;
          N_578                                     : out   std_logic;
          N_574                                     : out   std_logic;
          N_571                                     : out   std_logic;
          N_570                                     : out   std_logic;
          N_569                                     : out   std_logic;
          N_96                                      : out   std_logic;
          N_81                                      : out   std_logic;
          N_74                                      : out   std_logic;
          N_75                                      : out   std_logic;
          N_499                                     : out   std_logic;
          N_501                                     : out   std_logic;
          N_525                                     : out   std_logic;
          N_513                                     : out   std_logic;
          N_502                                     : out   std_logic;
          N_522                                     : out   std_logic;
          N_500                                     : out   std_logic;
          N_514                                     : out   std_logic;
          N_515                                     : out   std_logic;
          N_524                                     : out   std_logic;
          N_526                                     : out   std_logic;
          N_529                                     : out   std_logic;
          N_528                                     : out   std_logic;
          N_523                                     : out   std_logic;
          N_517                                     : out   std_logic;
          N_505                                     : out   std_logic;
          N_503                                     : out   std_logic;
          N_512                                     : out   std_logic;
          N_508                                     : out   std_logic;
          N_504                                     : out   std_logic;
          N_520                                     : out   std_logic;
          N_516                                     : out   std_logic;
          ren_pos                                   : out   std_logic;
          N_228                                     : out   std_logic;
          N_7                                       : out   std_logic;
          N_566                                     : out   std_logic;
          N_567                                     : out   std_logic;
          N_565                                     : out   std_logic;
          SHA256_Module_0_data_out_ready            : out   std_logic;
          AHB_slave_dummy_0_read_en                 : in    std_logic;
          SHA256_Module_0_error_o                   : out   std_logic;
          SHA256_Module_0_di_req_o                  : out   std_logic;
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic;
          sha256_system_sb_0_GPIO_9_M2F             : in    std_logic;
          SHA256_Module_0_data_available            : out   std_logic;
          sha256_system_sb_0_GPIO_1_M2F             : in    std_logic;
          AHB_slave_dummy_0_write_en                : in    std_logic;
          ce_i_i_2_i_0                              : out   std_logic;
          N_88_i_0                                  : out   std_logic;
          N_87_i_0                                  : out   std_logic
        );

end SHA256_Module;

architecture DEF_ARCH of SHA256_Module is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SHA256_BLOCK
    port( SHA256_BLOCK_0_H0_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o            : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o            : out   std_logic_vector(31 downto 0);
          AHB_slave_dummy_0_mem_wdata    : in    std_logic_vector(31 downto 0) := (others => 'U');
          waddr_in_net_0                 : in    std_logic_vector(4 downto 0) := (others => 'U');
          state_out_net_0                : out   std_logic_vector(0 to 0);
          sha256_system_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          SHA256_Module_0_di_req_o       : out   std_logic;
          SHA256_Module_0_do_valid_o     : out   std_logic;
          SHA256_Module_0_error_o        : out   std_logic;
          SHA256_Module_0_data_out_ready : out   std_logic;
          sha256_system_sb_0_GPIO_9_M2F  : in    std_logic := 'U';
          SHA256_Module_0_data_available : out   std_logic;
          sha256_system_sb_0_GPIO_1_M2F  : in    std_logic := 'U';
          AHB_slave_dummy_0_write_en     : in    std_logic := 'U';
          ce_i_i_2_i_0                   : out   std_logic;
          N_88_i_0                       : out   std_logic;
          N_87_i_0                       : out   std_logic
        );
  end component;

  component reg9_1x32
    port( result_addr_net_0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H0_o                       : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H1_o                       : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H2_o                       : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H3_o                       : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H4_o                       : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H5_o                       : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H6_o                       : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H7_o                       : in    std_logic_vector(31 downto 0) := (others => 'U');
          line_7_d0                                 : out   std_logic;
          line_10                                   : out   std_logic;
          line_11                                   : out   std_logic;
          line_20                                   : out   std_logic;
          line_28                                   : out   std_logic;
          line_31                                   : out   std_logic;
          line_0_7                                  : out   std_logic;
          line_0_10                                 : out   std_logic;
          line_0_11                                 : out   std_logic;
          line_0_20                                 : out   std_logic;
          line_0_28                                 : out   std_logic;
          line_0_31                                 : out   std_logic;
          line_1_7                                  : out   std_logic;
          line_1_10                                 : out   std_logic;
          line_1_11                                 : out   std_logic;
          line_1_20                                 : out   std_logic;
          line_1_28                                 : out   std_logic;
          line_1_31                                 : out   std_logic;
          line_2_7                                  : out   std_logic;
          line_2_10                                 : out   std_logic;
          line_2_11                                 : out   std_logic;
          line_2_20                                 : out   std_logic;
          line_2_28                                 : out   std_logic;
          line_2_31                                 : out   std_logic;
          line_3_7                                  : out   std_logic;
          line_3_10                                 : out   std_logic;
          line_3_11                                 : out   std_logic;
          line_3_20                                 : out   std_logic;
          line_3_28                                 : out   std_logic;
          line_3_31                                 : out   std_logic;
          line_4_7                                  : out   std_logic;
          line_4_10                                 : out   std_logic;
          line_4_11                                 : out   std_logic;
          line_4_20                                 : out   std_logic;
          line_4_28                                 : out   std_logic;
          line_4_31                                 : out   std_logic;
          line_5_7                                  : out   std_logic;
          line_5_10                                 : out   std_logic;
          line_5_11                                 : out   std_logic;
          line_5_20                                 : out   std_logic;
          line_5_28                                 : out   std_logic;
          line_5_31                                 : out   std_logic;
          line_6_7                                  : out   std_logic;
          line_6_10                                 : out   std_logic;
          line_6_11                                 : out   std_logic;
          line_6_20                                 : out   std_logic;
          line_6_28                                 : out   std_logic;
          line_6_31                                 : out   std_logic;
          line_7_28                                 : out   std_logic;
          line_7_20                                 : out   std_logic;
          line_7_11                                 : out   std_logic;
          line_7_10                                 : out   std_logic;
          line_7_7                                  : out   std_logic;
          N_568                                     : out   std_logic;
          N_579                                     : out   std_logic;
          N_580                                     : out   std_logic;
          N_581                                     : out   std_logic;
          N_583                                     : out   std_logic;
          N_588                                     : out   std_logic;
          N_589                                     : out   std_logic;
          N_590                                     : out   std_logic;
          N_591                                     : out   std_logic;
          N_592                                     : out   std_logic;
          N_595                                     : out   std_logic;
          N_594                                     : out   std_logic;
          N_586                                     : out   std_logic;
          N_582                                     : out   std_logic;
          N_578                                     : out   std_logic;
          N_574                                     : out   std_logic;
          N_571                                     : out   std_logic;
          N_570                                     : out   std_logic;
          N_569                                     : out   std_logic;
          N_96                                      : out   std_logic;
          N_81                                      : out   std_logic;
          N_74                                      : out   std_logic;
          N_75                                      : out   std_logic;
          N_499                                     : out   std_logic;
          N_501                                     : out   std_logic;
          N_525                                     : out   std_logic;
          N_513                                     : out   std_logic;
          N_502                                     : out   std_logic;
          N_522                                     : out   std_logic;
          N_500                                     : out   std_logic;
          N_514                                     : out   std_logic;
          N_515                                     : out   std_logic;
          N_524                                     : out   std_logic;
          N_526                                     : out   std_logic;
          N_529                                     : out   std_logic;
          N_528                                     : out   std_logic;
          N_523                                     : out   std_logic;
          N_517                                     : out   std_logic;
          N_505                                     : out   std_logic;
          N_503                                     : out   std_logic;
          N_512                                     : out   std_logic;
          N_508                                     : out   std_logic;
          N_504                                     : out   std_logic;
          N_520                                     : out   std_logic;
          N_516                                     : out   std_logic;
          ren_pos                                   : out   std_logic;
          N_228                                     : out   std_logic;
          N_7                                       : out   std_logic;
          N_566                                     : out   std_logic;
          N_567                                     : out   std_logic;
          N_565                                     : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK              : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready            : in    std_logic := 'U';
          AHB_slave_dummy_0_read_en                 : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o                : in    std_logic := 'U';
          prev_sig                                  : in    std_logic := 'U';
          SHA256_Module_0_error_o                   : in    std_logic := 'U';
          SHA256_Module_0_di_req_o                  : in    std_logic := 'U';
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic
        );
  end component;

  component limiter_1cycle
    port( prev_sig                     : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o   : in    std_logic := 'U'
        );
  end component;

    signal prev_sig, \SHA256_Module_0_do_valid_o\, 
        \SHA256_BLOCK_0_H0_o[0]\, \SHA256_BLOCK_0_H0_o[1]\, 
        \SHA256_BLOCK_0_H0_o[2]\, \SHA256_BLOCK_0_H0_o[3]\, 
        \SHA256_BLOCK_0_H0_o[4]\, \SHA256_BLOCK_0_H0_o[5]\, 
        \SHA256_BLOCK_0_H0_o[6]\, \SHA256_BLOCK_0_H0_o[7]\, 
        \SHA256_BLOCK_0_H0_o[8]\, \SHA256_BLOCK_0_H0_o[9]\, 
        \SHA256_BLOCK_0_H0_o[10]\, \SHA256_BLOCK_0_H0_o[11]\, 
        \SHA256_BLOCK_0_H0_o[12]\, \SHA256_BLOCK_0_H0_o[13]\, 
        \SHA256_BLOCK_0_H0_o[14]\, \SHA256_BLOCK_0_H0_o[15]\, 
        \SHA256_BLOCK_0_H0_o[16]\, \SHA256_BLOCK_0_H0_o[17]\, 
        \SHA256_BLOCK_0_H0_o[18]\, \SHA256_BLOCK_0_H0_o[19]\, 
        \SHA256_BLOCK_0_H0_o[20]\, \SHA256_BLOCK_0_H0_o[21]\, 
        \SHA256_BLOCK_0_H0_o[22]\, \SHA256_BLOCK_0_H0_o[23]\, 
        \SHA256_BLOCK_0_H0_o[24]\, \SHA256_BLOCK_0_H0_o[25]\, 
        \SHA256_BLOCK_0_H0_o[26]\, \SHA256_BLOCK_0_H0_o[27]\, 
        \SHA256_BLOCK_0_H0_o[28]\, \SHA256_BLOCK_0_H0_o[29]\, 
        \SHA256_BLOCK_0_H0_o[30]\, \SHA256_BLOCK_0_H0_o[31]\, 
        \SHA256_BLOCK_0_H1_o[0]\, \SHA256_BLOCK_0_H1_o[1]\, 
        \SHA256_BLOCK_0_H1_o[2]\, \SHA256_BLOCK_0_H1_o[3]\, 
        \SHA256_BLOCK_0_H1_o[4]\, \SHA256_BLOCK_0_H1_o[5]\, 
        \SHA256_BLOCK_0_H1_o[6]\, \SHA256_BLOCK_0_H1_o[7]\, 
        \SHA256_BLOCK_0_H1_o[8]\, \SHA256_BLOCK_0_H1_o[9]\, 
        \SHA256_BLOCK_0_H1_o[10]\, \SHA256_BLOCK_0_H1_o[11]\, 
        \SHA256_BLOCK_0_H1_o[12]\, \SHA256_BLOCK_0_H1_o[13]\, 
        \SHA256_BLOCK_0_H1_o[14]\, \SHA256_BLOCK_0_H1_o[15]\, 
        \SHA256_BLOCK_0_H1_o[16]\, \SHA256_BLOCK_0_H1_o[17]\, 
        \SHA256_BLOCK_0_H1_o[18]\, \SHA256_BLOCK_0_H1_o[19]\, 
        \SHA256_BLOCK_0_H1_o[20]\, \SHA256_BLOCK_0_H1_o[21]\, 
        \SHA256_BLOCK_0_H1_o[22]\, \SHA256_BLOCK_0_H1_o[23]\, 
        \SHA256_BLOCK_0_H1_o[24]\, \SHA256_BLOCK_0_H1_o[25]\, 
        \SHA256_BLOCK_0_H1_o[26]\, \SHA256_BLOCK_0_H1_o[27]\, 
        \SHA256_BLOCK_0_H1_o[28]\, \SHA256_BLOCK_0_H1_o[29]\, 
        \SHA256_BLOCK_0_H1_o[30]\, \SHA256_BLOCK_0_H1_o[31]\, 
        \SHA256_BLOCK_0_H2_o[0]\, \SHA256_BLOCK_0_H2_o[1]\, 
        \SHA256_BLOCK_0_H2_o[2]\, \SHA256_BLOCK_0_H2_o[3]\, 
        \SHA256_BLOCK_0_H2_o[4]\, \SHA256_BLOCK_0_H2_o[5]\, 
        \SHA256_BLOCK_0_H2_o[6]\, \SHA256_BLOCK_0_H2_o[7]\, 
        \SHA256_BLOCK_0_H2_o[8]\, \SHA256_BLOCK_0_H2_o[9]\, 
        \SHA256_BLOCK_0_H2_o[10]\, \SHA256_BLOCK_0_H2_o[11]\, 
        \SHA256_BLOCK_0_H2_o[12]\, \SHA256_BLOCK_0_H2_o[13]\, 
        \SHA256_BLOCK_0_H2_o[14]\, \SHA256_BLOCK_0_H2_o[15]\, 
        \SHA256_BLOCK_0_H2_o[16]\, \SHA256_BLOCK_0_H2_o[17]\, 
        \SHA256_BLOCK_0_H2_o[18]\, \SHA256_BLOCK_0_H2_o[19]\, 
        \SHA256_BLOCK_0_H2_o[20]\, \SHA256_BLOCK_0_H2_o[21]\, 
        \SHA256_BLOCK_0_H2_o[22]\, \SHA256_BLOCK_0_H2_o[23]\, 
        \SHA256_BLOCK_0_H2_o[24]\, \SHA256_BLOCK_0_H2_o[25]\, 
        \SHA256_BLOCK_0_H2_o[26]\, \SHA256_BLOCK_0_H2_o[27]\, 
        \SHA256_BLOCK_0_H2_o[28]\, \SHA256_BLOCK_0_H2_o[29]\, 
        \SHA256_BLOCK_0_H2_o[30]\, \SHA256_BLOCK_0_H2_o[31]\, 
        \SHA256_BLOCK_0_H3_o[0]\, \SHA256_BLOCK_0_H3_o[1]\, 
        \SHA256_BLOCK_0_H3_o[2]\, \SHA256_BLOCK_0_H3_o[3]\, 
        \SHA256_BLOCK_0_H3_o[4]\, \SHA256_BLOCK_0_H3_o[5]\, 
        \SHA256_BLOCK_0_H3_o[6]\, \SHA256_BLOCK_0_H3_o[7]\, 
        \SHA256_BLOCK_0_H3_o[8]\, \SHA256_BLOCK_0_H3_o[9]\, 
        \SHA256_BLOCK_0_H3_o[10]\, \SHA256_BLOCK_0_H3_o[11]\, 
        \SHA256_BLOCK_0_H3_o[12]\, \SHA256_BLOCK_0_H3_o[13]\, 
        \SHA256_BLOCK_0_H3_o[14]\, \SHA256_BLOCK_0_H3_o[15]\, 
        \SHA256_BLOCK_0_H3_o[16]\, \SHA256_BLOCK_0_H3_o[17]\, 
        \SHA256_BLOCK_0_H3_o[18]\, \SHA256_BLOCK_0_H3_o[19]\, 
        \SHA256_BLOCK_0_H3_o[20]\, \SHA256_BLOCK_0_H3_o[21]\, 
        \SHA256_BLOCK_0_H3_o[22]\, \SHA256_BLOCK_0_H3_o[23]\, 
        \SHA256_BLOCK_0_H3_o[24]\, \SHA256_BLOCK_0_H3_o[25]\, 
        \SHA256_BLOCK_0_H3_o[26]\, \SHA256_BLOCK_0_H3_o[27]\, 
        \SHA256_BLOCK_0_H3_o[28]\, \SHA256_BLOCK_0_H3_o[29]\, 
        \SHA256_BLOCK_0_H3_o[30]\, \SHA256_BLOCK_0_H3_o[31]\, 
        \SHA256_BLOCK_0_H4_o[0]\, \SHA256_BLOCK_0_H4_o[1]\, 
        \SHA256_BLOCK_0_H4_o[2]\, \SHA256_BLOCK_0_H4_o[3]\, 
        \SHA256_BLOCK_0_H4_o[4]\, \SHA256_BLOCK_0_H4_o[5]\, 
        \SHA256_BLOCK_0_H4_o[6]\, \SHA256_BLOCK_0_H4_o[7]\, 
        \SHA256_BLOCK_0_H4_o[8]\, \SHA256_BLOCK_0_H4_o[9]\, 
        \SHA256_BLOCK_0_H4_o[10]\, \SHA256_BLOCK_0_H4_o[11]\, 
        \SHA256_BLOCK_0_H4_o[12]\, \SHA256_BLOCK_0_H4_o[13]\, 
        \SHA256_BLOCK_0_H4_o[14]\, \SHA256_BLOCK_0_H4_o[15]\, 
        \SHA256_BLOCK_0_H4_o[16]\, \SHA256_BLOCK_0_H4_o[17]\, 
        \SHA256_BLOCK_0_H4_o[18]\, \SHA256_BLOCK_0_H4_o[19]\, 
        \SHA256_BLOCK_0_H4_o[20]\, \SHA256_BLOCK_0_H4_o[21]\, 
        \SHA256_BLOCK_0_H4_o[22]\, \SHA256_BLOCK_0_H4_o[23]\, 
        \SHA256_BLOCK_0_H4_o[24]\, \SHA256_BLOCK_0_H4_o[25]\, 
        \SHA256_BLOCK_0_H4_o[26]\, \SHA256_BLOCK_0_H4_o[27]\, 
        \SHA256_BLOCK_0_H4_o[28]\, \SHA256_BLOCK_0_H4_o[29]\, 
        \SHA256_BLOCK_0_H4_o[30]\, \SHA256_BLOCK_0_H4_o[31]\, 
        \SHA256_BLOCK_0_H5_o[0]\, \SHA256_BLOCK_0_H5_o[1]\, 
        \SHA256_BLOCK_0_H5_o[2]\, \SHA256_BLOCK_0_H5_o[3]\, 
        \SHA256_BLOCK_0_H5_o[4]\, \SHA256_BLOCK_0_H5_o[5]\, 
        \SHA256_BLOCK_0_H5_o[6]\, \SHA256_BLOCK_0_H5_o[7]\, 
        \SHA256_BLOCK_0_H5_o[8]\, \SHA256_BLOCK_0_H5_o[9]\, 
        \SHA256_BLOCK_0_H5_o[10]\, \SHA256_BLOCK_0_H5_o[11]\, 
        \SHA256_BLOCK_0_H5_o[12]\, \SHA256_BLOCK_0_H5_o[13]\, 
        \SHA256_BLOCK_0_H5_o[14]\, \SHA256_BLOCK_0_H5_o[15]\, 
        \SHA256_BLOCK_0_H5_o[16]\, \SHA256_BLOCK_0_H5_o[17]\, 
        \SHA256_BLOCK_0_H5_o[18]\, \SHA256_BLOCK_0_H5_o[19]\, 
        \SHA256_BLOCK_0_H5_o[20]\, \SHA256_BLOCK_0_H5_o[21]\, 
        \SHA256_BLOCK_0_H5_o[22]\, \SHA256_BLOCK_0_H5_o[23]\, 
        \SHA256_BLOCK_0_H5_o[24]\, \SHA256_BLOCK_0_H5_o[25]\, 
        \SHA256_BLOCK_0_H5_o[26]\, \SHA256_BLOCK_0_H5_o[27]\, 
        \SHA256_BLOCK_0_H5_o[28]\, \SHA256_BLOCK_0_H5_o[29]\, 
        \SHA256_BLOCK_0_H5_o[30]\, \SHA256_BLOCK_0_H5_o[31]\, 
        \SHA256_BLOCK_0_H6_o[0]\, \SHA256_BLOCK_0_H6_o[1]\, 
        \SHA256_BLOCK_0_H6_o[2]\, \SHA256_BLOCK_0_H6_o[3]\, 
        \SHA256_BLOCK_0_H6_o[4]\, \SHA256_BLOCK_0_H6_o[5]\, 
        \SHA256_BLOCK_0_H6_o[6]\, \SHA256_BLOCK_0_H6_o[7]\, 
        \SHA256_BLOCK_0_H6_o[8]\, \SHA256_BLOCK_0_H6_o[9]\, 
        \SHA256_BLOCK_0_H6_o[10]\, \SHA256_BLOCK_0_H6_o[11]\, 
        \SHA256_BLOCK_0_H6_o[12]\, \SHA256_BLOCK_0_H6_o[13]\, 
        \SHA256_BLOCK_0_H6_o[14]\, \SHA256_BLOCK_0_H6_o[15]\, 
        \SHA256_BLOCK_0_H6_o[16]\, \SHA256_BLOCK_0_H6_o[17]\, 
        \SHA256_BLOCK_0_H6_o[18]\, \SHA256_BLOCK_0_H6_o[19]\, 
        \SHA256_BLOCK_0_H6_o[20]\, \SHA256_BLOCK_0_H6_o[21]\, 
        \SHA256_BLOCK_0_H6_o[22]\, \SHA256_BLOCK_0_H6_o[23]\, 
        \SHA256_BLOCK_0_H6_o[24]\, \SHA256_BLOCK_0_H6_o[25]\, 
        \SHA256_BLOCK_0_H6_o[26]\, \SHA256_BLOCK_0_H6_o[27]\, 
        \SHA256_BLOCK_0_H6_o[28]\, \SHA256_BLOCK_0_H6_o[29]\, 
        \SHA256_BLOCK_0_H6_o[30]\, \SHA256_BLOCK_0_H6_o[31]\, 
        \SHA256_BLOCK_0_H7_o[0]\, \SHA256_BLOCK_0_H7_o[1]\, 
        \SHA256_BLOCK_0_H7_o[2]\, \SHA256_BLOCK_0_H7_o[3]\, 
        \SHA256_BLOCK_0_H7_o[4]\, \SHA256_BLOCK_0_H7_o[5]\, 
        \SHA256_BLOCK_0_H7_o[6]\, \SHA256_BLOCK_0_H7_o[7]\, 
        \SHA256_BLOCK_0_H7_o[8]\, \SHA256_BLOCK_0_H7_o[9]\, 
        \SHA256_BLOCK_0_H7_o[10]\, \SHA256_BLOCK_0_H7_o[11]\, 
        \SHA256_BLOCK_0_H7_o[12]\, \SHA256_BLOCK_0_H7_o[13]\, 
        \SHA256_BLOCK_0_H7_o[14]\, \SHA256_BLOCK_0_H7_o[15]\, 
        \SHA256_BLOCK_0_H7_o[16]\, \SHA256_BLOCK_0_H7_o[17]\, 
        \SHA256_BLOCK_0_H7_o[18]\, \SHA256_BLOCK_0_H7_o[19]\, 
        \SHA256_BLOCK_0_H7_o[20]\, \SHA256_BLOCK_0_H7_o[21]\, 
        \SHA256_BLOCK_0_H7_o[22]\, \SHA256_BLOCK_0_H7_o[23]\, 
        \SHA256_BLOCK_0_H7_o[24]\, \SHA256_BLOCK_0_H7_o[25]\, 
        \SHA256_BLOCK_0_H7_o[26]\, \SHA256_BLOCK_0_H7_o[27]\, 
        \SHA256_BLOCK_0_H7_o[28]\, \SHA256_BLOCK_0_H7_o[29]\, 
        \SHA256_BLOCK_0_H7_o[30]\, \SHA256_BLOCK_0_H7_o[31]\, 
        \SHA256_Module_0_data_out_ready\, 
        \SHA256_Module_0_error_o\, \SHA256_Module_0_di_req_o\, 
        GND_net_1, VCC_net_1 : std_logic;

    for all : SHA256_BLOCK
	Use entity work.SHA256_BLOCK(DEF_ARCH);
    for all : reg9_1x32
	Use entity work.reg9_1x32(DEF_ARCH);
    for all : limiter_1cycle
	Use entity work.limiter_1cycle(DEF_ARCH);
begin 

    SHA256_Module_0_do_valid_o <= \SHA256_Module_0_do_valid_o\;
    SHA256_Module_0_data_out_ready <= 
        \SHA256_Module_0_data_out_ready\;
    SHA256_Module_0_error_o <= \SHA256_Module_0_error_o\;
    SHA256_Module_0_di_req_o <= \SHA256_Module_0_di_req_o\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    SHA256_BLOCK_0 : SHA256_BLOCK
      port map(SHA256_BLOCK_0_H0_o(31) => 
        \SHA256_BLOCK_0_H0_o[31]\, SHA256_BLOCK_0_H0_o(30) => 
        \SHA256_BLOCK_0_H0_o[30]\, SHA256_BLOCK_0_H0_o(29) => 
        \SHA256_BLOCK_0_H0_o[29]\, SHA256_BLOCK_0_H0_o(28) => 
        \SHA256_BLOCK_0_H0_o[28]\, SHA256_BLOCK_0_H0_o(27) => 
        \SHA256_BLOCK_0_H0_o[27]\, SHA256_BLOCK_0_H0_o(26) => 
        \SHA256_BLOCK_0_H0_o[26]\, SHA256_BLOCK_0_H0_o(25) => 
        \SHA256_BLOCK_0_H0_o[25]\, SHA256_BLOCK_0_H0_o(24) => 
        \SHA256_BLOCK_0_H0_o[24]\, SHA256_BLOCK_0_H0_o(23) => 
        \SHA256_BLOCK_0_H0_o[23]\, SHA256_BLOCK_0_H0_o(22) => 
        \SHA256_BLOCK_0_H0_o[22]\, SHA256_BLOCK_0_H0_o(21) => 
        \SHA256_BLOCK_0_H0_o[21]\, SHA256_BLOCK_0_H0_o(20) => 
        \SHA256_BLOCK_0_H0_o[20]\, SHA256_BLOCK_0_H0_o(19) => 
        \SHA256_BLOCK_0_H0_o[19]\, SHA256_BLOCK_0_H0_o(18) => 
        \SHA256_BLOCK_0_H0_o[18]\, SHA256_BLOCK_0_H0_o(17) => 
        \SHA256_BLOCK_0_H0_o[17]\, SHA256_BLOCK_0_H0_o(16) => 
        \SHA256_BLOCK_0_H0_o[16]\, SHA256_BLOCK_0_H0_o(15) => 
        \SHA256_BLOCK_0_H0_o[15]\, SHA256_BLOCK_0_H0_o(14) => 
        \SHA256_BLOCK_0_H0_o[14]\, SHA256_BLOCK_0_H0_o(13) => 
        \SHA256_BLOCK_0_H0_o[13]\, SHA256_BLOCK_0_H0_o(12) => 
        \SHA256_BLOCK_0_H0_o[12]\, SHA256_BLOCK_0_H0_o(11) => 
        \SHA256_BLOCK_0_H0_o[11]\, SHA256_BLOCK_0_H0_o(10) => 
        \SHA256_BLOCK_0_H0_o[10]\, SHA256_BLOCK_0_H0_o(9) => 
        \SHA256_BLOCK_0_H0_o[9]\, SHA256_BLOCK_0_H0_o(8) => 
        \SHA256_BLOCK_0_H0_o[8]\, SHA256_BLOCK_0_H0_o(7) => 
        \SHA256_BLOCK_0_H0_o[7]\, SHA256_BLOCK_0_H0_o(6) => 
        \SHA256_BLOCK_0_H0_o[6]\, SHA256_BLOCK_0_H0_o(5) => 
        \SHA256_BLOCK_0_H0_o[5]\, SHA256_BLOCK_0_H0_o(4) => 
        \SHA256_BLOCK_0_H0_o[4]\, SHA256_BLOCK_0_H0_o(3) => 
        \SHA256_BLOCK_0_H0_o[3]\, SHA256_BLOCK_0_H0_o(2) => 
        \SHA256_BLOCK_0_H0_o[2]\, SHA256_BLOCK_0_H0_o(1) => 
        \SHA256_BLOCK_0_H0_o[1]\, SHA256_BLOCK_0_H0_o(0) => 
        \SHA256_BLOCK_0_H0_o[0]\, SHA256_BLOCK_0_H1_o(31) => 
        \SHA256_BLOCK_0_H1_o[31]\, SHA256_BLOCK_0_H1_o(30) => 
        \SHA256_BLOCK_0_H1_o[30]\, SHA256_BLOCK_0_H1_o(29) => 
        \SHA256_BLOCK_0_H1_o[29]\, SHA256_BLOCK_0_H1_o(28) => 
        \SHA256_BLOCK_0_H1_o[28]\, SHA256_BLOCK_0_H1_o(27) => 
        \SHA256_BLOCK_0_H1_o[27]\, SHA256_BLOCK_0_H1_o(26) => 
        \SHA256_BLOCK_0_H1_o[26]\, SHA256_BLOCK_0_H1_o(25) => 
        \SHA256_BLOCK_0_H1_o[25]\, SHA256_BLOCK_0_H1_o(24) => 
        \SHA256_BLOCK_0_H1_o[24]\, SHA256_BLOCK_0_H1_o(23) => 
        \SHA256_BLOCK_0_H1_o[23]\, SHA256_BLOCK_0_H1_o(22) => 
        \SHA256_BLOCK_0_H1_o[22]\, SHA256_BLOCK_0_H1_o(21) => 
        \SHA256_BLOCK_0_H1_o[21]\, SHA256_BLOCK_0_H1_o(20) => 
        \SHA256_BLOCK_0_H1_o[20]\, SHA256_BLOCK_0_H1_o(19) => 
        \SHA256_BLOCK_0_H1_o[19]\, SHA256_BLOCK_0_H1_o(18) => 
        \SHA256_BLOCK_0_H1_o[18]\, SHA256_BLOCK_0_H1_o(17) => 
        \SHA256_BLOCK_0_H1_o[17]\, SHA256_BLOCK_0_H1_o(16) => 
        \SHA256_BLOCK_0_H1_o[16]\, SHA256_BLOCK_0_H1_o(15) => 
        \SHA256_BLOCK_0_H1_o[15]\, SHA256_BLOCK_0_H1_o(14) => 
        \SHA256_BLOCK_0_H1_o[14]\, SHA256_BLOCK_0_H1_o(13) => 
        \SHA256_BLOCK_0_H1_o[13]\, SHA256_BLOCK_0_H1_o(12) => 
        \SHA256_BLOCK_0_H1_o[12]\, SHA256_BLOCK_0_H1_o(11) => 
        \SHA256_BLOCK_0_H1_o[11]\, SHA256_BLOCK_0_H1_o(10) => 
        \SHA256_BLOCK_0_H1_o[10]\, SHA256_BLOCK_0_H1_o(9) => 
        \SHA256_BLOCK_0_H1_o[9]\, SHA256_BLOCK_0_H1_o(8) => 
        \SHA256_BLOCK_0_H1_o[8]\, SHA256_BLOCK_0_H1_o(7) => 
        \SHA256_BLOCK_0_H1_o[7]\, SHA256_BLOCK_0_H1_o(6) => 
        \SHA256_BLOCK_0_H1_o[6]\, SHA256_BLOCK_0_H1_o(5) => 
        \SHA256_BLOCK_0_H1_o[5]\, SHA256_BLOCK_0_H1_o(4) => 
        \SHA256_BLOCK_0_H1_o[4]\, SHA256_BLOCK_0_H1_o(3) => 
        \SHA256_BLOCK_0_H1_o[3]\, SHA256_BLOCK_0_H1_o(2) => 
        \SHA256_BLOCK_0_H1_o[2]\, SHA256_BLOCK_0_H1_o(1) => 
        \SHA256_BLOCK_0_H1_o[1]\, SHA256_BLOCK_0_H1_o(0) => 
        \SHA256_BLOCK_0_H1_o[0]\, SHA256_BLOCK_0_H2_o(31) => 
        \SHA256_BLOCK_0_H2_o[31]\, SHA256_BLOCK_0_H2_o(30) => 
        \SHA256_BLOCK_0_H2_o[30]\, SHA256_BLOCK_0_H2_o(29) => 
        \SHA256_BLOCK_0_H2_o[29]\, SHA256_BLOCK_0_H2_o(28) => 
        \SHA256_BLOCK_0_H2_o[28]\, SHA256_BLOCK_0_H2_o(27) => 
        \SHA256_BLOCK_0_H2_o[27]\, SHA256_BLOCK_0_H2_o(26) => 
        \SHA256_BLOCK_0_H2_o[26]\, SHA256_BLOCK_0_H2_o(25) => 
        \SHA256_BLOCK_0_H2_o[25]\, SHA256_BLOCK_0_H2_o(24) => 
        \SHA256_BLOCK_0_H2_o[24]\, SHA256_BLOCK_0_H2_o(23) => 
        \SHA256_BLOCK_0_H2_o[23]\, SHA256_BLOCK_0_H2_o(22) => 
        \SHA256_BLOCK_0_H2_o[22]\, SHA256_BLOCK_0_H2_o(21) => 
        \SHA256_BLOCK_0_H2_o[21]\, SHA256_BLOCK_0_H2_o(20) => 
        \SHA256_BLOCK_0_H2_o[20]\, SHA256_BLOCK_0_H2_o(19) => 
        \SHA256_BLOCK_0_H2_o[19]\, SHA256_BLOCK_0_H2_o(18) => 
        \SHA256_BLOCK_0_H2_o[18]\, SHA256_BLOCK_0_H2_o(17) => 
        \SHA256_BLOCK_0_H2_o[17]\, SHA256_BLOCK_0_H2_o(16) => 
        \SHA256_BLOCK_0_H2_o[16]\, SHA256_BLOCK_0_H2_o(15) => 
        \SHA256_BLOCK_0_H2_o[15]\, SHA256_BLOCK_0_H2_o(14) => 
        \SHA256_BLOCK_0_H2_o[14]\, SHA256_BLOCK_0_H2_o(13) => 
        \SHA256_BLOCK_0_H2_o[13]\, SHA256_BLOCK_0_H2_o(12) => 
        \SHA256_BLOCK_0_H2_o[12]\, SHA256_BLOCK_0_H2_o(11) => 
        \SHA256_BLOCK_0_H2_o[11]\, SHA256_BLOCK_0_H2_o(10) => 
        \SHA256_BLOCK_0_H2_o[10]\, SHA256_BLOCK_0_H2_o(9) => 
        \SHA256_BLOCK_0_H2_o[9]\, SHA256_BLOCK_0_H2_o(8) => 
        \SHA256_BLOCK_0_H2_o[8]\, SHA256_BLOCK_0_H2_o(7) => 
        \SHA256_BLOCK_0_H2_o[7]\, SHA256_BLOCK_0_H2_o(6) => 
        \SHA256_BLOCK_0_H2_o[6]\, SHA256_BLOCK_0_H2_o(5) => 
        \SHA256_BLOCK_0_H2_o[5]\, SHA256_BLOCK_0_H2_o(4) => 
        \SHA256_BLOCK_0_H2_o[4]\, SHA256_BLOCK_0_H2_o(3) => 
        \SHA256_BLOCK_0_H2_o[3]\, SHA256_BLOCK_0_H2_o(2) => 
        \SHA256_BLOCK_0_H2_o[2]\, SHA256_BLOCK_0_H2_o(1) => 
        \SHA256_BLOCK_0_H2_o[1]\, SHA256_BLOCK_0_H2_o(0) => 
        \SHA256_BLOCK_0_H2_o[0]\, SHA256_BLOCK_0_H3_o(31) => 
        \SHA256_BLOCK_0_H3_o[31]\, SHA256_BLOCK_0_H3_o(30) => 
        \SHA256_BLOCK_0_H3_o[30]\, SHA256_BLOCK_0_H3_o(29) => 
        \SHA256_BLOCK_0_H3_o[29]\, SHA256_BLOCK_0_H3_o(28) => 
        \SHA256_BLOCK_0_H3_o[28]\, SHA256_BLOCK_0_H3_o(27) => 
        \SHA256_BLOCK_0_H3_o[27]\, SHA256_BLOCK_0_H3_o(26) => 
        \SHA256_BLOCK_0_H3_o[26]\, SHA256_BLOCK_0_H3_o(25) => 
        \SHA256_BLOCK_0_H3_o[25]\, SHA256_BLOCK_0_H3_o(24) => 
        \SHA256_BLOCK_0_H3_o[24]\, SHA256_BLOCK_0_H3_o(23) => 
        \SHA256_BLOCK_0_H3_o[23]\, SHA256_BLOCK_0_H3_o(22) => 
        \SHA256_BLOCK_0_H3_o[22]\, SHA256_BLOCK_0_H3_o(21) => 
        \SHA256_BLOCK_0_H3_o[21]\, SHA256_BLOCK_0_H3_o(20) => 
        \SHA256_BLOCK_0_H3_o[20]\, SHA256_BLOCK_0_H3_o(19) => 
        \SHA256_BLOCK_0_H3_o[19]\, SHA256_BLOCK_0_H3_o(18) => 
        \SHA256_BLOCK_0_H3_o[18]\, SHA256_BLOCK_0_H3_o(17) => 
        \SHA256_BLOCK_0_H3_o[17]\, SHA256_BLOCK_0_H3_o(16) => 
        \SHA256_BLOCK_0_H3_o[16]\, SHA256_BLOCK_0_H3_o(15) => 
        \SHA256_BLOCK_0_H3_o[15]\, SHA256_BLOCK_0_H3_o(14) => 
        \SHA256_BLOCK_0_H3_o[14]\, SHA256_BLOCK_0_H3_o(13) => 
        \SHA256_BLOCK_0_H3_o[13]\, SHA256_BLOCK_0_H3_o(12) => 
        \SHA256_BLOCK_0_H3_o[12]\, SHA256_BLOCK_0_H3_o(11) => 
        \SHA256_BLOCK_0_H3_o[11]\, SHA256_BLOCK_0_H3_o(10) => 
        \SHA256_BLOCK_0_H3_o[10]\, SHA256_BLOCK_0_H3_o(9) => 
        \SHA256_BLOCK_0_H3_o[9]\, SHA256_BLOCK_0_H3_o(8) => 
        \SHA256_BLOCK_0_H3_o[8]\, SHA256_BLOCK_0_H3_o(7) => 
        \SHA256_BLOCK_0_H3_o[7]\, SHA256_BLOCK_0_H3_o(6) => 
        \SHA256_BLOCK_0_H3_o[6]\, SHA256_BLOCK_0_H3_o(5) => 
        \SHA256_BLOCK_0_H3_o[5]\, SHA256_BLOCK_0_H3_o(4) => 
        \SHA256_BLOCK_0_H3_o[4]\, SHA256_BLOCK_0_H3_o(3) => 
        \SHA256_BLOCK_0_H3_o[3]\, SHA256_BLOCK_0_H3_o(2) => 
        \SHA256_BLOCK_0_H3_o[2]\, SHA256_BLOCK_0_H3_o(1) => 
        \SHA256_BLOCK_0_H3_o[1]\, SHA256_BLOCK_0_H3_o(0) => 
        \SHA256_BLOCK_0_H3_o[0]\, SHA256_BLOCK_0_H4_o(31) => 
        \SHA256_BLOCK_0_H4_o[31]\, SHA256_BLOCK_0_H4_o(30) => 
        \SHA256_BLOCK_0_H4_o[30]\, SHA256_BLOCK_0_H4_o(29) => 
        \SHA256_BLOCK_0_H4_o[29]\, SHA256_BLOCK_0_H4_o(28) => 
        \SHA256_BLOCK_0_H4_o[28]\, SHA256_BLOCK_0_H4_o(27) => 
        \SHA256_BLOCK_0_H4_o[27]\, SHA256_BLOCK_0_H4_o(26) => 
        \SHA256_BLOCK_0_H4_o[26]\, SHA256_BLOCK_0_H4_o(25) => 
        \SHA256_BLOCK_0_H4_o[25]\, SHA256_BLOCK_0_H4_o(24) => 
        \SHA256_BLOCK_0_H4_o[24]\, SHA256_BLOCK_0_H4_o(23) => 
        \SHA256_BLOCK_0_H4_o[23]\, SHA256_BLOCK_0_H4_o(22) => 
        \SHA256_BLOCK_0_H4_o[22]\, SHA256_BLOCK_0_H4_o(21) => 
        \SHA256_BLOCK_0_H4_o[21]\, SHA256_BLOCK_0_H4_o(20) => 
        \SHA256_BLOCK_0_H4_o[20]\, SHA256_BLOCK_0_H4_o(19) => 
        \SHA256_BLOCK_0_H4_o[19]\, SHA256_BLOCK_0_H4_o(18) => 
        \SHA256_BLOCK_0_H4_o[18]\, SHA256_BLOCK_0_H4_o(17) => 
        \SHA256_BLOCK_0_H4_o[17]\, SHA256_BLOCK_0_H4_o(16) => 
        \SHA256_BLOCK_0_H4_o[16]\, SHA256_BLOCK_0_H4_o(15) => 
        \SHA256_BLOCK_0_H4_o[15]\, SHA256_BLOCK_0_H4_o(14) => 
        \SHA256_BLOCK_0_H4_o[14]\, SHA256_BLOCK_0_H4_o(13) => 
        \SHA256_BLOCK_0_H4_o[13]\, SHA256_BLOCK_0_H4_o(12) => 
        \SHA256_BLOCK_0_H4_o[12]\, SHA256_BLOCK_0_H4_o(11) => 
        \SHA256_BLOCK_0_H4_o[11]\, SHA256_BLOCK_0_H4_o(10) => 
        \SHA256_BLOCK_0_H4_o[10]\, SHA256_BLOCK_0_H4_o(9) => 
        \SHA256_BLOCK_0_H4_o[9]\, SHA256_BLOCK_0_H4_o(8) => 
        \SHA256_BLOCK_0_H4_o[8]\, SHA256_BLOCK_0_H4_o(7) => 
        \SHA256_BLOCK_0_H4_o[7]\, SHA256_BLOCK_0_H4_o(6) => 
        \SHA256_BLOCK_0_H4_o[6]\, SHA256_BLOCK_0_H4_o(5) => 
        \SHA256_BLOCK_0_H4_o[5]\, SHA256_BLOCK_0_H4_o(4) => 
        \SHA256_BLOCK_0_H4_o[4]\, SHA256_BLOCK_0_H4_o(3) => 
        \SHA256_BLOCK_0_H4_o[3]\, SHA256_BLOCK_0_H4_o(2) => 
        \SHA256_BLOCK_0_H4_o[2]\, SHA256_BLOCK_0_H4_o(1) => 
        \SHA256_BLOCK_0_H4_o[1]\, SHA256_BLOCK_0_H4_o(0) => 
        \SHA256_BLOCK_0_H4_o[0]\, SHA256_BLOCK_0_H5_o(31) => 
        \SHA256_BLOCK_0_H5_o[31]\, SHA256_BLOCK_0_H5_o(30) => 
        \SHA256_BLOCK_0_H5_o[30]\, SHA256_BLOCK_0_H5_o(29) => 
        \SHA256_BLOCK_0_H5_o[29]\, SHA256_BLOCK_0_H5_o(28) => 
        \SHA256_BLOCK_0_H5_o[28]\, SHA256_BLOCK_0_H5_o(27) => 
        \SHA256_BLOCK_0_H5_o[27]\, SHA256_BLOCK_0_H5_o(26) => 
        \SHA256_BLOCK_0_H5_o[26]\, SHA256_BLOCK_0_H5_o(25) => 
        \SHA256_BLOCK_0_H5_o[25]\, SHA256_BLOCK_0_H5_o(24) => 
        \SHA256_BLOCK_0_H5_o[24]\, SHA256_BLOCK_0_H5_o(23) => 
        \SHA256_BLOCK_0_H5_o[23]\, SHA256_BLOCK_0_H5_o(22) => 
        \SHA256_BLOCK_0_H5_o[22]\, SHA256_BLOCK_0_H5_o(21) => 
        \SHA256_BLOCK_0_H5_o[21]\, SHA256_BLOCK_0_H5_o(20) => 
        \SHA256_BLOCK_0_H5_o[20]\, SHA256_BLOCK_0_H5_o(19) => 
        \SHA256_BLOCK_0_H5_o[19]\, SHA256_BLOCK_0_H5_o(18) => 
        \SHA256_BLOCK_0_H5_o[18]\, SHA256_BLOCK_0_H5_o(17) => 
        \SHA256_BLOCK_0_H5_o[17]\, SHA256_BLOCK_0_H5_o(16) => 
        \SHA256_BLOCK_0_H5_o[16]\, SHA256_BLOCK_0_H5_o(15) => 
        \SHA256_BLOCK_0_H5_o[15]\, SHA256_BLOCK_0_H5_o(14) => 
        \SHA256_BLOCK_0_H5_o[14]\, SHA256_BLOCK_0_H5_o(13) => 
        \SHA256_BLOCK_0_H5_o[13]\, SHA256_BLOCK_0_H5_o(12) => 
        \SHA256_BLOCK_0_H5_o[12]\, SHA256_BLOCK_0_H5_o(11) => 
        \SHA256_BLOCK_0_H5_o[11]\, SHA256_BLOCK_0_H5_o(10) => 
        \SHA256_BLOCK_0_H5_o[10]\, SHA256_BLOCK_0_H5_o(9) => 
        \SHA256_BLOCK_0_H5_o[9]\, SHA256_BLOCK_0_H5_o(8) => 
        \SHA256_BLOCK_0_H5_o[8]\, SHA256_BLOCK_0_H5_o(7) => 
        \SHA256_BLOCK_0_H5_o[7]\, SHA256_BLOCK_0_H5_o(6) => 
        \SHA256_BLOCK_0_H5_o[6]\, SHA256_BLOCK_0_H5_o(5) => 
        \SHA256_BLOCK_0_H5_o[5]\, SHA256_BLOCK_0_H5_o(4) => 
        \SHA256_BLOCK_0_H5_o[4]\, SHA256_BLOCK_0_H5_o(3) => 
        \SHA256_BLOCK_0_H5_o[3]\, SHA256_BLOCK_0_H5_o(2) => 
        \SHA256_BLOCK_0_H5_o[2]\, SHA256_BLOCK_0_H5_o(1) => 
        \SHA256_BLOCK_0_H5_o[1]\, SHA256_BLOCK_0_H5_o(0) => 
        \SHA256_BLOCK_0_H5_o[0]\, SHA256_BLOCK_0_H6_o(31) => 
        \SHA256_BLOCK_0_H6_o[31]\, SHA256_BLOCK_0_H6_o(30) => 
        \SHA256_BLOCK_0_H6_o[30]\, SHA256_BLOCK_0_H6_o(29) => 
        \SHA256_BLOCK_0_H6_o[29]\, SHA256_BLOCK_0_H6_o(28) => 
        \SHA256_BLOCK_0_H6_o[28]\, SHA256_BLOCK_0_H6_o(27) => 
        \SHA256_BLOCK_0_H6_o[27]\, SHA256_BLOCK_0_H6_o(26) => 
        \SHA256_BLOCK_0_H6_o[26]\, SHA256_BLOCK_0_H6_o(25) => 
        \SHA256_BLOCK_0_H6_o[25]\, SHA256_BLOCK_0_H6_o(24) => 
        \SHA256_BLOCK_0_H6_o[24]\, SHA256_BLOCK_0_H6_o(23) => 
        \SHA256_BLOCK_0_H6_o[23]\, SHA256_BLOCK_0_H6_o(22) => 
        \SHA256_BLOCK_0_H6_o[22]\, SHA256_BLOCK_0_H6_o(21) => 
        \SHA256_BLOCK_0_H6_o[21]\, SHA256_BLOCK_0_H6_o(20) => 
        \SHA256_BLOCK_0_H6_o[20]\, SHA256_BLOCK_0_H6_o(19) => 
        \SHA256_BLOCK_0_H6_o[19]\, SHA256_BLOCK_0_H6_o(18) => 
        \SHA256_BLOCK_0_H6_o[18]\, SHA256_BLOCK_0_H6_o(17) => 
        \SHA256_BLOCK_0_H6_o[17]\, SHA256_BLOCK_0_H6_o(16) => 
        \SHA256_BLOCK_0_H6_o[16]\, SHA256_BLOCK_0_H6_o(15) => 
        \SHA256_BLOCK_0_H6_o[15]\, SHA256_BLOCK_0_H6_o(14) => 
        \SHA256_BLOCK_0_H6_o[14]\, SHA256_BLOCK_0_H6_o(13) => 
        \SHA256_BLOCK_0_H6_o[13]\, SHA256_BLOCK_0_H6_o(12) => 
        \SHA256_BLOCK_0_H6_o[12]\, SHA256_BLOCK_0_H6_o(11) => 
        \SHA256_BLOCK_0_H6_o[11]\, SHA256_BLOCK_0_H6_o(10) => 
        \SHA256_BLOCK_0_H6_o[10]\, SHA256_BLOCK_0_H6_o(9) => 
        \SHA256_BLOCK_0_H6_o[9]\, SHA256_BLOCK_0_H6_o(8) => 
        \SHA256_BLOCK_0_H6_o[8]\, SHA256_BLOCK_0_H6_o(7) => 
        \SHA256_BLOCK_0_H6_o[7]\, SHA256_BLOCK_0_H6_o(6) => 
        \SHA256_BLOCK_0_H6_o[6]\, SHA256_BLOCK_0_H6_o(5) => 
        \SHA256_BLOCK_0_H6_o[5]\, SHA256_BLOCK_0_H6_o(4) => 
        \SHA256_BLOCK_0_H6_o[4]\, SHA256_BLOCK_0_H6_o(3) => 
        \SHA256_BLOCK_0_H6_o[3]\, SHA256_BLOCK_0_H6_o(2) => 
        \SHA256_BLOCK_0_H6_o[2]\, SHA256_BLOCK_0_H6_o(1) => 
        \SHA256_BLOCK_0_H6_o[1]\, SHA256_BLOCK_0_H6_o(0) => 
        \SHA256_BLOCK_0_H6_o[0]\, SHA256_BLOCK_0_H7_o(31) => 
        \SHA256_BLOCK_0_H7_o[31]\, SHA256_BLOCK_0_H7_o(30) => 
        \SHA256_BLOCK_0_H7_o[30]\, SHA256_BLOCK_0_H7_o(29) => 
        \SHA256_BLOCK_0_H7_o[29]\, SHA256_BLOCK_0_H7_o(28) => 
        \SHA256_BLOCK_0_H7_o[28]\, SHA256_BLOCK_0_H7_o(27) => 
        \SHA256_BLOCK_0_H7_o[27]\, SHA256_BLOCK_0_H7_o(26) => 
        \SHA256_BLOCK_0_H7_o[26]\, SHA256_BLOCK_0_H7_o(25) => 
        \SHA256_BLOCK_0_H7_o[25]\, SHA256_BLOCK_0_H7_o(24) => 
        \SHA256_BLOCK_0_H7_o[24]\, SHA256_BLOCK_0_H7_o(23) => 
        \SHA256_BLOCK_0_H7_o[23]\, SHA256_BLOCK_0_H7_o(22) => 
        \SHA256_BLOCK_0_H7_o[22]\, SHA256_BLOCK_0_H7_o(21) => 
        \SHA256_BLOCK_0_H7_o[21]\, SHA256_BLOCK_0_H7_o(20) => 
        \SHA256_BLOCK_0_H7_o[20]\, SHA256_BLOCK_0_H7_o(19) => 
        \SHA256_BLOCK_0_H7_o[19]\, SHA256_BLOCK_0_H7_o(18) => 
        \SHA256_BLOCK_0_H7_o[18]\, SHA256_BLOCK_0_H7_o(17) => 
        \SHA256_BLOCK_0_H7_o[17]\, SHA256_BLOCK_0_H7_o(16) => 
        \SHA256_BLOCK_0_H7_o[16]\, SHA256_BLOCK_0_H7_o(15) => 
        \SHA256_BLOCK_0_H7_o[15]\, SHA256_BLOCK_0_H7_o(14) => 
        \SHA256_BLOCK_0_H7_o[14]\, SHA256_BLOCK_0_H7_o(13) => 
        \SHA256_BLOCK_0_H7_o[13]\, SHA256_BLOCK_0_H7_o(12) => 
        \SHA256_BLOCK_0_H7_o[12]\, SHA256_BLOCK_0_H7_o(11) => 
        \SHA256_BLOCK_0_H7_o[11]\, SHA256_BLOCK_0_H7_o(10) => 
        \SHA256_BLOCK_0_H7_o[10]\, SHA256_BLOCK_0_H7_o(9) => 
        \SHA256_BLOCK_0_H7_o[9]\, SHA256_BLOCK_0_H7_o(8) => 
        \SHA256_BLOCK_0_H7_o[8]\, SHA256_BLOCK_0_H7_o(7) => 
        \SHA256_BLOCK_0_H7_o[7]\, SHA256_BLOCK_0_H7_o(6) => 
        \SHA256_BLOCK_0_H7_o[6]\, SHA256_BLOCK_0_H7_o(5) => 
        \SHA256_BLOCK_0_H7_o[5]\, SHA256_BLOCK_0_H7_o(4) => 
        \SHA256_BLOCK_0_H7_o[4]\, SHA256_BLOCK_0_H7_o(3) => 
        \SHA256_BLOCK_0_H7_o[3]\, SHA256_BLOCK_0_H7_o(2) => 
        \SHA256_BLOCK_0_H7_o[2]\, SHA256_BLOCK_0_H7_o(1) => 
        \SHA256_BLOCK_0_H7_o[1]\, SHA256_BLOCK_0_H7_o(0) => 
        \SHA256_BLOCK_0_H7_o[0]\, AHB_slave_dummy_0_mem_wdata(31)
         => AHB_slave_dummy_0_mem_wdata(31), 
        AHB_slave_dummy_0_mem_wdata(30) => 
        AHB_slave_dummy_0_mem_wdata(30), 
        AHB_slave_dummy_0_mem_wdata(29) => 
        AHB_slave_dummy_0_mem_wdata(29), 
        AHB_slave_dummy_0_mem_wdata(28) => 
        AHB_slave_dummy_0_mem_wdata(28), 
        AHB_slave_dummy_0_mem_wdata(27) => 
        AHB_slave_dummy_0_mem_wdata(27), 
        AHB_slave_dummy_0_mem_wdata(26) => 
        AHB_slave_dummy_0_mem_wdata(26), 
        AHB_slave_dummy_0_mem_wdata(25) => 
        AHB_slave_dummy_0_mem_wdata(25), 
        AHB_slave_dummy_0_mem_wdata(24) => 
        AHB_slave_dummy_0_mem_wdata(24), 
        AHB_slave_dummy_0_mem_wdata(23) => 
        AHB_slave_dummy_0_mem_wdata(23), 
        AHB_slave_dummy_0_mem_wdata(22) => 
        AHB_slave_dummy_0_mem_wdata(22), 
        AHB_slave_dummy_0_mem_wdata(21) => 
        AHB_slave_dummy_0_mem_wdata(21), 
        AHB_slave_dummy_0_mem_wdata(20) => 
        AHB_slave_dummy_0_mem_wdata(20), 
        AHB_slave_dummy_0_mem_wdata(19) => 
        AHB_slave_dummy_0_mem_wdata(19), 
        AHB_slave_dummy_0_mem_wdata(18) => 
        AHB_slave_dummy_0_mem_wdata(18), 
        AHB_slave_dummy_0_mem_wdata(17) => 
        AHB_slave_dummy_0_mem_wdata(17), 
        AHB_slave_dummy_0_mem_wdata(16) => 
        AHB_slave_dummy_0_mem_wdata(16), 
        AHB_slave_dummy_0_mem_wdata(15) => 
        AHB_slave_dummy_0_mem_wdata(15), 
        AHB_slave_dummy_0_mem_wdata(14) => 
        AHB_slave_dummy_0_mem_wdata(14), 
        AHB_slave_dummy_0_mem_wdata(13) => 
        AHB_slave_dummy_0_mem_wdata(13), 
        AHB_slave_dummy_0_mem_wdata(12) => 
        AHB_slave_dummy_0_mem_wdata(12), 
        AHB_slave_dummy_0_mem_wdata(11) => 
        AHB_slave_dummy_0_mem_wdata(11), 
        AHB_slave_dummy_0_mem_wdata(10) => 
        AHB_slave_dummy_0_mem_wdata(10), 
        AHB_slave_dummy_0_mem_wdata(9) => 
        AHB_slave_dummy_0_mem_wdata(9), 
        AHB_slave_dummy_0_mem_wdata(8) => 
        AHB_slave_dummy_0_mem_wdata(8), 
        AHB_slave_dummy_0_mem_wdata(7) => 
        AHB_slave_dummy_0_mem_wdata(7), 
        AHB_slave_dummy_0_mem_wdata(6) => 
        AHB_slave_dummy_0_mem_wdata(6), 
        AHB_slave_dummy_0_mem_wdata(5) => 
        AHB_slave_dummy_0_mem_wdata(5), 
        AHB_slave_dummy_0_mem_wdata(4) => 
        AHB_slave_dummy_0_mem_wdata(4), 
        AHB_slave_dummy_0_mem_wdata(3) => 
        AHB_slave_dummy_0_mem_wdata(3), 
        AHB_slave_dummy_0_mem_wdata(2) => 
        AHB_slave_dummy_0_mem_wdata(2), 
        AHB_slave_dummy_0_mem_wdata(1) => 
        AHB_slave_dummy_0_mem_wdata(1), 
        AHB_slave_dummy_0_mem_wdata(0) => 
        AHB_slave_dummy_0_mem_wdata(0), waddr_in_net_0(4) => 
        waddr_in_net_0(4), waddr_in_net_0(3) => waddr_in_net_0(3), 
        waddr_in_net_0(2) => waddr_in_net_0(2), waddr_in_net_0(1)
         => waddr_in_net_0(1), waddr_in_net_0(0) => 
        waddr_in_net_0(0), state_out_net_0(0) => 
        state_out_net_0(0), sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, SHA256_Module_0_di_req_o
         => \SHA256_Module_0_di_req_o\, 
        SHA256_Module_0_do_valid_o => 
        \SHA256_Module_0_do_valid_o\, SHA256_Module_0_error_o => 
        \SHA256_Module_0_error_o\, SHA256_Module_0_data_out_ready
         => \SHA256_Module_0_data_out_ready\, 
        sha256_system_sb_0_GPIO_9_M2F => 
        sha256_system_sb_0_GPIO_9_M2F, 
        SHA256_Module_0_data_available => 
        SHA256_Module_0_data_available, 
        sha256_system_sb_0_GPIO_1_M2F => 
        sha256_system_sb_0_GPIO_1_M2F, AHB_slave_dummy_0_write_en
         => AHB_slave_dummy_0_write_en, ce_i_i_2_i_0 => 
        ce_i_i_2_i_0, N_88_i_0 => N_88_i_0, N_87_i_0 => N_87_i_0);
    
    reg9_1x32_0 : reg9_1x32
      port map(result_addr_net_0(3) => result_addr_net_0(3), 
        result_addr_net_0(2) => result_addr_net_0(2), 
        result_addr_net_0(1) => result_addr_net_0(1), 
        result_addr_net_0(0) => result_addr_net_0(0), 
        SHA256_BLOCK_0_H0_o(31) => \SHA256_BLOCK_0_H0_o[31]\, 
        SHA256_BLOCK_0_H0_o(30) => \SHA256_BLOCK_0_H0_o[30]\, 
        SHA256_BLOCK_0_H0_o(29) => \SHA256_BLOCK_0_H0_o[29]\, 
        SHA256_BLOCK_0_H0_o(28) => \SHA256_BLOCK_0_H0_o[28]\, 
        SHA256_BLOCK_0_H0_o(27) => \SHA256_BLOCK_0_H0_o[27]\, 
        SHA256_BLOCK_0_H0_o(26) => \SHA256_BLOCK_0_H0_o[26]\, 
        SHA256_BLOCK_0_H0_o(25) => \SHA256_BLOCK_0_H0_o[25]\, 
        SHA256_BLOCK_0_H0_o(24) => \SHA256_BLOCK_0_H0_o[24]\, 
        SHA256_BLOCK_0_H0_o(23) => \SHA256_BLOCK_0_H0_o[23]\, 
        SHA256_BLOCK_0_H0_o(22) => \SHA256_BLOCK_0_H0_o[22]\, 
        SHA256_BLOCK_0_H0_o(21) => \SHA256_BLOCK_0_H0_o[21]\, 
        SHA256_BLOCK_0_H0_o(20) => \SHA256_BLOCK_0_H0_o[20]\, 
        SHA256_BLOCK_0_H0_o(19) => \SHA256_BLOCK_0_H0_o[19]\, 
        SHA256_BLOCK_0_H0_o(18) => \SHA256_BLOCK_0_H0_o[18]\, 
        SHA256_BLOCK_0_H0_o(17) => \SHA256_BLOCK_0_H0_o[17]\, 
        SHA256_BLOCK_0_H0_o(16) => \SHA256_BLOCK_0_H0_o[16]\, 
        SHA256_BLOCK_0_H0_o(15) => \SHA256_BLOCK_0_H0_o[15]\, 
        SHA256_BLOCK_0_H0_o(14) => \SHA256_BLOCK_0_H0_o[14]\, 
        SHA256_BLOCK_0_H0_o(13) => \SHA256_BLOCK_0_H0_o[13]\, 
        SHA256_BLOCK_0_H0_o(12) => \SHA256_BLOCK_0_H0_o[12]\, 
        SHA256_BLOCK_0_H0_o(11) => \SHA256_BLOCK_0_H0_o[11]\, 
        SHA256_BLOCK_0_H0_o(10) => \SHA256_BLOCK_0_H0_o[10]\, 
        SHA256_BLOCK_0_H0_o(9) => \SHA256_BLOCK_0_H0_o[9]\, 
        SHA256_BLOCK_0_H0_o(8) => \SHA256_BLOCK_0_H0_o[8]\, 
        SHA256_BLOCK_0_H0_o(7) => \SHA256_BLOCK_0_H0_o[7]\, 
        SHA256_BLOCK_0_H0_o(6) => \SHA256_BLOCK_0_H0_o[6]\, 
        SHA256_BLOCK_0_H0_o(5) => \SHA256_BLOCK_0_H0_o[5]\, 
        SHA256_BLOCK_0_H0_o(4) => \SHA256_BLOCK_0_H0_o[4]\, 
        SHA256_BLOCK_0_H0_o(3) => \SHA256_BLOCK_0_H0_o[3]\, 
        SHA256_BLOCK_0_H0_o(2) => \SHA256_BLOCK_0_H0_o[2]\, 
        SHA256_BLOCK_0_H0_o(1) => \SHA256_BLOCK_0_H0_o[1]\, 
        SHA256_BLOCK_0_H0_o(0) => \SHA256_BLOCK_0_H0_o[0]\, 
        SHA256_BLOCK_0_H1_o(31) => \SHA256_BLOCK_0_H1_o[31]\, 
        SHA256_BLOCK_0_H1_o(30) => \SHA256_BLOCK_0_H1_o[30]\, 
        SHA256_BLOCK_0_H1_o(29) => \SHA256_BLOCK_0_H1_o[29]\, 
        SHA256_BLOCK_0_H1_o(28) => \SHA256_BLOCK_0_H1_o[28]\, 
        SHA256_BLOCK_0_H1_o(27) => \SHA256_BLOCK_0_H1_o[27]\, 
        SHA256_BLOCK_0_H1_o(26) => \SHA256_BLOCK_0_H1_o[26]\, 
        SHA256_BLOCK_0_H1_o(25) => \SHA256_BLOCK_0_H1_o[25]\, 
        SHA256_BLOCK_0_H1_o(24) => \SHA256_BLOCK_0_H1_o[24]\, 
        SHA256_BLOCK_0_H1_o(23) => \SHA256_BLOCK_0_H1_o[23]\, 
        SHA256_BLOCK_0_H1_o(22) => \SHA256_BLOCK_0_H1_o[22]\, 
        SHA256_BLOCK_0_H1_o(21) => \SHA256_BLOCK_0_H1_o[21]\, 
        SHA256_BLOCK_0_H1_o(20) => \SHA256_BLOCK_0_H1_o[20]\, 
        SHA256_BLOCK_0_H1_o(19) => \SHA256_BLOCK_0_H1_o[19]\, 
        SHA256_BLOCK_0_H1_o(18) => \SHA256_BLOCK_0_H1_o[18]\, 
        SHA256_BLOCK_0_H1_o(17) => \SHA256_BLOCK_0_H1_o[17]\, 
        SHA256_BLOCK_0_H1_o(16) => \SHA256_BLOCK_0_H1_o[16]\, 
        SHA256_BLOCK_0_H1_o(15) => \SHA256_BLOCK_0_H1_o[15]\, 
        SHA256_BLOCK_0_H1_o(14) => \SHA256_BLOCK_0_H1_o[14]\, 
        SHA256_BLOCK_0_H1_o(13) => \SHA256_BLOCK_0_H1_o[13]\, 
        SHA256_BLOCK_0_H1_o(12) => \SHA256_BLOCK_0_H1_o[12]\, 
        SHA256_BLOCK_0_H1_o(11) => \SHA256_BLOCK_0_H1_o[11]\, 
        SHA256_BLOCK_0_H1_o(10) => \SHA256_BLOCK_0_H1_o[10]\, 
        SHA256_BLOCK_0_H1_o(9) => \SHA256_BLOCK_0_H1_o[9]\, 
        SHA256_BLOCK_0_H1_o(8) => \SHA256_BLOCK_0_H1_o[8]\, 
        SHA256_BLOCK_0_H1_o(7) => \SHA256_BLOCK_0_H1_o[7]\, 
        SHA256_BLOCK_0_H1_o(6) => \SHA256_BLOCK_0_H1_o[6]\, 
        SHA256_BLOCK_0_H1_o(5) => \SHA256_BLOCK_0_H1_o[5]\, 
        SHA256_BLOCK_0_H1_o(4) => \SHA256_BLOCK_0_H1_o[4]\, 
        SHA256_BLOCK_0_H1_o(3) => \SHA256_BLOCK_0_H1_o[3]\, 
        SHA256_BLOCK_0_H1_o(2) => \SHA256_BLOCK_0_H1_o[2]\, 
        SHA256_BLOCK_0_H1_o(1) => \SHA256_BLOCK_0_H1_o[1]\, 
        SHA256_BLOCK_0_H1_o(0) => \SHA256_BLOCK_0_H1_o[0]\, 
        SHA256_BLOCK_0_H2_o(31) => \SHA256_BLOCK_0_H2_o[31]\, 
        SHA256_BLOCK_0_H2_o(30) => \SHA256_BLOCK_0_H2_o[30]\, 
        SHA256_BLOCK_0_H2_o(29) => \SHA256_BLOCK_0_H2_o[29]\, 
        SHA256_BLOCK_0_H2_o(28) => \SHA256_BLOCK_0_H2_o[28]\, 
        SHA256_BLOCK_0_H2_o(27) => \SHA256_BLOCK_0_H2_o[27]\, 
        SHA256_BLOCK_0_H2_o(26) => \SHA256_BLOCK_0_H2_o[26]\, 
        SHA256_BLOCK_0_H2_o(25) => \SHA256_BLOCK_0_H2_o[25]\, 
        SHA256_BLOCK_0_H2_o(24) => \SHA256_BLOCK_0_H2_o[24]\, 
        SHA256_BLOCK_0_H2_o(23) => \SHA256_BLOCK_0_H2_o[23]\, 
        SHA256_BLOCK_0_H2_o(22) => \SHA256_BLOCK_0_H2_o[22]\, 
        SHA256_BLOCK_0_H2_o(21) => \SHA256_BLOCK_0_H2_o[21]\, 
        SHA256_BLOCK_0_H2_o(20) => \SHA256_BLOCK_0_H2_o[20]\, 
        SHA256_BLOCK_0_H2_o(19) => \SHA256_BLOCK_0_H2_o[19]\, 
        SHA256_BLOCK_0_H2_o(18) => \SHA256_BLOCK_0_H2_o[18]\, 
        SHA256_BLOCK_0_H2_o(17) => \SHA256_BLOCK_0_H2_o[17]\, 
        SHA256_BLOCK_0_H2_o(16) => \SHA256_BLOCK_0_H2_o[16]\, 
        SHA256_BLOCK_0_H2_o(15) => \SHA256_BLOCK_0_H2_o[15]\, 
        SHA256_BLOCK_0_H2_o(14) => \SHA256_BLOCK_0_H2_o[14]\, 
        SHA256_BLOCK_0_H2_o(13) => \SHA256_BLOCK_0_H2_o[13]\, 
        SHA256_BLOCK_0_H2_o(12) => \SHA256_BLOCK_0_H2_o[12]\, 
        SHA256_BLOCK_0_H2_o(11) => \SHA256_BLOCK_0_H2_o[11]\, 
        SHA256_BLOCK_0_H2_o(10) => \SHA256_BLOCK_0_H2_o[10]\, 
        SHA256_BLOCK_0_H2_o(9) => \SHA256_BLOCK_0_H2_o[9]\, 
        SHA256_BLOCK_0_H2_o(8) => \SHA256_BLOCK_0_H2_o[8]\, 
        SHA256_BLOCK_0_H2_o(7) => \SHA256_BLOCK_0_H2_o[7]\, 
        SHA256_BLOCK_0_H2_o(6) => \SHA256_BLOCK_0_H2_o[6]\, 
        SHA256_BLOCK_0_H2_o(5) => \SHA256_BLOCK_0_H2_o[5]\, 
        SHA256_BLOCK_0_H2_o(4) => \SHA256_BLOCK_0_H2_o[4]\, 
        SHA256_BLOCK_0_H2_o(3) => \SHA256_BLOCK_0_H2_o[3]\, 
        SHA256_BLOCK_0_H2_o(2) => \SHA256_BLOCK_0_H2_o[2]\, 
        SHA256_BLOCK_0_H2_o(1) => \SHA256_BLOCK_0_H2_o[1]\, 
        SHA256_BLOCK_0_H2_o(0) => \SHA256_BLOCK_0_H2_o[0]\, 
        SHA256_BLOCK_0_H3_o(31) => \SHA256_BLOCK_0_H3_o[31]\, 
        SHA256_BLOCK_0_H3_o(30) => \SHA256_BLOCK_0_H3_o[30]\, 
        SHA256_BLOCK_0_H3_o(29) => \SHA256_BLOCK_0_H3_o[29]\, 
        SHA256_BLOCK_0_H3_o(28) => \SHA256_BLOCK_0_H3_o[28]\, 
        SHA256_BLOCK_0_H3_o(27) => \SHA256_BLOCK_0_H3_o[27]\, 
        SHA256_BLOCK_0_H3_o(26) => \SHA256_BLOCK_0_H3_o[26]\, 
        SHA256_BLOCK_0_H3_o(25) => \SHA256_BLOCK_0_H3_o[25]\, 
        SHA256_BLOCK_0_H3_o(24) => \SHA256_BLOCK_0_H3_o[24]\, 
        SHA256_BLOCK_0_H3_o(23) => \SHA256_BLOCK_0_H3_o[23]\, 
        SHA256_BLOCK_0_H3_o(22) => \SHA256_BLOCK_0_H3_o[22]\, 
        SHA256_BLOCK_0_H3_o(21) => \SHA256_BLOCK_0_H3_o[21]\, 
        SHA256_BLOCK_0_H3_o(20) => \SHA256_BLOCK_0_H3_o[20]\, 
        SHA256_BLOCK_0_H3_o(19) => \SHA256_BLOCK_0_H3_o[19]\, 
        SHA256_BLOCK_0_H3_o(18) => \SHA256_BLOCK_0_H3_o[18]\, 
        SHA256_BLOCK_0_H3_o(17) => \SHA256_BLOCK_0_H3_o[17]\, 
        SHA256_BLOCK_0_H3_o(16) => \SHA256_BLOCK_0_H3_o[16]\, 
        SHA256_BLOCK_0_H3_o(15) => \SHA256_BLOCK_0_H3_o[15]\, 
        SHA256_BLOCK_0_H3_o(14) => \SHA256_BLOCK_0_H3_o[14]\, 
        SHA256_BLOCK_0_H3_o(13) => \SHA256_BLOCK_0_H3_o[13]\, 
        SHA256_BLOCK_0_H3_o(12) => \SHA256_BLOCK_0_H3_o[12]\, 
        SHA256_BLOCK_0_H3_o(11) => \SHA256_BLOCK_0_H3_o[11]\, 
        SHA256_BLOCK_0_H3_o(10) => \SHA256_BLOCK_0_H3_o[10]\, 
        SHA256_BLOCK_0_H3_o(9) => \SHA256_BLOCK_0_H3_o[9]\, 
        SHA256_BLOCK_0_H3_o(8) => \SHA256_BLOCK_0_H3_o[8]\, 
        SHA256_BLOCK_0_H3_o(7) => \SHA256_BLOCK_0_H3_o[7]\, 
        SHA256_BLOCK_0_H3_o(6) => \SHA256_BLOCK_0_H3_o[6]\, 
        SHA256_BLOCK_0_H3_o(5) => \SHA256_BLOCK_0_H3_o[5]\, 
        SHA256_BLOCK_0_H3_o(4) => \SHA256_BLOCK_0_H3_o[4]\, 
        SHA256_BLOCK_0_H3_o(3) => \SHA256_BLOCK_0_H3_o[3]\, 
        SHA256_BLOCK_0_H3_o(2) => \SHA256_BLOCK_0_H3_o[2]\, 
        SHA256_BLOCK_0_H3_o(1) => \SHA256_BLOCK_0_H3_o[1]\, 
        SHA256_BLOCK_0_H3_o(0) => \SHA256_BLOCK_0_H3_o[0]\, 
        SHA256_BLOCK_0_H4_o(31) => \SHA256_BLOCK_0_H4_o[31]\, 
        SHA256_BLOCK_0_H4_o(30) => \SHA256_BLOCK_0_H4_o[30]\, 
        SHA256_BLOCK_0_H4_o(29) => \SHA256_BLOCK_0_H4_o[29]\, 
        SHA256_BLOCK_0_H4_o(28) => \SHA256_BLOCK_0_H4_o[28]\, 
        SHA256_BLOCK_0_H4_o(27) => \SHA256_BLOCK_0_H4_o[27]\, 
        SHA256_BLOCK_0_H4_o(26) => \SHA256_BLOCK_0_H4_o[26]\, 
        SHA256_BLOCK_0_H4_o(25) => \SHA256_BLOCK_0_H4_o[25]\, 
        SHA256_BLOCK_0_H4_o(24) => \SHA256_BLOCK_0_H4_o[24]\, 
        SHA256_BLOCK_0_H4_o(23) => \SHA256_BLOCK_0_H4_o[23]\, 
        SHA256_BLOCK_0_H4_o(22) => \SHA256_BLOCK_0_H4_o[22]\, 
        SHA256_BLOCK_0_H4_o(21) => \SHA256_BLOCK_0_H4_o[21]\, 
        SHA256_BLOCK_0_H4_o(20) => \SHA256_BLOCK_0_H4_o[20]\, 
        SHA256_BLOCK_0_H4_o(19) => \SHA256_BLOCK_0_H4_o[19]\, 
        SHA256_BLOCK_0_H4_o(18) => \SHA256_BLOCK_0_H4_o[18]\, 
        SHA256_BLOCK_0_H4_o(17) => \SHA256_BLOCK_0_H4_o[17]\, 
        SHA256_BLOCK_0_H4_o(16) => \SHA256_BLOCK_0_H4_o[16]\, 
        SHA256_BLOCK_0_H4_o(15) => \SHA256_BLOCK_0_H4_o[15]\, 
        SHA256_BLOCK_0_H4_o(14) => \SHA256_BLOCK_0_H4_o[14]\, 
        SHA256_BLOCK_0_H4_o(13) => \SHA256_BLOCK_0_H4_o[13]\, 
        SHA256_BLOCK_0_H4_o(12) => \SHA256_BLOCK_0_H4_o[12]\, 
        SHA256_BLOCK_0_H4_o(11) => \SHA256_BLOCK_0_H4_o[11]\, 
        SHA256_BLOCK_0_H4_o(10) => \SHA256_BLOCK_0_H4_o[10]\, 
        SHA256_BLOCK_0_H4_o(9) => \SHA256_BLOCK_0_H4_o[9]\, 
        SHA256_BLOCK_0_H4_o(8) => \SHA256_BLOCK_0_H4_o[8]\, 
        SHA256_BLOCK_0_H4_o(7) => \SHA256_BLOCK_0_H4_o[7]\, 
        SHA256_BLOCK_0_H4_o(6) => \SHA256_BLOCK_0_H4_o[6]\, 
        SHA256_BLOCK_0_H4_o(5) => \SHA256_BLOCK_0_H4_o[5]\, 
        SHA256_BLOCK_0_H4_o(4) => \SHA256_BLOCK_0_H4_o[4]\, 
        SHA256_BLOCK_0_H4_o(3) => \SHA256_BLOCK_0_H4_o[3]\, 
        SHA256_BLOCK_0_H4_o(2) => \SHA256_BLOCK_0_H4_o[2]\, 
        SHA256_BLOCK_0_H4_o(1) => \SHA256_BLOCK_0_H4_o[1]\, 
        SHA256_BLOCK_0_H4_o(0) => \SHA256_BLOCK_0_H4_o[0]\, 
        SHA256_BLOCK_0_H5_o(31) => \SHA256_BLOCK_0_H5_o[31]\, 
        SHA256_BLOCK_0_H5_o(30) => \SHA256_BLOCK_0_H5_o[30]\, 
        SHA256_BLOCK_0_H5_o(29) => \SHA256_BLOCK_0_H5_o[29]\, 
        SHA256_BLOCK_0_H5_o(28) => \SHA256_BLOCK_0_H5_o[28]\, 
        SHA256_BLOCK_0_H5_o(27) => \SHA256_BLOCK_0_H5_o[27]\, 
        SHA256_BLOCK_0_H5_o(26) => \SHA256_BLOCK_0_H5_o[26]\, 
        SHA256_BLOCK_0_H5_o(25) => \SHA256_BLOCK_0_H5_o[25]\, 
        SHA256_BLOCK_0_H5_o(24) => \SHA256_BLOCK_0_H5_o[24]\, 
        SHA256_BLOCK_0_H5_o(23) => \SHA256_BLOCK_0_H5_o[23]\, 
        SHA256_BLOCK_0_H5_o(22) => \SHA256_BLOCK_0_H5_o[22]\, 
        SHA256_BLOCK_0_H5_o(21) => \SHA256_BLOCK_0_H5_o[21]\, 
        SHA256_BLOCK_0_H5_o(20) => \SHA256_BLOCK_0_H5_o[20]\, 
        SHA256_BLOCK_0_H5_o(19) => \SHA256_BLOCK_0_H5_o[19]\, 
        SHA256_BLOCK_0_H5_o(18) => \SHA256_BLOCK_0_H5_o[18]\, 
        SHA256_BLOCK_0_H5_o(17) => \SHA256_BLOCK_0_H5_o[17]\, 
        SHA256_BLOCK_0_H5_o(16) => \SHA256_BLOCK_0_H5_o[16]\, 
        SHA256_BLOCK_0_H5_o(15) => \SHA256_BLOCK_0_H5_o[15]\, 
        SHA256_BLOCK_0_H5_o(14) => \SHA256_BLOCK_0_H5_o[14]\, 
        SHA256_BLOCK_0_H5_o(13) => \SHA256_BLOCK_0_H5_o[13]\, 
        SHA256_BLOCK_0_H5_o(12) => \SHA256_BLOCK_0_H5_o[12]\, 
        SHA256_BLOCK_0_H5_o(11) => \SHA256_BLOCK_0_H5_o[11]\, 
        SHA256_BLOCK_0_H5_o(10) => \SHA256_BLOCK_0_H5_o[10]\, 
        SHA256_BLOCK_0_H5_o(9) => \SHA256_BLOCK_0_H5_o[9]\, 
        SHA256_BLOCK_0_H5_o(8) => \SHA256_BLOCK_0_H5_o[8]\, 
        SHA256_BLOCK_0_H5_o(7) => \SHA256_BLOCK_0_H5_o[7]\, 
        SHA256_BLOCK_0_H5_o(6) => \SHA256_BLOCK_0_H5_o[6]\, 
        SHA256_BLOCK_0_H5_o(5) => \SHA256_BLOCK_0_H5_o[5]\, 
        SHA256_BLOCK_0_H5_o(4) => \SHA256_BLOCK_0_H5_o[4]\, 
        SHA256_BLOCK_0_H5_o(3) => \SHA256_BLOCK_0_H5_o[3]\, 
        SHA256_BLOCK_0_H5_o(2) => \SHA256_BLOCK_0_H5_o[2]\, 
        SHA256_BLOCK_0_H5_o(1) => \SHA256_BLOCK_0_H5_o[1]\, 
        SHA256_BLOCK_0_H5_o(0) => \SHA256_BLOCK_0_H5_o[0]\, 
        SHA256_BLOCK_0_H6_o(31) => \SHA256_BLOCK_0_H6_o[31]\, 
        SHA256_BLOCK_0_H6_o(30) => \SHA256_BLOCK_0_H6_o[30]\, 
        SHA256_BLOCK_0_H6_o(29) => \SHA256_BLOCK_0_H6_o[29]\, 
        SHA256_BLOCK_0_H6_o(28) => \SHA256_BLOCK_0_H6_o[28]\, 
        SHA256_BLOCK_0_H6_o(27) => \SHA256_BLOCK_0_H6_o[27]\, 
        SHA256_BLOCK_0_H6_o(26) => \SHA256_BLOCK_0_H6_o[26]\, 
        SHA256_BLOCK_0_H6_o(25) => \SHA256_BLOCK_0_H6_o[25]\, 
        SHA256_BLOCK_0_H6_o(24) => \SHA256_BLOCK_0_H6_o[24]\, 
        SHA256_BLOCK_0_H6_o(23) => \SHA256_BLOCK_0_H6_o[23]\, 
        SHA256_BLOCK_0_H6_o(22) => \SHA256_BLOCK_0_H6_o[22]\, 
        SHA256_BLOCK_0_H6_o(21) => \SHA256_BLOCK_0_H6_o[21]\, 
        SHA256_BLOCK_0_H6_o(20) => \SHA256_BLOCK_0_H6_o[20]\, 
        SHA256_BLOCK_0_H6_o(19) => \SHA256_BLOCK_0_H6_o[19]\, 
        SHA256_BLOCK_0_H6_o(18) => \SHA256_BLOCK_0_H6_o[18]\, 
        SHA256_BLOCK_0_H6_o(17) => \SHA256_BLOCK_0_H6_o[17]\, 
        SHA256_BLOCK_0_H6_o(16) => \SHA256_BLOCK_0_H6_o[16]\, 
        SHA256_BLOCK_0_H6_o(15) => \SHA256_BLOCK_0_H6_o[15]\, 
        SHA256_BLOCK_0_H6_o(14) => \SHA256_BLOCK_0_H6_o[14]\, 
        SHA256_BLOCK_0_H6_o(13) => \SHA256_BLOCK_0_H6_o[13]\, 
        SHA256_BLOCK_0_H6_o(12) => \SHA256_BLOCK_0_H6_o[12]\, 
        SHA256_BLOCK_0_H6_o(11) => \SHA256_BLOCK_0_H6_o[11]\, 
        SHA256_BLOCK_0_H6_o(10) => \SHA256_BLOCK_0_H6_o[10]\, 
        SHA256_BLOCK_0_H6_o(9) => \SHA256_BLOCK_0_H6_o[9]\, 
        SHA256_BLOCK_0_H6_o(8) => \SHA256_BLOCK_0_H6_o[8]\, 
        SHA256_BLOCK_0_H6_o(7) => \SHA256_BLOCK_0_H6_o[7]\, 
        SHA256_BLOCK_0_H6_o(6) => \SHA256_BLOCK_0_H6_o[6]\, 
        SHA256_BLOCK_0_H6_o(5) => \SHA256_BLOCK_0_H6_o[5]\, 
        SHA256_BLOCK_0_H6_o(4) => \SHA256_BLOCK_0_H6_o[4]\, 
        SHA256_BLOCK_0_H6_o(3) => \SHA256_BLOCK_0_H6_o[3]\, 
        SHA256_BLOCK_0_H6_o(2) => \SHA256_BLOCK_0_H6_o[2]\, 
        SHA256_BLOCK_0_H6_o(1) => \SHA256_BLOCK_0_H6_o[1]\, 
        SHA256_BLOCK_0_H6_o(0) => \SHA256_BLOCK_0_H6_o[0]\, 
        SHA256_BLOCK_0_H7_o(31) => \SHA256_BLOCK_0_H7_o[31]\, 
        SHA256_BLOCK_0_H7_o(30) => \SHA256_BLOCK_0_H7_o[30]\, 
        SHA256_BLOCK_0_H7_o(29) => \SHA256_BLOCK_0_H7_o[29]\, 
        SHA256_BLOCK_0_H7_o(28) => \SHA256_BLOCK_0_H7_o[28]\, 
        SHA256_BLOCK_0_H7_o(27) => \SHA256_BLOCK_0_H7_o[27]\, 
        SHA256_BLOCK_0_H7_o(26) => \SHA256_BLOCK_0_H7_o[26]\, 
        SHA256_BLOCK_0_H7_o(25) => \SHA256_BLOCK_0_H7_o[25]\, 
        SHA256_BLOCK_0_H7_o(24) => \SHA256_BLOCK_0_H7_o[24]\, 
        SHA256_BLOCK_0_H7_o(23) => \SHA256_BLOCK_0_H7_o[23]\, 
        SHA256_BLOCK_0_H7_o(22) => \SHA256_BLOCK_0_H7_o[22]\, 
        SHA256_BLOCK_0_H7_o(21) => \SHA256_BLOCK_0_H7_o[21]\, 
        SHA256_BLOCK_0_H7_o(20) => \SHA256_BLOCK_0_H7_o[20]\, 
        SHA256_BLOCK_0_H7_o(19) => \SHA256_BLOCK_0_H7_o[19]\, 
        SHA256_BLOCK_0_H7_o(18) => \SHA256_BLOCK_0_H7_o[18]\, 
        SHA256_BLOCK_0_H7_o(17) => \SHA256_BLOCK_0_H7_o[17]\, 
        SHA256_BLOCK_0_H7_o(16) => \SHA256_BLOCK_0_H7_o[16]\, 
        SHA256_BLOCK_0_H7_o(15) => \SHA256_BLOCK_0_H7_o[15]\, 
        SHA256_BLOCK_0_H7_o(14) => \SHA256_BLOCK_0_H7_o[14]\, 
        SHA256_BLOCK_0_H7_o(13) => \SHA256_BLOCK_0_H7_o[13]\, 
        SHA256_BLOCK_0_H7_o(12) => \SHA256_BLOCK_0_H7_o[12]\, 
        SHA256_BLOCK_0_H7_o(11) => \SHA256_BLOCK_0_H7_o[11]\, 
        SHA256_BLOCK_0_H7_o(10) => \SHA256_BLOCK_0_H7_o[10]\, 
        SHA256_BLOCK_0_H7_o(9) => \SHA256_BLOCK_0_H7_o[9]\, 
        SHA256_BLOCK_0_H7_o(8) => \SHA256_BLOCK_0_H7_o[8]\, 
        SHA256_BLOCK_0_H7_o(7) => \SHA256_BLOCK_0_H7_o[7]\, 
        SHA256_BLOCK_0_H7_o(6) => \SHA256_BLOCK_0_H7_o[6]\, 
        SHA256_BLOCK_0_H7_o(5) => \SHA256_BLOCK_0_H7_o[5]\, 
        SHA256_BLOCK_0_H7_o(4) => \SHA256_BLOCK_0_H7_o[4]\, 
        SHA256_BLOCK_0_H7_o(3) => \SHA256_BLOCK_0_H7_o[3]\, 
        SHA256_BLOCK_0_H7_o(2) => \SHA256_BLOCK_0_H7_o[2]\, 
        SHA256_BLOCK_0_H7_o(1) => \SHA256_BLOCK_0_H7_o[1]\, 
        SHA256_BLOCK_0_H7_o(0) => \SHA256_BLOCK_0_H7_o[0]\, 
        line_7_d0 => line_0_d0, line_10 => line_3_d0, line_11 => 
        line_4_d0, line_20 => line_13, line_28 => line_21, 
        line_31 => line_24, line_0_7 => line_0_0, line_0_10 => 
        line_0_3, line_0_11 => line_0_4, line_0_20 => line_0_13, 
        line_0_28 => line_0_21, line_0_31 => line_0_24, line_1_7
         => line_1_0, line_1_10 => line_1_3, line_1_11 => 
        line_1_4, line_1_20 => line_1_13, line_1_28 => line_1_21, 
        line_1_31 => line_1_24, line_2_7 => line_2_0, line_2_10
         => line_2_3, line_2_11 => line_2_4, line_2_20 => 
        line_2_13, line_2_28 => line_2_21, line_2_31 => line_2_24, 
        line_3_7 => line_3_0, line_3_10 => line_3_3, line_3_11
         => line_3_4, line_3_20 => line_3_13, line_3_28 => 
        line_3_21, line_3_31 => line_3_24, line_4_7 => line_4_0, 
        line_4_10 => line_4_3, line_4_11 => line_4_4, line_4_20
         => line_4_13, line_4_28 => line_4_21, line_4_31 => 
        line_4_24, line_5_7 => line_5_0, line_5_10 => line_5_3, 
        line_5_11 => line_5_4, line_5_20 => line_5_13, line_5_28
         => line_5_21, line_5_31 => line_5_24, line_6_7 => 
        line_6_0, line_6_10 => line_6_3, line_6_11 => line_6_4, 
        line_6_20 => line_6_13, line_6_28 => line_6_21, line_6_31
         => line_6_24, line_7_28 => line_7_21, line_7_20 => 
        line_7_13, line_7_11 => line_7_4, line_7_10 => line_7_3, 
        line_7_7 => line_7_0, N_568 => N_568, N_579 => N_579, 
        N_580 => N_580, N_581 => N_581, N_583 => N_583, N_588 => 
        N_588, N_589 => N_589, N_590 => N_590, N_591 => N_591, 
        N_592 => N_592, N_595 => N_595, N_594 => N_594, N_586 => 
        N_586, N_582 => N_582, N_578 => N_578, N_574 => N_574, 
        N_571 => N_571, N_570 => N_570, N_569 => N_569, N_96 => 
        N_96, N_81 => N_81, N_74 => N_74, N_75 => N_75, N_499 => 
        N_499, N_501 => N_501, N_525 => N_525, N_513 => N_513, 
        N_502 => N_502, N_522 => N_522, N_500 => N_500, N_514 => 
        N_514, N_515 => N_515, N_524 => N_524, N_526 => N_526, 
        N_529 => N_529, N_528 => N_528, N_523 => N_523, N_517 => 
        N_517, N_505 => N_505, N_503 => N_503, N_512 => N_512, 
        N_508 => N_508, N_504 => N_504, N_520 => N_520, N_516 => 
        N_516, ren_pos => ren_pos, N_228 => N_228, N_7 => N_7, 
        N_566 => N_566, N_567 => N_567, N_565 => N_565, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, 
        SHA256_Module_0_data_out_ready => 
        \SHA256_Module_0_data_out_ready\, 
        AHB_slave_dummy_0_read_en => AHB_slave_dummy_0_read_en, 
        SHA256_Module_0_do_valid_o => 
        \SHA256_Module_0_do_valid_o\, prev_sig => prev_sig, 
        SHA256_Module_0_error_o => \SHA256_Module_0_error_o\, 
        SHA256_Module_0_di_req_o => \SHA256_Module_0_di_req_o\, 
        SHA256_Module_0_data_available_lastbank_8 => 
        SHA256_Module_0_data_available_lastbank_8);
    
    limiter_1cycle_0 : limiter_1cycle
      port map(prev_sig => prev_sig, sha256_system_sb_0_FIC_0_CLK
         => sha256_system_sb_0_FIC_0_CLK, 
        SHA256_Module_0_do_valid_o => 
        \SHA256_Module_0_do_valid_o\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity AHB_slave_dummy is

    port( waddr_in_net_0                                     : out   std_logic_vector(4 downto 0);
          result_addr_net_0                                  : out   std_logic_vector(3 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS : in    std_logic_vector(1 to 1);
          arbRegSMCurrentState                               : in    std_logic_vector(15 downto 14);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR  : in    std_logic_vector(25 downto 24);
          sha256_system_sb_0_POWER_ON_RESET_N                : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                       : in    std_logic;
          N_118                                              : in    std_logic;
          N_117                                              : in    std_logic;
          N_116                                              : in    std_logic;
          N_115                                              : in    std_logic;
          N_114                                              : in    std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY             : out   std_logic;
          AHB_slave_dummy_0_write_en                         : out   std_logic;
          AHB_slave_dummy_0_read_en                          : out   std_logic;
          N_119                                              : in    std_logic;
          masterRegAddrSel                                   : in    std_logic;
          regHTRANS                                          : in    std_logic;
          N_165                                              : in    std_logic;
          N_14_i                                             : in    std_logic;
          N_164                                              : in    std_logic;
          defSlaveSMCurrentState                             : in    std_logic;
          N_31                                               : in    std_logic
        );

end AHB_slave_dummy;

architecture DEF_ARCH of AHB_slave_dummy is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, lsram_waddr_0_sqmuxa, GND_net_1, N_58_i_0, 
        \sha256_system_sb_0_AMBA_SLAVE_0_HREADY\, \ready_ldmx\, 
        N_157_i_0, \AHB_slave_dummy_0_write_en\, \write_en_ldmx\, 
        \AHB_slave_dummy_0_read_en\, \read_en_ldmx\, \hwrite_r\, 
        N_62_i_0, \FSM[0]_net_1\, \FSM[1]_net_1\, \FSM_ns[1]\, 
        lsram_raddr_1_sqmuxa_i_o2_4_a3_0, 
        \lsram_raddr_1_sqmuxa_i_o2_4_a4\, 
        \lsram_waddr_0_sqmuxa_0_a2_1\, 
        \lsram_raddr_1_sqmuxa_i_o2_1_0\, 
        \lsram_raddr_1_sqmuxa_i_o2_1_2\, N_97, N_100 : std_logic;

begin 

    sha256_system_sb_0_AMBA_SLAVE_0_HREADY <= 
        \sha256_system_sb_0_AMBA_SLAVE_0_HREADY\;
    AHB_slave_dummy_0_write_en <= \AHB_slave_dummy_0_write_en\;
    AHB_slave_dummy_0_read_en <= \AHB_slave_dummy_0_read_en\;

    lsram_waddr_0_sqmuxa_0_a2_1 : CFG3
      generic map(INIT => x"04")

      port map(A => \FSM[0]_net_1\, B => N_119, C => 
        \FSM[1]_net_1\, Y => \lsram_waddr_0_sqmuxa_0_a2_1\);
    
    ready_ldmx : CFG4
      generic map(INIT => x"F4A0")

      port map(A => \FSM_ns[1]\, B => N_119, C => \FSM[0]_net_1\, 
        D => \sha256_system_sb_0_AMBA_SLAVE_0_HREADY\, Y => 
        \ready_ldmx\);
    
    lsram_raddr_1_sqmuxa_i_o2_1_2 : CFG4
      generic map(INIT => x"EEEA")

      port map(A => \lsram_raddr_1_sqmuxa_i_o2_1_0\, B => 
        lsram_raddr_1_sqmuxa_i_o2_4_a3_0, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(25), D
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(24), 
        Y => \lsram_raddr_1_sqmuxa_i_o2_1_2\);
    
    \lsram_raddr[2]\ : SLE
      port map(D => N_116, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_58_i_0, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => result_addr_net_0(2));
    
    hwrite_r : SLE
      port map(D => N_119, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_62_i_0, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \hwrite_r\);
    
    \FSM[1]\ : SLE
      port map(D => \FSM_ns[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \FSM[1]_net_1\);
    
    \lsram_waddr[0]\ : SLE
      port map(D => N_118, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => lsram_waddr_0_sqmuxa, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => waddr_in_net_0(0));
    
    lsram_raddr_1_sqmuxa_i_o2_RNI9R3M_0 : CFG2
      generic map(INIT => x"1")

      port map(A => N_100, B => \FSM[0]_net_1\, Y => N_62_i_0);
    
    write_en_ldmx : CFG4
      generic map(INIT => x"CC54")

      port map(A => \FSM[0]_net_1\, B => 
        \AHB_slave_dummy_0_write_en\, C => N_119, D => 
        \FSM_ns[1]\, Y => \write_en_ldmx\);
    
    lsram_raddr_1_sqmuxa_i_o2_4_a4 : CFG3
      generic map(INIT => x"51")

      port map(A => N_165, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), C
         => masterRegAddrSel, Y => 
        \lsram_raddr_1_sqmuxa_i_o2_4_a4\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \lsram_raddr[1]\ : SLE
      port map(D => N_117, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_58_i_0, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => result_addr_net_0(1));
    
    lsram_raddr_1_sqmuxa_i_o2_1 : CFG4
      generic map(INIT => x"FFBA")

      port map(A => \lsram_raddr_1_sqmuxa_i_o2_1_2\, B => N_164, 
        C => lsram_raddr_1_sqmuxa_i_o2_4_a3_0, D => 
        \lsram_raddr_1_sqmuxa_i_o2_4_a4\, Y => N_97);
    
    \lsram_waddr[1]\ : SLE
      port map(D => N_117, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => lsram_waddr_0_sqmuxa, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => waddr_in_net_0(1));
    
    \lsram_raddr[0]\ : SLE
      port map(D => N_118, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_58_i_0, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => result_addr_net_0(0));
    
    lsram_raddr_1_sqmuxa_i_o2 : CFG4
      generic map(INIT => x"FCFE")

      port map(A => N_31, B => N_97, C => \FSM[1]_net_1\, D => 
        defSlaveSMCurrentState, Y => N_100);
    
    \lsram_waddr[3]\ : SLE
      port map(D => N_115, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => lsram_waddr_0_sqmuxa, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => waddr_in_net_0(3));
    
    \FSM_ns_0_a2_0_a2[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \FSM[0]_net_1\, B => \hwrite_r\, Y => 
        \FSM_ns[1]\);
    
    \FSM[0]\ : SLE
      port map(D => N_62_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \FSM[0]_net_1\);
    
    lsram_raddr_1_sqmuxa_i_o2_RNI7O441 : CFG3
      generic map(INIT => x"01")

      port map(A => N_100, B => \FSM[0]_net_1\, C => N_119, Y => 
        N_58_i_0);
    
    lsram_raddr_1_sqmuxa_i_o2_1_0 : CFG4
      generic map(INIT => x"3337")

      port map(A => N_14_i, B => 
        \sha256_system_sb_0_AMBA_SLAVE_0_HREADY\, C => 
        arbRegSMCurrentState(15), D => arbRegSMCurrentState(14), 
        Y => \lsram_raddr_1_sqmuxa_i_o2_1_0\);
    
    write_en : SLE
      port map(D => \write_en_ldmx\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_157_i_0, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AHB_slave_dummy_0_write_en\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    lsram_raddr_1_sqmuxa_i_o2_RNI9R3M : CFG2
      generic map(INIT => x"D")

      port map(A => N_100, B => \FSM[0]_net_1\, Y => N_157_i_0);
    
    read_en : SLE
      port map(D => \read_en_ldmx\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_157_i_0, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AHB_slave_dummy_0_read_en\);
    
    ready : SLE
      port map(D => \ready_ldmx\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_157_i_0, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sha256_system_sb_0_AMBA_SLAVE_0_HREADY\);
    
    lsram_waddr_0_sqmuxa_0_a2 : CFG4
      generic map(INIT => x"0B00")

      port map(A => defSlaveSMCurrentState, B => N_31, C => N_97, 
        D => \lsram_waddr_0_sqmuxa_0_a2_1\, Y => 
        lsram_waddr_0_sqmuxa);
    
    \lsram_raddr[3]\ : SLE
      port map(D => N_115, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_58_i_0, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => result_addr_net_0(3));
    
    \lsram_waddr[4]\ : SLE
      port map(D => N_114, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => lsram_waddr_0_sqmuxa, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => waddr_in_net_0(4));
    
    \lsram_waddr[2]\ : SLE
      port map(D => N_116, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => lsram_waddr_0_sqmuxa, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => waddr_in_net_0(2));
    
    read_en_ldmx : CFG4
      generic map(INIT => x"55CD")

      port map(A => \FSM[0]_net_1\, B => 
        \AHB_slave_dummy_0_read_en\, C => N_119, D => \FSM_ns[1]\, 
        Y => \read_en_ldmx\);
    
    lsram_raddr_1_sqmuxa_i_o2_4_a1_0 : CFG3
      generic map(INIT => x"15")

      port map(A => arbRegSMCurrentState(15), B => 
        masterRegAddrSel, C => regHTRANS, Y => 
        lsram_raddr_1_sqmuxa_i_o2_4_a3_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_system_sb_MSS is

    port( result_addr_net_0                                    : in    std_logic_vector(2 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : out   std_logic_vector(1 to 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : out   std_logic_vector(31 downto 0);
          state_out_net_0                                      : in    std_logic_vector(0 to 0);
          line_4_d0                                            : in    std_logic;
          line_21                                              : in    std_logic;
          line_3_d0                                            : in    std_logic;
          line_13                                              : in    std_logic;
          line_0_d0                                            : in    std_logic;
          line_24                                              : in    std_logic;
          line_0_4                                             : in    std_logic;
          line_0_21                                            : in    std_logic;
          line_0_3                                             : in    std_logic;
          line_0_13                                            : in    std_logic;
          line_0_0                                             : in    std_logic;
          line_0_24                                            : in    std_logic;
          line_1_4                                             : in    std_logic;
          line_1_21                                            : in    std_logic;
          line_1_3                                             : in    std_logic;
          line_1_13                                            : in    std_logic;
          line_1_0                                             : in    std_logic;
          line_1_24                                            : in    std_logic;
          line_2_4                                             : in    std_logic;
          line_2_21                                            : in    std_logic;
          line_2_3                                             : in    std_logic;
          line_2_13                                            : in    std_logic;
          line_2_0                                             : in    std_logic;
          line_2_24                                            : in    std_logic;
          line_3_3                                             : in    std_logic;
          line_3_21                                            : in    std_logic;
          line_3_0                                             : in    std_logic;
          line_3_4                                             : in    std_logic;
          line_3_24                                            : in    std_logic;
          line_3_13                                            : in    std_logic;
          line_4_3                                             : in    std_logic;
          line_4_21                                            : in    std_logic;
          line_4_0                                             : in    std_logic;
          line_4_4                                             : in    std_logic;
          line_4_24                                            : in    std_logic;
          line_4_13                                            : in    std_logic;
          line_5_3                                             : in    std_logic;
          line_5_21                                            : in    std_logic;
          line_5_0                                             : in    std_logic;
          line_5_4                                             : in    std_logic;
          line_5_24                                            : in    std_logic;
          line_5_13                                            : in    std_logic;
          line_6_3                                             : in    std_logic;
          line_6_21                                            : in    std_logic;
          line_6_0                                             : in    std_logic;
          line_6_4                                             : in    std_logic;
          line_6_24                                            : in    std_logic;
          line_6_13                                            : in    std_logic;
          line_7_3                                             : in    std_logic;
          line_7_0                                             : in    std_logic;
          line_7_13                                            : in    std_logic;
          line_7_4                                             : in    std_logic;
          line_7_21                                            : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_26 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_27 : out   std_logic;
          N_96                                                 : in    std_logic;
          hready_m_xhdl339                                     : in    std_logic;
          ren_pos                                              : in    std_logic;
          N_516                                                : in    std_logic;
          N_582                                                : in    std_logic;
          N_520                                                : in    std_logic;
          N_586                                                : in    std_logic;
          N_504                                                : in    std_logic;
          N_570                                                : in    std_logic;
          N_508                                                : in    std_logic;
          N_574                                                : in    std_logic;
          N_512                                                : in    std_logic;
          N_578                                                : in    std_logic;
          N_503                                                : in    std_logic;
          N_569                                                : in    std_logic;
          N_505                                                : in    std_logic;
          N_571                                                : in    std_logic;
          N_517                                                : in    std_logic;
          N_583                                                : in    std_logic;
          N_523                                                : in    std_logic;
          N_589                                                : in    std_logic;
          N_528                                                : in    std_logic;
          N_594                                                : in    std_logic;
          N_529                                                : in    std_logic;
          N_595                                                : in    std_logic;
          N_526                                                : in    std_logic;
          N_592                                                : in    std_logic;
          N_524                                                : in    std_logic;
          N_590                                                : in    std_logic;
          N_515                                                : in    std_logic;
          N_581                                                : in    std_logic;
          N_514                                                : in    std_logic;
          N_580                                                : in    std_logic;
          N_522                                                : in    std_logic;
          N_588                                                : in    std_logic;
          N_502                                                : in    std_logic;
          N_568                                                : in    std_logic;
          N_513                                                : in    std_logic;
          N_579                                                : in    std_logic;
          N_525                                                : in    std_logic;
          N_591                                                : in    std_logic;
          N_500                                                : in    std_logic;
          N_566                                                : in    std_logic;
          N_501                                                : in    std_logic;
          N_567                                                : in    std_logic;
          N_499                                                : in    std_logic;
          N_565                                                : in    std_logic;
          N_74                                                 : in    std_logic;
          N_228                                                : in    std_logic;
          N_81                                                 : in    std_logic;
          N_7                                                  : in    std_logic;
          N_75                                                 : in    std_logic;
          N_274                                                : in    std_logic;
          N_273                                                : in    std_logic;
          N_59                                                 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N      : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : out   std_logic;
          sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F           : out   std_logic;
          sha256_system_sb_0_GPIO_1_M2F                        : out   std_logic;
          GPIO_0_M2F_c                                         : out   std_logic;
          sha256_system_sb_0_GPIO_9_M2F                        : out   std_logic;
          N_23_i_0                                             : in    std_logic;
          N_31                                                 : in    std_logic;
          FIC_0_LOCK                                           : in    std_logic;
          N_87_i_0                                             : in    std_logic;
          N_88_i_0                                             : in    std_logic;
          ce_i_i_2_i_0                                         : in    std_logic;
          SHA256_Module_0_data_available_lastbank_8            : in    std_logic;
          SHA256_Module_0_di_req_o                             : in    std_logic;
          SHA256_Module_0_data_out_ready                       : in    std_logic;
          SHA256_Module_0_do_valid_o                           : in    std_logic;
          SHA256_Module_0_data_available                       : in    std_logic;
          SHA256_Module_0_error_o                              : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic
        );

end sha256_system_sb_MSS;

architecture DEF_ARCH of sha256_system_sb_MSS is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MSS_060

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MGPIO0B_IN                              : in    std_logic := 'U';
          MGPIO10B_IN                             : in    std_logic := 'U';
          MGPIO1B_IN                              : in    std_logic := 'U';
          MGPIO25A_IN                             : in    std_logic := 'U';
          MGPIO26A_IN                             : in    std_logic := 'U';
          MGPIO27A_IN                             : in    std_logic := 'U';
          MGPIO28A_IN                             : in    std_logic := 'U';
          MGPIO29A_IN                             : in    std_logic := 'U';
          MGPIO2B_IN                              : in    std_logic := 'U';
          MGPIO30A_IN                             : in    std_logic := 'U';
          MGPIO31A_IN                             : in    std_logic := 'U';
          MGPIO3B_IN                              : in    std_logic := 'U';
          MGPIO4B_IN                              : in    std_logic := 'U';
          MGPIO5B_IN                              : in    std_logic := 'U';
          MGPIO6B_IN                              : in    std_logic := 'U';
          MGPIO7B_IN                              : in    std_logic := 'U';
          MGPIO8B_IN                              : in    std_logic := 'U';
          MGPIO9B_IN                              : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_CTS_MGPIO13B_IN                 : in    std_logic := 'U';
          MMUART1_DCD_MGPIO16B_IN                 : in    std_logic := 'U';
          MMUART1_DSR_MGPIO14B_IN                 : in    std_logic := 'U';
          MMUART1_DTR_MGPIO12B_IN                 : in    std_logic := 'U';
          MMUART1_RI_MGPIO15B_IN                  : in    std_logic := 'U';
          MMUART1_RTS_MGPIO11B_IN                 : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI0_SS4_MGPIO19A_IN                    : in    std_logic := 'U';
          SPI0_SS5_MGPIO20A_IN                    : in    std_logic := 'U';
          SPI0_SS6_MGPIO21A_IN                    : in    std_logic := 'U';
          SPI0_SS7_MGPIO22A_IN                    : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          USBD_DATA0_IN                           : in    std_logic := 'U';
          USBD_DATA1_IN                           : in    std_logic := 'U';
          USBD_DATA2_IN                           : in    std_logic := 'U';
          USBD_DATA3_IN                           : in    std_logic := 'U';
          USBD_DATA4_IN                           : in    std_logic := 'U';
          USBD_DATA5_IN                           : in    std_logic := 'U';
          USBD_DATA6_IN                           : in    std_logic := 'U';
          USBD_DATA7_MGPIO23B_IN                  : in    std_logic := 'U';
          USBD_DIR_IN                             : in    std_logic := 'U';
          USBD_NXT_IN                             : in    std_logic := 'U';
          USBD_STP_IN                             : in    std_logic := 'U';
          USBD_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MGPIO0B_OUT                             : out   std_logic;
          MGPIO10B_OUT                            : out   std_logic;
          MGPIO1B_OUT                             : out   std_logic;
          MGPIO25A_OUT                            : out   std_logic;
          MGPIO26A_OUT                            : out   std_logic;
          MGPIO27A_OUT                            : out   std_logic;
          MGPIO28A_OUT                            : out   std_logic;
          MGPIO29A_OUT                            : out   std_logic;
          MGPIO2B_OUT                             : out   std_logic;
          MGPIO30A_OUT                            : out   std_logic;
          MGPIO31A_OUT                            : out   std_logic;
          MGPIO3B_OUT                             : out   std_logic;
          MGPIO4B_OUT                             : out   std_logic;
          MGPIO5B_OUT                             : out   std_logic;
          MGPIO6B_OUT                             : out   std_logic;
          MGPIO7B_OUT                             : out   std_logic;
          MGPIO8B_OUT                             : out   std_logic;
          MGPIO9B_OUT                             : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_CTS_MGPIO13B_OUT                : out   std_logic;
          MMUART1_DCD_MGPIO16B_OUT                : out   std_logic;
          MMUART1_DSR_MGPIO14B_OUT                : out   std_logic;
          MMUART1_DTR_MGPIO12B_OUT                : out   std_logic;
          MMUART1_RI_MGPIO15B_OUT                 : out   std_logic;
          MMUART1_RTS_MGPIO11B_OUT                : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI0_SS4_MGPIO19A_OUT                   : out   std_logic;
          SPI0_SS5_MGPIO20A_OUT                   : out   std_logic;
          SPI0_SS6_MGPIO21A_OUT                   : out   std_logic;
          SPI0_SS7_MGPIO22A_OUT                   : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          USBD_DATA0_OUT                          : out   std_logic;
          USBD_DATA1_OUT                          : out   std_logic;
          USBD_DATA2_OUT                          : out   std_logic;
          USBD_DATA3_OUT                          : out   std_logic;
          USBD_DATA4_OUT                          : out   std_logic;
          USBD_DATA5_OUT                          : out   std_logic;
          USBD_DATA6_OUT                          : out   std_logic;
          USBD_DATA7_MGPIO23B_OUT                 : out   std_logic;
          USBD_DIR_OUT                            : out   std_logic;
          USBD_NXT_OUT                            : out   std_logic;
          USBD_STP_OUT                            : out   std_logic;
          USBD_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MGPIO0B_OE                              : out   std_logic;
          MGPIO10B_OE                             : out   std_logic;
          MGPIO1B_OE                              : out   std_logic;
          MGPIO25A_OE                             : out   std_logic;
          MGPIO26A_OE                             : out   std_logic;
          MGPIO27A_OE                             : out   std_logic;
          MGPIO28A_OE                             : out   std_logic;
          MGPIO29A_OE                             : out   std_logic;
          MGPIO2B_OE                              : out   std_logic;
          MGPIO30A_OE                             : out   std_logic;
          MGPIO31A_OE                             : out   std_logic;
          MGPIO3B_OE                              : out   std_logic;
          MGPIO4B_OE                              : out   std_logic;
          MGPIO5B_OE                              : out   std_logic;
          MGPIO6B_OE                              : out   std_logic;
          MGPIO7B_OE                              : out   std_logic;
          MGPIO8B_OE                              : out   std_logic;
          MGPIO9B_OE                              : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_CTS_MGPIO13B_OE                 : out   std_logic;
          MMUART1_DCD_MGPIO16B_OE                 : out   std_logic;
          MMUART1_DSR_MGPIO14B_OE                 : out   std_logic;
          MMUART1_DTR_MGPIO12B_OE                 : out   std_logic;
          MMUART1_RI_MGPIO15B_OE                  : out   std_logic;
          MMUART1_RTS_MGPIO11B_OE                 : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI0_SS4_MGPIO19A_OE                    : out   std_logic;
          SPI0_SS5_MGPIO20A_OE                    : out   std_logic;
          SPI0_SS6_MGPIO21A_OE                    : out   std_logic;
          SPI0_SS7_MGPIO22A_OE                    : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic;
          USBD_DATA0_OE                           : out   std_logic;
          USBD_DATA1_OE                           : out   std_logic;
          USBD_DATA2_OE                           : out   std_logic;
          USBD_DATA3_OE                           : out   std_logic;
          USBD_DATA4_OE                           : out   std_logic;
          USBD_DATA5_OE                           : out   std_logic;
          USBD_DATA6_OE                           : out   std_logic;
          USBD_DATA7_MGPIO23B_OE                  : out   std_logic;
          USBD_DIR_OE                             : out   std_logic;
          USBD_NXT_OE                             : out   std_logic;
          USBD_STP_OE                             : out   std_logic;
          USBD_XCLK_OE                            : out   std_logic
        );
  end component;

    signal \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[11]\, N_243, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[28]\, N_252, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[10]\, N_188, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[10]\, N_196, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[20]\, N_199, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[7]\, N_240, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[28]\, N_249, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[31]\, N_208, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[7]\, N_237, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[11]\, N_246, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[31]\, N_205, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[20]\, N_202, 
        \AMBA_SLAVE_0_HRDATA_S0_m[22]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[17]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[21]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[5]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[9]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[13]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[4]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[6]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[18]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[24]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[29]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[30]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[27]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[25]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[16]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[15]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[23]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[3]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[14]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[26]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[1]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[2]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[0]\, N_34_i_0, N_35_i_0, 
        N_25_i_0, \AMBA_SLAVE_0_HRDATA_S0_m_0_0[10]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_0[7]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_0[20]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_0[11]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_0[28]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[31]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[7]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[11]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[28]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[10]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[20]\, VCC_net_1, GND_net_1
         : std_logic;
    signal nc228, nc203, nc265, nc216, nc194, nc151, nc23, nc175, 
        nc250, nc58, nc116, nc74, nc133, nc238, nc167, nc84, nc39, 
        nc72, nc256, nc212, nc205, nc82, nc145, nc181, nc160, 
        nc57, nc156, nc280, nc125, nc211, nc73, nc107, nc329, 
        nc66, nc83, nc9, nc252, nc171, nc54, nc286, nc307, nc135, 
        nc41, nc100, nc270, nc52, nc251, nc186, nc29, nc269, 
        nc118, nc60, nc141, nc311, nc276, nc193, nc214, nc298, 
        nc282, nc240, nc45, nc53, nc121, nc176, nc220, nc158, 
        nc281, nc209, nc246, nc162, nc11, nc272, nc131, nc254, 
        nc267, nc96, nc79, nc226, nc146, nc230, nc89, nc119, nc48, 
        nc271, nc213, nc300, nc126, nc195, nc188, nc242, nc15, 
        nc308, nc236, nc102, nc304, nc3, nc207, nc47, nc90, nc284, 
        nc222, nc159, nc136, nc241, nc253, nc178, nc306, nc215, 
        nc59, nc221, nc232, nc274, nc18, nc44, nc117, nc189, 
        nc164, nc148, nc42, nc231, nc191, nc255, nc283, nc317, 
        nc290, nc17, nc2, nc302, nc110, nc128, nc244, nc321, nc43, 
        nc179, nc157, nc36, nc224, nc296, nc273, nc61, nc104, 
        nc138, nc14, nc285, nc303, nc150, nc331, nc196, nc234, 
        nc149, nc12, nc219, nc30, nc243, nc187, nc65, nc7, nc292, 
        nc129, nc275, nc8, nc223, nc13, nc305, nc180, nc26, nc291, 
        nc177, nc139, nc310, nc259, nc245, nc233, nc163, nc318, 
        nc268, nc112, nc68, nc49, nc314, nc217, nc170, nc91, 
        nc225, nc5, nc20, nc198, nc147, nc316, nc67, nc289, nc294, 
        nc152, nc127, nc103, nc235, nc76, nc208, nc140, nc257, 
        nc86, nc95, nc327, nc120, nc165, nc279, nc137, nc64, nc19, 
        nc312, nc70, nc182, nc62, nc199, nc80, nc130, nc287, nc98, 
        nc293, nc249, nc114, nc56, nc105, nc63, nc313, nc309, 
        nc172, nc229, nc277, nc97, nc161, nc31, nc295, nc154, 
        nc50, nc260, nc239, nc142, nc320, nc315, nc247, nc94, 
        nc197, nc328, nc122, nc266, nc35, nc324, nc4, nc227, nc92, 
        nc101, nc330, nc184, nc200, nc190, nc166, nc326, nc132, 
        nc334, nc21, nc237, nc93, nc262, nc69, nc206, nc174, nc38, 
        nc113, nc218, nc106, nc261, nc25, nc1, nc322, nc299, nc37, 
        nc202, nc144, nc153, nc46, nc258, nc71, nc124, nc332, 
        nc81, nc201, nc168, nc323, nc34, nc28, nc115, nc264, 
        nc192, nc319, nc134, nc32, nc40, nc297, nc99, nc75, nc183, 
        nc333, nc288, nc85, nc27, nc108, nc325, nc16, nc155, nc51, 
        nc301, nc33, nc204, nc173, nc278, nc169, nc78, nc263, 
        nc24, nc88, nc111, nc55, nc10, nc22, nc210, nc185, nc143, 
        nc248, nc77, nc6, nc109, nc87, nc123 : std_logic;

begin 


    MSS_ADLIB_INST_RNO_20 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_520, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_586, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[21]\);
    
    MSS_ADLIB_INST_RNO_40 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_3_21, B => line_4_21, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[28]\, D => 
        result_addr_net_0(1), Y => N_249);
    
    MSS_ADLIB_INST_RNO_23 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_523, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_589, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[24]\);
    
    MSS_ADLIB_INST_RNO_35 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_274, B => N_273, C => line_7_21, D => N_252, 
        Y => \AMBA_SLAVE_0_HRDATA_S0_m_0_0[28]\);
    
    MSS_ADLIB_INST_RNO_43 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_0_d0, B => line_0_0, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[7]\, D => 
        result_addr_net_0(1), Y => N_240);
    
    MSS_ADLIB_INST_RNO_29 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_529, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_595, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[30]\);
    
    MSS_ADLIB_INST_RNO_34 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_274, B => N_273, C => line_7_13, D => N_202, 
        Y => \AMBA_SLAVE_0_HRDATA_S0_m_0_0[20]\);
    
    MSS_ADLIB_INST_RNO_21 : CFG3
      generic map(INIT => x"80")

      port map(A => N_96, B => hready_m_xhdl339, C => ren_pos, Y
         => \AMBA_SLAVE_0_HRDATA_S0_m[22]\);
    
    MSS_ADLIB_INST_RNO_49 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_3, B => line_2_3, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[10]\);
    
    MSS_ADLIB_INST_RNO_41 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_24, B => line_0_24, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[31]\, D => 
        result_addr_net_0(1), Y => N_208);
    
    MSS_ADLIB_INST_RNO : CFG4
      generic map(INIT => x"B080")

      port map(A => N_499, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_565, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[0]\);
    
    MSS_ADLIB_INST_RNO_22 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_522, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_588, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[23]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    MSS_ADLIB_INST_RNO_36 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_3_0, B => line_4_0, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[7]\, D => 
        result_addr_net_0(1), Y => N_237);
    
    MSS_ADLIB_INST_RNO_50 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_4, B => line_2_4, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[11]\);
    
    MSS_ADLIB_INST_RNO_42 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_3_24, B => line_4_24, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[31]\, D => 
        result_addr_net_0(1), Y => N_205);
    
    MSS_ADLIB_INST_RNO_53 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_24, B => line_2_24, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[31]\);
    
    MSS_ADLIB_INST_RNO_27 : CFG3
      generic map(INIT => x"EC")

      port map(A => N_59, B => \AMBA_SLAVE_0_HRDATA_S0_m_0_0[28]\, 
        C => N_249, Y => \AMBA_SLAVE_0_HRDATA_S0_m[28]\);
    
    MSS_ADLIB_INST_RNO_10 : CFG3
      generic map(INIT => x"EC")

      port map(A => N_59, B => \AMBA_SLAVE_0_HRDATA_S0_m_0_0[11]\, 
        C => N_243, Y => \AMBA_SLAVE_0_HRDATA_S0_m[11]\);
    
    MSS_ADLIB_INST_RNO_38 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_4_d0, B => line_0_4, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[11]\, D => 
        result_addr_net_0(1), Y => N_243);
    
    MSS_ADLIB_INST_RNO_59 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_21, B => line_2_21, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[28]\);
    
    MSS_ADLIB_INST_RNO_47 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_21, B => line_0_21, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[28]\, D => 
        result_addr_net_0(1), Y => N_252);
    
    MSS_ADLIB_INST_RNO_13 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_513, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_579, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[14]\);
    
    MSS_ADLIB_INST_RNO_51 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_13, B => line_2_13, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[20]\);
    
    MSS_ADLIB_INST_RNO_19 : CFG3
      generic map(INIT => x"EC")

      port map(A => N_59, B => \AMBA_SLAVE_0_HRDATA_S0_m_0_0[20]\, 
        C => N_199, Y => \AMBA_SLAVE_0_HRDATA_S0_m[20]\);
    
    MSS_ADLIB_INST_RNO_11 : CFG3
      generic map(INIT => x"80")

      port map(A => N_81, B => hready_m_xhdl339, C => ren_pos, Y
         => N_35_i_0);
    
    MSS_ADLIB_INST_RNO_52 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_21, B => line_6_21, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[28]\);
    
    MSS_ADLIB_INST_RNO_12 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_512, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_578, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[13]\);
    
    MSS_ADLIB_INST_RNO_2 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_502, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_568, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[3]\);
    
    MSS_ADLIB_INST_RNO_57 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_4, B => line_6_4, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[11]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    MSS_ADLIB_INST_RNO_4 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_504, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_570, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[5]\);
    
    MSS_ADLIB_INST_RNO_17 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_517, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_583, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[18]\);
    
    MSS_ADLIB_INST_RNO_7 : CFG4
      generic map(INIT => x"C404")

      port map(A => N_7, B => hready_m_xhdl339, C => 
        result_addr_net_0(0), D => N_75, Y => N_25_i_0);
    
    MSS_ADLIB_INST : MSS_060

              generic map(INIT => "00" & x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C000000006092C0104003FFFFE4000000000000100000000F0F15C00000182DFFC010842108421000001FE34001FF8000000400000000020891007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem", RTC_MAIN_XTL_FREQ => 0.0,
         DDR_CLK_FREQ => 100.0)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => OPEN, CAN_TX_EBL_MGPIO4A_H2F_A
         => OPEN, CAN_TX_EBL_MGPIO4A_H2F_B => OPEN, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => OPEN, CLK_CONFIG_APB => OPEN, COMMS_INT => OPEN, 
        CONFIG_PRESET_N => 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        EDAC_ERROR(7) => nc228, EDAC_ERROR(6) => nc203, 
        EDAC_ERROR(5) => nc265, EDAC_ERROR(4) => nc216, 
        EDAC_ERROR(3) => nc194, EDAC_ERROR(2) => nc151, 
        EDAC_ERROR(1) => nc23, EDAC_ERROR(0) => nc175, 
        F_FM0_RDATA(31) => nc250, F_FM0_RDATA(30) => nc58, 
        F_FM0_RDATA(29) => nc116, F_FM0_RDATA(28) => nc74, 
        F_FM0_RDATA(27) => nc133, F_FM0_RDATA(26) => nc238, 
        F_FM0_RDATA(25) => nc167, F_FM0_RDATA(24) => nc84, 
        F_FM0_RDATA(23) => nc39, F_FM0_RDATA(22) => nc72, 
        F_FM0_RDATA(21) => nc256, F_FM0_RDATA(20) => nc212, 
        F_FM0_RDATA(19) => nc205, F_FM0_RDATA(18) => nc82, 
        F_FM0_RDATA(17) => nc145, F_FM0_RDATA(16) => nc181, 
        F_FM0_RDATA(15) => nc160, F_FM0_RDATA(14) => nc57, 
        F_FM0_RDATA(13) => nc156, F_FM0_RDATA(12) => nc280, 
        F_FM0_RDATA(11) => nc125, F_FM0_RDATA(10) => nc211, 
        F_FM0_RDATA(9) => nc73, F_FM0_RDATA(8) => nc107, 
        F_FM0_RDATA(7) => nc329, F_FM0_RDATA(6) => nc66, 
        F_FM0_RDATA(5) => nc83, F_FM0_RDATA(4) => nc9, 
        F_FM0_RDATA(3) => nc252, F_FM0_RDATA(2) => nc171, 
        F_FM0_RDATA(1) => nc54, F_FM0_RDATA(0) => nc286, 
        F_FM0_READYOUT => OPEN, F_FM0_RESP => OPEN, 
        F_HM0_ADDR(31) => nc307, F_HM0_ADDR(30) => nc135, 
        F_HM0_ADDR(29) => nc41, F_HM0_ADDR(28) => nc100, 
        F_HM0_ADDR(27) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_27, 
        F_HM0_ADDR(26) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_26, 
        F_HM0_ADDR(25) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, 
        F_HM0_ADDR(24) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        F_HM0_ADDR(23) => nc270, F_HM0_ADDR(22) => nc52, 
        F_HM0_ADDR(21) => nc251, F_HM0_ADDR(20) => nc186, 
        F_HM0_ADDR(19) => nc29, F_HM0_ADDR(18) => nc269, 
        F_HM0_ADDR(17) => nc118, F_HM0_ADDR(16) => nc60, 
        F_HM0_ADDR(15) => nc141, F_HM0_ADDR(14) => nc311, 
        F_HM0_ADDR(13) => nc276, F_HM0_ADDR(12) => nc193, 
        F_HM0_ADDR(11) => nc214, F_HM0_ADDR(10) => nc298, 
        F_HM0_ADDR(9) => nc282, F_HM0_ADDR(8) => nc240, 
        F_HM0_ADDR(7) => nc45, F_HM0_ADDR(6) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        F_HM0_ADDR(5) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        F_HM0_ADDR(4) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        F_HM0_ADDR(3) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        F_HM0_ADDR(2) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        F_HM0_ADDR(1) => nc53, F_HM0_ADDR(0) => nc121, 
        F_HM0_ENABLE => OPEN, F_HM0_SEL => OPEN, F_HM0_SIZE(1)
         => nc176, F_HM0_SIZE(0) => nc220, F_HM0_TRANS1 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        F_HM0_WDATA(31) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        F_HM0_WDATA(30) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        F_HM0_WDATA(29) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        F_HM0_WDATA(28) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        F_HM0_WDATA(27) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        F_HM0_WDATA(26) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        F_HM0_WDATA(25) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        F_HM0_WDATA(24) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        F_HM0_WDATA(23) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        F_HM0_WDATA(22) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        F_HM0_WDATA(21) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        F_HM0_WDATA(20) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        F_HM0_WDATA(19) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        F_HM0_WDATA(18) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        F_HM0_WDATA(17) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        F_HM0_WDATA(16) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        F_HM0_WDATA(15) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        F_HM0_WDATA(14) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        F_HM0_WDATA(13) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        F_HM0_WDATA(12) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        F_HM0_WDATA(11) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        F_HM0_WDATA(10) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        F_HM0_WDATA(9) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        F_HM0_WDATA(8) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        F_HM0_WDATA(7) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        F_HM0_WDATA(6) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        F_HM0_WDATA(5) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        F_HM0_WDATA(4) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        F_HM0_WDATA(3) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        F_HM0_WDATA(2) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        F_HM0_WDATA(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        F_HM0_WDATA(0) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        F_HM0_WRITE => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        FAB_CHRGVBUS => OPEN, FAB_DISCHRGVBUS => OPEN, 
        FAB_DMPULLDOWN => OPEN, FAB_DPPULLDOWN => OPEN, 
        FAB_DRVVBUS => OPEN, FAB_IDPULLUP => OPEN, FAB_OPMODE(1)
         => nc158, FAB_OPMODE(0) => nc281, FAB_SUSPENDM => OPEN, 
        FAB_TERMSEL => OPEN, FAB_TXVALID => OPEN, FAB_VCONTROL(3)
         => nc209, FAB_VCONTROL(2) => nc246, FAB_VCONTROL(1) => 
        nc162, FAB_VCONTROL(0) => nc11, FAB_VCONTROLLOADM => OPEN, 
        FAB_XCVRSEL(1) => nc272, FAB_XCVRSEL(0) => nc131, 
        FAB_XDATAOUT(7) => nc254, FAB_XDATAOUT(6) => nc267, 
        FAB_XDATAOUT(5) => nc96, FAB_XDATAOUT(4) => nc79, 
        FAB_XDATAOUT(3) => nc226, FAB_XDATAOUT(2) => nc146, 
        FAB_XDATAOUT(1) => nc230, FAB_XDATAOUT(0) => nc89, 
        FACC_GLMUX_SEL => OPEN, FIC32_0_MASTER(1) => nc119, 
        FIC32_0_MASTER(0) => nc48, FIC32_1_MASTER(1) => nc271, 
        FIC32_1_MASTER(0) => nc213, FPGA_RESET_N => 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, GTX_CLK => 
        OPEN, H2F_INTERRUPT(15) => nc300, H2F_INTERRUPT(14) => 
        nc126, H2F_INTERRUPT(13) => nc195, H2F_INTERRUPT(12) => 
        nc188, H2F_INTERRUPT(11) => nc242, H2F_INTERRUPT(10) => 
        nc15, H2F_INTERRUPT(9) => nc308, H2F_INTERRUPT(8) => 
        nc236, H2F_INTERRUPT(7) => nc102, H2F_INTERRUPT(6) => 
        nc304, H2F_INTERRUPT(5) => nc3, H2F_INTERRUPT(4) => nc207, 
        H2F_INTERRUPT(3) => nc47, H2F_INTERRUPT(2) => nc90, 
        H2F_INTERRUPT(1) => nc284, H2F_INTERRUPT(0) => nc222, 
        H2F_NMI => OPEN, H2FCALIB => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_A => OPEN, I2C0_SCL_MGPIO31B_H2F_B
         => OPEN, I2C0_SDA_MGPIO30B_H2F_A => OPEN, 
        I2C0_SDA_MGPIO30B_H2F_B => OPEN, I2C1_SCL_MGPIO1A_H2F_A
         => OPEN, I2C1_SCL_MGPIO1A_H2F_B => 
        sha256_system_sb_0_GPIO_1_M2F, I2C1_SDA_MGPIO0A_H2F_A => 
        OPEN, I2C1_SDA_MGPIO0A_H2F_B => GPIO_0_M2F_c, MDCF => 
        OPEN, MDOENF => OPEN, MDOF => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_A => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => OPEN, MPLL_LOCK => OPEN, 
        PER2_FABRIC_PADDR(15) => nc159, PER2_FABRIC_PADDR(14) => 
        nc136, PER2_FABRIC_PADDR(13) => nc241, 
        PER2_FABRIC_PADDR(12) => nc253, PER2_FABRIC_PADDR(11) => 
        nc178, PER2_FABRIC_PADDR(10) => nc306, 
        PER2_FABRIC_PADDR(9) => nc215, PER2_FABRIC_PADDR(8) => 
        nc59, PER2_FABRIC_PADDR(7) => nc221, PER2_FABRIC_PADDR(6)
         => nc232, PER2_FABRIC_PADDR(5) => nc274, 
        PER2_FABRIC_PADDR(4) => nc18, PER2_FABRIC_PADDR(3) => 
        nc44, PER2_FABRIC_PADDR(2) => nc117, PER2_FABRIC_PENABLE
         => OPEN, PER2_FABRIC_PSEL => OPEN, 
        PER2_FABRIC_PWDATA(31) => nc189, PER2_FABRIC_PWDATA(30)
         => nc164, PER2_FABRIC_PWDATA(29) => nc148, 
        PER2_FABRIC_PWDATA(28) => nc42, PER2_FABRIC_PWDATA(27)
         => nc231, PER2_FABRIC_PWDATA(26) => nc191, 
        PER2_FABRIC_PWDATA(25) => nc255, PER2_FABRIC_PWDATA(24)
         => nc283, PER2_FABRIC_PWDATA(23) => nc317, 
        PER2_FABRIC_PWDATA(22) => nc290, PER2_FABRIC_PWDATA(21)
         => nc17, PER2_FABRIC_PWDATA(20) => nc2, 
        PER2_FABRIC_PWDATA(19) => nc302, PER2_FABRIC_PWDATA(18)
         => nc110, PER2_FABRIC_PWDATA(17) => nc128, 
        PER2_FABRIC_PWDATA(16) => nc244, PER2_FABRIC_PWDATA(15)
         => nc321, PER2_FABRIC_PWDATA(14) => nc43, 
        PER2_FABRIC_PWDATA(13) => nc179, PER2_FABRIC_PWDATA(12)
         => nc157, PER2_FABRIC_PWDATA(11) => nc36, 
        PER2_FABRIC_PWDATA(10) => nc224, PER2_FABRIC_PWDATA(9)
         => nc296, PER2_FABRIC_PWDATA(8) => nc273, 
        PER2_FABRIC_PWDATA(7) => nc61, PER2_FABRIC_PWDATA(6) => 
        nc104, PER2_FABRIC_PWDATA(5) => nc138, 
        PER2_FABRIC_PWDATA(4) => nc14, PER2_FABRIC_PWDATA(3) => 
        nc285, PER2_FABRIC_PWDATA(2) => nc303, 
        PER2_FABRIC_PWDATA(1) => nc150, PER2_FABRIC_PWDATA(0) => 
        nc331, PER2_FABRIC_PWRITE => OPEN, RTC_MATCH => OPEN, 
        SLEEPDEEP => OPEN, SLEEPHOLDACK => OPEN, SLEEPING => OPEN, 
        SMBALERT_NO0 => OPEN, SMBALERT_NO1 => OPEN, SMBSUS_NO0
         => OPEN, SMBSUS_NO1 => OPEN, SPI0_CLK_OUT => OPEN, 
        SPI0_SDI_MGPIO5A_H2F_A => OPEN, SPI0_SDI_MGPIO5A_H2F_B
         => OPEN, SPI0_SDO_MGPIO6A_H2F_A => OPEN, 
        SPI0_SDO_MGPIO6A_H2F_B => OPEN, SPI0_SS0_MGPIO7A_H2F_A
         => OPEN, SPI0_SS0_MGPIO7A_H2F_B => OPEN, 
        SPI0_SS1_MGPIO8A_H2F_A => OPEN, SPI0_SS1_MGPIO8A_H2F_B
         => OPEN, SPI0_SS2_MGPIO9A_H2F_A => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_B => sha256_system_sb_0_GPIO_9_M2F, 
        SPI0_SS3_MGPIO10A_H2F_A => OPEN, SPI0_SS3_MGPIO10A_H2F_B
         => OPEN, SPI0_SS4_MGPIO19A_H2F_A => OPEN, 
        SPI0_SS5_MGPIO20A_H2F_A => OPEN, SPI0_SS6_MGPIO21A_H2F_A
         => OPEN, SPI0_SS7_MGPIO22A_H2F_A => OPEN, SPI1_CLK_OUT
         => OPEN, SPI1_SDI_MGPIO11A_H2F_A => OPEN, 
        SPI1_SDI_MGPIO11A_H2F_B => OPEN, SPI1_SDO_MGPIO12A_H2F_A
         => OPEN, SPI1_SDO_MGPIO12A_H2F_B => OPEN, 
        SPI1_SS0_MGPIO13A_H2F_A => OPEN, SPI1_SS0_MGPIO13A_H2F_B
         => OPEN, SPI1_SS1_MGPIO14A_H2F_A => OPEN, 
        SPI1_SS1_MGPIO14A_H2F_B => OPEN, SPI1_SS2_MGPIO15A_H2F_A
         => OPEN, SPI1_SS2_MGPIO15A_H2F_B => OPEN, 
        SPI1_SS3_MGPIO16A_H2F_A => OPEN, SPI1_SS3_MGPIO16A_H2F_B
         => OPEN, SPI1_SS4_MGPIO17A_H2F_A => OPEN, 
        SPI1_SS5_MGPIO18A_H2F_A => OPEN, SPI1_SS6_MGPIO23A_H2F_A
         => OPEN, SPI1_SS7_MGPIO24A_H2F_A => OPEN, TCGF(9) => 
        nc196, TCGF(8) => nc234, TCGF(7) => nc149, TCGF(6) => 
        nc12, TCGF(5) => nc219, TCGF(4) => nc30, TCGF(3) => nc243, 
        TCGF(2) => nc187, TCGF(1) => nc65, TCGF(0) => nc7, 
        TRACECLK => OPEN, TRACEDATA(3) => nc292, TRACEDATA(2) => 
        nc129, TRACEDATA(1) => nc275, TRACEDATA(0) => nc8, TX_CLK
         => OPEN, TX_ENF => OPEN, TX_ERRF => OPEN, TXCTL_EN_RIF
         => OPEN, TXD_RIF(3) => nc223, TXD_RIF(2) => nc13, 
        TXD_RIF(1) => nc305, TXD_RIF(0) => nc180, TXDF(7) => nc26, 
        TXDF(6) => nc291, TXDF(5) => nc177, TXDF(4) => nc139, 
        TXDF(3) => nc310, TXDF(2) => nc259, TXDF(1) => nc245, 
        TXDF(0) => nc233, TXEV => OPEN, WDOGTIMEOUT => OPEN, 
        F_ARREADY_HREADYOUT1 => OPEN, F_AWREADY_HREADYOUT0 => 
        OPEN, F_BID(3) => nc163, F_BID(2) => nc318, F_BID(1) => 
        nc268, F_BID(0) => nc112, F_BRESP_HRESP0(1) => nc68, 
        F_BRESP_HRESP0(0) => nc49, F_BVALID => OPEN, 
        F_RDATA_HRDATA01(63) => nc314, F_RDATA_HRDATA01(62) => 
        nc217, F_RDATA_HRDATA01(61) => nc170, 
        F_RDATA_HRDATA01(60) => nc91, F_RDATA_HRDATA01(59) => 
        nc225, F_RDATA_HRDATA01(58) => nc5, F_RDATA_HRDATA01(57)
         => nc20, F_RDATA_HRDATA01(56) => nc198, 
        F_RDATA_HRDATA01(55) => nc147, F_RDATA_HRDATA01(54) => 
        nc316, F_RDATA_HRDATA01(53) => nc67, F_RDATA_HRDATA01(52)
         => nc289, F_RDATA_HRDATA01(51) => nc294, 
        F_RDATA_HRDATA01(50) => nc152, F_RDATA_HRDATA01(49) => 
        nc127, F_RDATA_HRDATA01(48) => nc103, 
        F_RDATA_HRDATA01(47) => nc235, F_RDATA_HRDATA01(46) => 
        nc76, F_RDATA_HRDATA01(45) => nc208, F_RDATA_HRDATA01(44)
         => nc140, F_RDATA_HRDATA01(43) => nc257, 
        F_RDATA_HRDATA01(42) => nc86, F_RDATA_HRDATA01(41) => 
        nc95, F_RDATA_HRDATA01(40) => nc327, F_RDATA_HRDATA01(39)
         => nc120, F_RDATA_HRDATA01(38) => nc165, 
        F_RDATA_HRDATA01(37) => nc279, F_RDATA_HRDATA01(36) => 
        nc137, F_RDATA_HRDATA01(35) => nc64, F_RDATA_HRDATA01(34)
         => nc19, F_RDATA_HRDATA01(33) => nc312, 
        F_RDATA_HRDATA01(32) => nc70, F_RDATA_HRDATA01(31) => 
        nc182, F_RDATA_HRDATA01(30) => nc62, F_RDATA_HRDATA01(29)
         => nc199, F_RDATA_HRDATA01(28) => nc80, 
        F_RDATA_HRDATA01(27) => nc130, F_RDATA_HRDATA01(26) => 
        nc287, F_RDATA_HRDATA01(25) => nc98, F_RDATA_HRDATA01(24)
         => nc293, F_RDATA_HRDATA01(23) => nc249, 
        F_RDATA_HRDATA01(22) => nc114, F_RDATA_HRDATA01(21) => 
        nc56, F_RDATA_HRDATA01(20) => nc105, F_RDATA_HRDATA01(19)
         => nc63, F_RDATA_HRDATA01(18) => nc313, 
        F_RDATA_HRDATA01(17) => nc309, F_RDATA_HRDATA01(16) => 
        nc172, F_RDATA_HRDATA01(15) => nc229, 
        F_RDATA_HRDATA01(14) => nc277, F_RDATA_HRDATA01(13) => 
        nc97, F_RDATA_HRDATA01(12) => nc161, F_RDATA_HRDATA01(11)
         => nc31, F_RDATA_HRDATA01(10) => nc295, 
        F_RDATA_HRDATA01(9) => nc154, F_RDATA_HRDATA01(8) => nc50, 
        F_RDATA_HRDATA01(7) => nc260, F_RDATA_HRDATA01(6) => 
        nc239, F_RDATA_HRDATA01(5) => nc142, F_RDATA_HRDATA01(4)
         => nc320, F_RDATA_HRDATA01(3) => nc315, 
        F_RDATA_HRDATA01(2) => nc247, F_RDATA_HRDATA01(1) => nc94, 
        F_RDATA_HRDATA01(0) => nc197, F_RID(3) => nc328, F_RID(2)
         => nc122, F_RID(1) => nc266, F_RID(0) => nc35, F_RLAST
         => OPEN, F_RRESP_HRESP1(1) => nc324, F_RRESP_HRESP1(0)
         => nc4, F_RVALID => OPEN, F_WREADY => OPEN, 
        MDDR_FABRIC_PRDATA(15) => nc227, MDDR_FABRIC_PRDATA(14)
         => nc92, MDDR_FABRIC_PRDATA(13) => nc101, 
        MDDR_FABRIC_PRDATA(12) => nc330, MDDR_FABRIC_PRDATA(11)
         => nc184, MDDR_FABRIC_PRDATA(10) => nc200, 
        MDDR_FABRIC_PRDATA(9) => nc190, MDDR_FABRIC_PRDATA(8) => 
        nc166, MDDR_FABRIC_PRDATA(7) => nc326, 
        MDDR_FABRIC_PRDATA(6) => nc132, MDDR_FABRIC_PRDATA(5) => 
        nc334, MDDR_FABRIC_PRDATA(4) => nc21, 
        MDDR_FABRIC_PRDATA(3) => nc237, MDDR_FABRIC_PRDATA(2) => 
        nc93, MDDR_FABRIC_PRDATA(1) => nc262, 
        MDDR_FABRIC_PRDATA(0) => nc69, MDDR_FABRIC_PREADY => OPEN, 
        MDDR_FABRIC_PSLVERR => OPEN, CAN_RXBUS_F2H_SCP => 
        VCC_net_1, CAN_TX_EBL_F2H_SCP => VCC_net_1, 
        CAN_TXBUS_F2H_SCP => VCC_net_1, COLF => VCC_net_1, CRSF
         => VCC_net_1, F2_DMAREADY(1) => VCC_net_1, 
        F2_DMAREADY(0) => VCC_net_1, F2H_INTERRUPT(15) => 
        GND_net_1, F2H_INTERRUPT(14) => GND_net_1, 
        F2H_INTERRUPT(13) => GND_net_1, F2H_INTERRUPT(12) => 
        GND_net_1, F2H_INTERRUPT(11) => GND_net_1, 
        F2H_INTERRUPT(10) => GND_net_1, F2H_INTERRUPT(9) => 
        GND_net_1, F2H_INTERRUPT(8) => GND_net_1, 
        F2H_INTERRUPT(7) => GND_net_1, F2H_INTERRUPT(6) => 
        GND_net_1, F2H_INTERRUPT(5) => GND_net_1, 
        F2H_INTERRUPT(4) => GND_net_1, F2H_INTERRUPT(3) => 
        GND_net_1, F2H_INTERRUPT(2) => GND_net_1, 
        F2H_INTERRUPT(1) => GND_net_1, F2H_INTERRUPT(0) => 
        GND_net_1, F2HCALIB => VCC_net_1, F_DMAREADY(1) => 
        VCC_net_1, F_DMAREADY(0) => VCC_net_1, F_FM0_ADDR(31) => 
        GND_net_1, F_FM0_ADDR(30) => GND_net_1, F_FM0_ADDR(29)
         => GND_net_1, F_FM0_ADDR(28) => GND_net_1, 
        F_FM0_ADDR(27) => GND_net_1, F_FM0_ADDR(26) => GND_net_1, 
        F_FM0_ADDR(25) => GND_net_1, F_FM0_ADDR(24) => GND_net_1, 
        F_FM0_ADDR(23) => GND_net_1, F_FM0_ADDR(22) => GND_net_1, 
        F_FM0_ADDR(21) => GND_net_1, F_FM0_ADDR(20) => GND_net_1, 
        F_FM0_ADDR(19) => GND_net_1, F_FM0_ADDR(18) => GND_net_1, 
        F_FM0_ADDR(17) => GND_net_1, F_FM0_ADDR(16) => GND_net_1, 
        F_FM0_ADDR(15) => GND_net_1, F_FM0_ADDR(14) => GND_net_1, 
        F_FM0_ADDR(13) => GND_net_1, F_FM0_ADDR(12) => GND_net_1, 
        F_FM0_ADDR(11) => GND_net_1, F_FM0_ADDR(10) => GND_net_1, 
        F_FM0_ADDR(9) => GND_net_1, F_FM0_ADDR(8) => GND_net_1, 
        F_FM0_ADDR(7) => GND_net_1, F_FM0_ADDR(6) => GND_net_1, 
        F_FM0_ADDR(5) => GND_net_1, F_FM0_ADDR(4) => GND_net_1, 
        F_FM0_ADDR(3) => GND_net_1, F_FM0_ADDR(2) => GND_net_1, 
        F_FM0_ADDR(1) => GND_net_1, F_FM0_ADDR(0) => GND_net_1, 
        F_FM0_ENABLE => GND_net_1, F_FM0_MASTLOCK => GND_net_1, 
        F_FM0_READY => VCC_net_1, F_FM0_SEL => GND_net_1, 
        F_FM0_SIZE(1) => GND_net_1, F_FM0_SIZE(0) => GND_net_1, 
        F_FM0_TRANS1 => GND_net_1, F_FM0_WDATA(31) => GND_net_1, 
        F_FM0_WDATA(30) => GND_net_1, F_FM0_WDATA(29) => 
        GND_net_1, F_FM0_WDATA(28) => GND_net_1, F_FM0_WDATA(27)
         => GND_net_1, F_FM0_WDATA(26) => GND_net_1, 
        F_FM0_WDATA(25) => GND_net_1, F_FM0_WDATA(24) => 
        GND_net_1, F_FM0_WDATA(23) => GND_net_1, F_FM0_WDATA(22)
         => GND_net_1, F_FM0_WDATA(21) => GND_net_1, 
        F_FM0_WDATA(20) => GND_net_1, F_FM0_WDATA(19) => 
        GND_net_1, F_FM0_WDATA(18) => GND_net_1, F_FM0_WDATA(17)
         => GND_net_1, F_FM0_WDATA(16) => GND_net_1, 
        F_FM0_WDATA(15) => GND_net_1, F_FM0_WDATA(14) => 
        GND_net_1, F_FM0_WDATA(13) => GND_net_1, F_FM0_WDATA(12)
         => GND_net_1, F_FM0_WDATA(11) => GND_net_1, 
        F_FM0_WDATA(10) => GND_net_1, F_FM0_WDATA(9) => GND_net_1, 
        F_FM0_WDATA(8) => GND_net_1, F_FM0_WDATA(7) => GND_net_1, 
        F_FM0_WDATA(6) => GND_net_1, F_FM0_WDATA(5) => GND_net_1, 
        F_FM0_WDATA(4) => GND_net_1, F_FM0_WDATA(3) => GND_net_1, 
        F_FM0_WDATA(2) => GND_net_1, F_FM0_WDATA(1) => GND_net_1, 
        F_FM0_WDATA(0) => GND_net_1, F_FM0_WRITE => GND_net_1, 
        F_HM0_RDATA(31) => \AMBA_SLAVE_0_HRDATA_S0_m[31]\, 
        F_HM0_RDATA(30) => \AMBA_SLAVE_0_HRDATA_S0_m[30]\, 
        F_HM0_RDATA(29) => \AMBA_SLAVE_0_HRDATA_S0_m[29]\, 
        F_HM0_RDATA(28) => \AMBA_SLAVE_0_HRDATA_S0_m[28]\, 
        F_HM0_RDATA(27) => \AMBA_SLAVE_0_HRDATA_S0_m[27]\, 
        F_HM0_RDATA(26) => \AMBA_SLAVE_0_HRDATA_S0_m[26]\, 
        F_HM0_RDATA(25) => \AMBA_SLAVE_0_HRDATA_S0_m[25]\, 
        F_HM0_RDATA(24) => \AMBA_SLAVE_0_HRDATA_S0_m[24]\, 
        F_HM0_RDATA(23) => \AMBA_SLAVE_0_HRDATA_S0_m[23]\, 
        F_HM0_RDATA(22) => \AMBA_SLAVE_0_HRDATA_S0_m[22]\, 
        F_HM0_RDATA(21) => \AMBA_SLAVE_0_HRDATA_S0_m[21]\, 
        F_HM0_RDATA(20) => \AMBA_SLAVE_0_HRDATA_S0_m[20]\, 
        F_HM0_RDATA(19) => N_34_i_0, F_HM0_RDATA(18) => 
        \AMBA_SLAVE_0_HRDATA_S0_m[18]\, F_HM0_RDATA(17) => 
        \AMBA_SLAVE_0_HRDATA_S0_m[17]\, F_HM0_RDATA(16) => 
        \AMBA_SLAVE_0_HRDATA_S0_m[16]\, F_HM0_RDATA(15) => 
        \AMBA_SLAVE_0_HRDATA_S0_m[15]\, F_HM0_RDATA(14) => 
        \AMBA_SLAVE_0_HRDATA_S0_m[14]\, F_HM0_RDATA(13) => 
        \AMBA_SLAVE_0_HRDATA_S0_m[13]\, F_HM0_RDATA(12) => 
        N_35_i_0, F_HM0_RDATA(11) => 
        \AMBA_SLAVE_0_HRDATA_S0_m[11]\, F_HM0_RDATA(10) => 
        \AMBA_SLAVE_0_HRDATA_S0_m[10]\, F_HM0_RDATA(9) => 
        \AMBA_SLAVE_0_HRDATA_S0_m[9]\, F_HM0_RDATA(8) => N_25_i_0, 
        F_HM0_RDATA(7) => \AMBA_SLAVE_0_HRDATA_S0_m[7]\, 
        F_HM0_RDATA(6) => \AMBA_SLAVE_0_HRDATA_S0_m[6]\, 
        F_HM0_RDATA(5) => \AMBA_SLAVE_0_HRDATA_S0_m[5]\, 
        F_HM0_RDATA(4) => \AMBA_SLAVE_0_HRDATA_S0_m[4]\, 
        F_HM0_RDATA(3) => \AMBA_SLAVE_0_HRDATA_S0_m[3]\, 
        F_HM0_RDATA(2) => \AMBA_SLAVE_0_HRDATA_S0_m[2]\, 
        F_HM0_RDATA(1) => \AMBA_SLAVE_0_HRDATA_S0_m[1]\, 
        F_HM0_RDATA(0) => \AMBA_SLAVE_0_HRDATA_S0_m[0]\, 
        F_HM0_READY => N_23_i_0, F_HM0_RESP => N_31, FAB_AVALID
         => VCC_net_1, FAB_HOSTDISCON => VCC_net_1, FAB_IDDIG => 
        VCC_net_1, FAB_LINESTATE(1) => VCC_net_1, 
        FAB_LINESTATE(0) => VCC_net_1, FAB_M3_RESET_N => 
        VCC_net_1, FAB_PLL_LOCK => FIC_0_LOCK, FAB_RXACTIVE => 
        VCC_net_1, FAB_RXERROR => VCC_net_1, FAB_RXVALID => 
        VCC_net_1, FAB_RXVALIDH => GND_net_1, FAB_SESSEND => 
        VCC_net_1, FAB_TXREADY => VCC_net_1, FAB_VBUSVALID => 
        VCC_net_1, FAB_VSTATUS(7) => VCC_net_1, FAB_VSTATUS(6)
         => VCC_net_1, FAB_VSTATUS(5) => VCC_net_1, 
        FAB_VSTATUS(4) => VCC_net_1, FAB_VSTATUS(3) => VCC_net_1, 
        FAB_VSTATUS(2) => VCC_net_1, FAB_VSTATUS(1) => VCC_net_1, 
        FAB_VSTATUS(0) => VCC_net_1, FAB_XDATAIN(7) => VCC_net_1, 
        FAB_XDATAIN(6) => VCC_net_1, FAB_XDATAIN(5) => VCC_net_1, 
        FAB_XDATAIN(4) => VCC_net_1, FAB_XDATAIN(3) => VCC_net_1, 
        FAB_XDATAIN(2) => VCC_net_1, FAB_XDATAIN(1) => VCC_net_1, 
        FAB_XDATAIN(0) => VCC_net_1, GTX_CLKPF => VCC_net_1, 
        I2C0_BCLK => VCC_net_1, I2C0_SCL_F2H_SCP => VCC_net_1, 
        I2C0_SDA_F2H_SCP => VCC_net_1, I2C1_BCLK => VCC_net_1, 
        I2C1_SCL_F2H_SCP => VCC_net_1, I2C1_SDA_F2H_SCP => 
        VCC_net_1, MDIF => VCC_net_1, MGPIO0A_F2H_GPIN => 
        VCC_net_1, MGPIO10A_F2H_GPIN => state_out_net_0(0), 
        MGPIO11A_F2H_GPIN => N_87_i_0, MGPIO11B_F2H_GPIN => 
        VCC_net_1, MGPIO12A_F2H_GPIN => N_88_i_0, 
        MGPIO13A_F2H_GPIN => VCC_net_1, MGPIO14A_F2H_GPIN => 
        VCC_net_1, MGPIO15A_F2H_GPIN => VCC_net_1, 
        MGPIO16A_F2H_GPIN => VCC_net_1, MGPIO17B_F2H_GPIN => 
        VCC_net_1, MGPIO18B_F2H_GPIN => VCC_net_1, 
        MGPIO19B_F2H_GPIN => VCC_net_1, MGPIO1A_F2H_GPIN => 
        VCC_net_1, MGPIO20B_F2H_GPIN => VCC_net_1, 
        MGPIO21B_F2H_GPIN => VCC_net_1, MGPIO22B_F2H_GPIN => 
        VCC_net_1, MGPIO24B_F2H_GPIN => VCC_net_1, 
        MGPIO25B_F2H_GPIN => VCC_net_1, MGPIO26B_F2H_GPIN => 
        VCC_net_1, MGPIO27B_F2H_GPIN => VCC_net_1, 
        MGPIO28B_F2H_GPIN => VCC_net_1, MGPIO29B_F2H_GPIN => 
        VCC_net_1, MGPIO2A_F2H_GPIN => ce_i_i_2_i_0, 
        MGPIO30B_F2H_GPIN => VCC_net_1, MGPIO31B_F2H_GPIN => 
        VCC_net_1, MGPIO3A_F2H_GPIN => 
        SHA256_Module_0_data_available_lastbank_8, 
        MGPIO4A_F2H_GPIN => SHA256_Module_0_di_req_o, 
        MGPIO5A_F2H_GPIN => SHA256_Module_0_data_out_ready, 
        MGPIO6A_F2H_GPIN => SHA256_Module_0_do_valid_o, 
        MGPIO7A_F2H_GPIN => SHA256_Module_0_data_available, 
        MGPIO8A_F2H_GPIN => SHA256_Module_0_error_o, 
        MGPIO9A_F2H_GPIN => VCC_net_1, MMUART0_CTS_F2H_SCP => 
        VCC_net_1, MMUART0_DCD_F2H_SCP => VCC_net_1, 
        MMUART0_DSR_F2H_SCP => VCC_net_1, MMUART0_DTR_F2H_SCP => 
        VCC_net_1, MMUART0_RI_F2H_SCP => VCC_net_1, 
        MMUART0_RTS_F2H_SCP => VCC_net_1, MMUART0_RXD_F2H_SCP => 
        VCC_net_1, MMUART0_SCK_F2H_SCP => VCC_net_1, 
        MMUART0_TXD_F2H_SCP => VCC_net_1, MMUART1_CTS_F2H_SCP => 
        VCC_net_1, MMUART1_DCD_F2H_SCP => VCC_net_1, 
        MMUART1_DSR_F2H_SCP => VCC_net_1, MMUART1_RI_F2H_SCP => 
        VCC_net_1, MMUART1_RTS_F2H_SCP => VCC_net_1, 
        MMUART1_RXD_F2H_SCP => VCC_net_1, MMUART1_SCK_F2H_SCP => 
        VCC_net_1, MMUART1_TXD_F2H_SCP => VCC_net_1, 
        PER2_FABRIC_PRDATA(31) => GND_net_1, 
        PER2_FABRIC_PRDATA(30) => GND_net_1, 
        PER2_FABRIC_PRDATA(29) => GND_net_1, 
        PER2_FABRIC_PRDATA(28) => GND_net_1, 
        PER2_FABRIC_PRDATA(27) => GND_net_1, 
        PER2_FABRIC_PRDATA(26) => GND_net_1, 
        PER2_FABRIC_PRDATA(25) => GND_net_1, 
        PER2_FABRIC_PRDATA(24) => GND_net_1, 
        PER2_FABRIC_PRDATA(23) => GND_net_1, 
        PER2_FABRIC_PRDATA(22) => GND_net_1, 
        PER2_FABRIC_PRDATA(21) => GND_net_1, 
        PER2_FABRIC_PRDATA(20) => GND_net_1, 
        PER2_FABRIC_PRDATA(19) => GND_net_1, 
        PER2_FABRIC_PRDATA(18) => GND_net_1, 
        PER2_FABRIC_PRDATA(17) => GND_net_1, 
        PER2_FABRIC_PRDATA(16) => GND_net_1, 
        PER2_FABRIC_PRDATA(15) => GND_net_1, 
        PER2_FABRIC_PRDATA(14) => GND_net_1, 
        PER2_FABRIC_PRDATA(13) => GND_net_1, 
        PER2_FABRIC_PRDATA(12) => GND_net_1, 
        PER2_FABRIC_PRDATA(11) => GND_net_1, 
        PER2_FABRIC_PRDATA(10) => GND_net_1, 
        PER2_FABRIC_PRDATA(9) => GND_net_1, PER2_FABRIC_PRDATA(8)
         => GND_net_1, PER2_FABRIC_PRDATA(7) => GND_net_1, 
        PER2_FABRIC_PRDATA(6) => GND_net_1, PER2_FABRIC_PRDATA(5)
         => GND_net_1, PER2_FABRIC_PRDATA(4) => GND_net_1, 
        PER2_FABRIC_PRDATA(3) => GND_net_1, PER2_FABRIC_PRDATA(2)
         => GND_net_1, PER2_FABRIC_PRDATA(1) => GND_net_1, 
        PER2_FABRIC_PRDATA(0) => GND_net_1, PER2_FABRIC_PREADY
         => VCC_net_1, PER2_FABRIC_PSLVERR => GND_net_1, RCGF(9)
         => VCC_net_1, RCGF(8) => VCC_net_1, RCGF(7) => VCC_net_1, 
        RCGF(6) => VCC_net_1, RCGF(5) => VCC_net_1, RCGF(4) => 
        VCC_net_1, RCGF(3) => VCC_net_1, RCGF(2) => VCC_net_1, 
        RCGF(1) => VCC_net_1, RCGF(0) => VCC_net_1, RX_CLKPF => 
        VCC_net_1, RX_DVF => VCC_net_1, RX_ERRF => VCC_net_1, 
        RX_EV => VCC_net_1, RXDF(7) => VCC_net_1, RXDF(6) => 
        VCC_net_1, RXDF(5) => VCC_net_1, RXDF(4) => VCC_net_1, 
        RXDF(3) => VCC_net_1, RXDF(2) => VCC_net_1, RXDF(1) => 
        VCC_net_1, RXDF(0) => VCC_net_1, SLEEPHOLDREQ => 
        GND_net_1, SMBALERT_NI0 => VCC_net_1, SMBALERT_NI1 => 
        VCC_net_1, SMBSUS_NI0 => VCC_net_1, SMBSUS_NI1 => 
        VCC_net_1, SPI0_CLK_IN => VCC_net_1, SPI0_SDI_F2H_SCP => 
        VCC_net_1, SPI0_SDO_F2H_SCP => VCC_net_1, 
        SPI0_SS0_F2H_SCP => VCC_net_1, SPI0_SS1_F2H_SCP => 
        VCC_net_1, SPI0_SS2_F2H_SCP => VCC_net_1, 
        SPI0_SS3_F2H_SCP => VCC_net_1, SPI1_CLK_IN => VCC_net_1, 
        SPI1_SDI_F2H_SCP => VCC_net_1, SPI1_SDO_F2H_SCP => 
        VCC_net_1, SPI1_SS0_F2H_SCP => VCC_net_1, 
        SPI1_SS1_F2H_SCP => VCC_net_1, SPI1_SS2_F2H_SCP => 
        VCC_net_1, SPI1_SS3_F2H_SCP => VCC_net_1, TX_CLKPF => 
        VCC_net_1, USER_MSS_GPIO_RESET_N => VCC_net_1, 
        USER_MSS_RESET_N => VCC_net_1, XCLK_FAB => VCC_net_1, 
        CLK_BASE => sha256_system_sb_0_FIC_0_CLK, CLK_MDDR_APB
         => VCC_net_1, F_ARADDR_HADDR1(31) => VCC_net_1, 
        F_ARADDR_HADDR1(30) => VCC_net_1, F_ARADDR_HADDR1(29) => 
        VCC_net_1, F_ARADDR_HADDR1(28) => VCC_net_1, 
        F_ARADDR_HADDR1(27) => VCC_net_1, F_ARADDR_HADDR1(26) => 
        VCC_net_1, F_ARADDR_HADDR1(25) => VCC_net_1, 
        F_ARADDR_HADDR1(24) => VCC_net_1, F_ARADDR_HADDR1(23) => 
        VCC_net_1, F_ARADDR_HADDR1(22) => VCC_net_1, 
        F_ARADDR_HADDR1(21) => VCC_net_1, F_ARADDR_HADDR1(20) => 
        VCC_net_1, F_ARADDR_HADDR1(19) => VCC_net_1, 
        F_ARADDR_HADDR1(18) => VCC_net_1, F_ARADDR_HADDR1(17) => 
        VCC_net_1, F_ARADDR_HADDR1(16) => VCC_net_1, 
        F_ARADDR_HADDR1(15) => VCC_net_1, F_ARADDR_HADDR1(14) => 
        VCC_net_1, F_ARADDR_HADDR1(13) => VCC_net_1, 
        F_ARADDR_HADDR1(12) => VCC_net_1, F_ARADDR_HADDR1(11) => 
        VCC_net_1, F_ARADDR_HADDR1(10) => VCC_net_1, 
        F_ARADDR_HADDR1(9) => VCC_net_1, F_ARADDR_HADDR1(8) => 
        VCC_net_1, F_ARADDR_HADDR1(7) => VCC_net_1, 
        F_ARADDR_HADDR1(6) => VCC_net_1, F_ARADDR_HADDR1(5) => 
        VCC_net_1, F_ARADDR_HADDR1(4) => VCC_net_1, 
        F_ARADDR_HADDR1(3) => VCC_net_1, F_ARADDR_HADDR1(2) => 
        VCC_net_1, F_ARADDR_HADDR1(1) => VCC_net_1, 
        F_ARADDR_HADDR1(0) => VCC_net_1, F_ARBURST_HTRANS1(1) => 
        GND_net_1, F_ARBURST_HTRANS1(0) => GND_net_1, 
        F_ARID_HSEL1(3) => GND_net_1, F_ARID_HSEL1(2) => 
        GND_net_1, F_ARID_HSEL1(1) => GND_net_1, F_ARID_HSEL1(0)
         => GND_net_1, F_ARLEN_HBURST1(3) => GND_net_1, 
        F_ARLEN_HBURST1(2) => GND_net_1, F_ARLEN_HBURST1(1) => 
        GND_net_1, F_ARLEN_HBURST1(0) => GND_net_1, 
        F_ARLOCK_HMASTLOCK1(1) => GND_net_1, 
        F_ARLOCK_HMASTLOCK1(0) => GND_net_1, F_ARSIZE_HSIZE1(1)
         => GND_net_1, F_ARSIZE_HSIZE1(0) => GND_net_1, 
        F_ARVALID_HWRITE1 => GND_net_1, F_AWADDR_HADDR0(31) => 
        VCC_net_1, F_AWADDR_HADDR0(30) => VCC_net_1, 
        F_AWADDR_HADDR0(29) => VCC_net_1, F_AWADDR_HADDR0(28) => 
        VCC_net_1, F_AWADDR_HADDR0(27) => VCC_net_1, 
        F_AWADDR_HADDR0(26) => VCC_net_1, F_AWADDR_HADDR0(25) => 
        VCC_net_1, F_AWADDR_HADDR0(24) => VCC_net_1, 
        F_AWADDR_HADDR0(23) => VCC_net_1, F_AWADDR_HADDR0(22) => 
        VCC_net_1, F_AWADDR_HADDR0(21) => VCC_net_1, 
        F_AWADDR_HADDR0(20) => VCC_net_1, F_AWADDR_HADDR0(19) => 
        VCC_net_1, F_AWADDR_HADDR0(18) => VCC_net_1, 
        F_AWADDR_HADDR0(17) => VCC_net_1, F_AWADDR_HADDR0(16) => 
        VCC_net_1, F_AWADDR_HADDR0(15) => VCC_net_1, 
        F_AWADDR_HADDR0(14) => VCC_net_1, F_AWADDR_HADDR0(13) => 
        VCC_net_1, F_AWADDR_HADDR0(12) => VCC_net_1, 
        F_AWADDR_HADDR0(11) => VCC_net_1, F_AWADDR_HADDR0(10) => 
        VCC_net_1, F_AWADDR_HADDR0(9) => VCC_net_1, 
        F_AWADDR_HADDR0(8) => VCC_net_1, F_AWADDR_HADDR0(7) => 
        VCC_net_1, F_AWADDR_HADDR0(6) => VCC_net_1, 
        F_AWADDR_HADDR0(5) => VCC_net_1, F_AWADDR_HADDR0(4) => 
        VCC_net_1, F_AWADDR_HADDR0(3) => VCC_net_1, 
        F_AWADDR_HADDR0(2) => VCC_net_1, F_AWADDR_HADDR0(1) => 
        VCC_net_1, F_AWADDR_HADDR0(0) => VCC_net_1, 
        F_AWBURST_HTRANS0(1) => GND_net_1, F_AWBURST_HTRANS0(0)
         => GND_net_1, F_AWID_HSEL0(3) => GND_net_1, 
        F_AWID_HSEL0(2) => GND_net_1, F_AWID_HSEL0(1) => 
        GND_net_1, F_AWID_HSEL0(0) => GND_net_1, 
        F_AWLEN_HBURST0(3) => GND_net_1, F_AWLEN_HBURST0(2) => 
        GND_net_1, F_AWLEN_HBURST0(1) => GND_net_1, 
        F_AWLEN_HBURST0(0) => GND_net_1, F_AWLOCK_HMASTLOCK0(1)
         => GND_net_1, F_AWLOCK_HMASTLOCK0(0) => GND_net_1, 
        F_AWSIZE_HSIZE0(1) => GND_net_1, F_AWSIZE_HSIZE0(0) => 
        GND_net_1, F_AWVALID_HWRITE0 => GND_net_1, F_BREADY => 
        GND_net_1, F_RMW_AXI => GND_net_1, F_RREADY => GND_net_1, 
        F_WDATA_HWDATA01(63) => VCC_net_1, F_WDATA_HWDATA01(62)
         => VCC_net_1, F_WDATA_HWDATA01(61) => VCC_net_1, 
        F_WDATA_HWDATA01(60) => VCC_net_1, F_WDATA_HWDATA01(59)
         => VCC_net_1, F_WDATA_HWDATA01(58) => VCC_net_1, 
        F_WDATA_HWDATA01(57) => VCC_net_1, F_WDATA_HWDATA01(56)
         => VCC_net_1, F_WDATA_HWDATA01(55) => VCC_net_1, 
        F_WDATA_HWDATA01(54) => VCC_net_1, F_WDATA_HWDATA01(53)
         => VCC_net_1, F_WDATA_HWDATA01(52) => VCC_net_1, 
        F_WDATA_HWDATA01(51) => VCC_net_1, F_WDATA_HWDATA01(50)
         => VCC_net_1, F_WDATA_HWDATA01(49) => VCC_net_1, 
        F_WDATA_HWDATA01(48) => VCC_net_1, F_WDATA_HWDATA01(47)
         => VCC_net_1, F_WDATA_HWDATA01(46) => VCC_net_1, 
        F_WDATA_HWDATA01(45) => VCC_net_1, F_WDATA_HWDATA01(44)
         => VCC_net_1, F_WDATA_HWDATA01(43) => VCC_net_1, 
        F_WDATA_HWDATA01(42) => VCC_net_1, F_WDATA_HWDATA01(41)
         => VCC_net_1, F_WDATA_HWDATA01(40) => VCC_net_1, 
        F_WDATA_HWDATA01(39) => VCC_net_1, F_WDATA_HWDATA01(38)
         => VCC_net_1, F_WDATA_HWDATA01(37) => VCC_net_1, 
        F_WDATA_HWDATA01(36) => VCC_net_1, F_WDATA_HWDATA01(35)
         => VCC_net_1, F_WDATA_HWDATA01(34) => VCC_net_1, 
        F_WDATA_HWDATA01(33) => VCC_net_1, F_WDATA_HWDATA01(32)
         => VCC_net_1, F_WDATA_HWDATA01(31) => VCC_net_1, 
        F_WDATA_HWDATA01(30) => VCC_net_1, F_WDATA_HWDATA01(29)
         => VCC_net_1, F_WDATA_HWDATA01(28) => VCC_net_1, 
        F_WDATA_HWDATA01(27) => VCC_net_1, F_WDATA_HWDATA01(26)
         => VCC_net_1, F_WDATA_HWDATA01(25) => VCC_net_1, 
        F_WDATA_HWDATA01(24) => VCC_net_1, F_WDATA_HWDATA01(23)
         => VCC_net_1, F_WDATA_HWDATA01(22) => VCC_net_1, 
        F_WDATA_HWDATA01(21) => VCC_net_1, F_WDATA_HWDATA01(20)
         => VCC_net_1, F_WDATA_HWDATA01(19) => VCC_net_1, 
        F_WDATA_HWDATA01(18) => VCC_net_1, F_WDATA_HWDATA01(17)
         => VCC_net_1, F_WDATA_HWDATA01(16) => VCC_net_1, 
        F_WDATA_HWDATA01(15) => VCC_net_1, F_WDATA_HWDATA01(14)
         => VCC_net_1, F_WDATA_HWDATA01(13) => VCC_net_1, 
        F_WDATA_HWDATA01(12) => VCC_net_1, F_WDATA_HWDATA01(11)
         => VCC_net_1, F_WDATA_HWDATA01(10) => VCC_net_1, 
        F_WDATA_HWDATA01(9) => VCC_net_1, F_WDATA_HWDATA01(8) => 
        VCC_net_1, F_WDATA_HWDATA01(7) => VCC_net_1, 
        F_WDATA_HWDATA01(6) => VCC_net_1, F_WDATA_HWDATA01(5) => 
        VCC_net_1, F_WDATA_HWDATA01(4) => VCC_net_1, 
        F_WDATA_HWDATA01(3) => VCC_net_1, F_WDATA_HWDATA01(2) => 
        VCC_net_1, F_WDATA_HWDATA01(1) => VCC_net_1, 
        F_WDATA_HWDATA01(0) => VCC_net_1, F_WID_HREADY01(3) => 
        GND_net_1, F_WID_HREADY01(2) => GND_net_1, 
        F_WID_HREADY01(1) => GND_net_1, F_WID_HREADY01(0) => 
        GND_net_1, F_WLAST => GND_net_1, F_WSTRB(7) => GND_net_1, 
        F_WSTRB(6) => GND_net_1, F_WSTRB(5) => GND_net_1, 
        F_WSTRB(4) => GND_net_1, F_WSTRB(3) => GND_net_1, 
        F_WSTRB(2) => GND_net_1, F_WSTRB(1) => GND_net_1, 
        F_WSTRB(0) => GND_net_1, F_WVALID => GND_net_1, 
        FPGA_MDDR_ARESET_N => VCC_net_1, MDDR_FABRIC_PADDR(10)
         => VCC_net_1, MDDR_FABRIC_PADDR(9) => VCC_net_1, 
        MDDR_FABRIC_PADDR(8) => VCC_net_1, MDDR_FABRIC_PADDR(7)
         => VCC_net_1, MDDR_FABRIC_PADDR(6) => VCC_net_1, 
        MDDR_FABRIC_PADDR(5) => VCC_net_1, MDDR_FABRIC_PADDR(4)
         => VCC_net_1, MDDR_FABRIC_PADDR(3) => VCC_net_1, 
        MDDR_FABRIC_PADDR(2) => VCC_net_1, MDDR_FABRIC_PENABLE
         => VCC_net_1, MDDR_FABRIC_PSEL => VCC_net_1, 
        MDDR_FABRIC_PWDATA(15) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(14) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(13) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(12) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(11) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(10) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(9) => VCC_net_1, MDDR_FABRIC_PWDATA(8)
         => VCC_net_1, MDDR_FABRIC_PWDATA(7) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(6) => VCC_net_1, MDDR_FABRIC_PWDATA(5)
         => VCC_net_1, MDDR_FABRIC_PWDATA(4) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(3) => VCC_net_1, MDDR_FABRIC_PWDATA(2)
         => VCC_net_1, MDDR_FABRIC_PWDATA(1) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(0) => VCC_net_1, MDDR_FABRIC_PWRITE
         => VCC_net_1, PRESET_N => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => GND_net_1, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => GND_net_1, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => GND_net_1, DM_IN(2)
         => GND_net_1, DM_IN(1) => GND_net_1, DM_IN(0) => 
        GND_net_1, DRAM_DQ_IN(17) => GND_net_1, DRAM_DQ_IN(16)
         => GND_net_1, DRAM_DQ_IN(15) => GND_net_1, 
        DRAM_DQ_IN(14) => GND_net_1, DRAM_DQ_IN(13) => GND_net_1, 
        DRAM_DQ_IN(12) => GND_net_1, DRAM_DQ_IN(11) => GND_net_1, 
        DRAM_DQ_IN(10) => GND_net_1, DRAM_DQ_IN(9) => GND_net_1, 
        DRAM_DQ_IN(8) => GND_net_1, DRAM_DQ_IN(7) => GND_net_1, 
        DRAM_DQ_IN(6) => GND_net_1, DRAM_DQ_IN(5) => GND_net_1, 
        DRAM_DQ_IN(4) => GND_net_1, DRAM_DQ_IN(3) => GND_net_1, 
        DRAM_DQ_IN(2) => GND_net_1, DRAM_DQ_IN(1) => GND_net_1, 
        DRAM_DQ_IN(0) => GND_net_1, DRAM_DQS_IN(2) => GND_net_1, 
        DRAM_DQS_IN(1) => GND_net_1, DRAM_DQS_IN(0) => GND_net_1, 
        DRAM_FIFO_WE_IN(1) => GND_net_1, DRAM_FIFO_WE_IN(0) => 
        GND_net_1, I2C0_SCL_USBC_DATA1_MGPIO31B_IN => GND_net_1, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => GND_net_1, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => GND_net_1, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => GND_net_1, MGPIO0B_IN
         => GND_net_1, MGPIO10B_IN => GND_net_1, MGPIO1B_IN => 
        GND_net_1, MGPIO25A_IN => GND_net_1, MGPIO26A_IN => 
        GND_net_1, MGPIO27A_IN => GND_net_1, MGPIO28A_IN => 
        GND_net_1, MGPIO29A_IN => GND_net_1, MGPIO2B_IN => 
        GND_net_1, MGPIO30A_IN => GND_net_1, MGPIO31A_IN => 
        GND_net_1, MGPIO3B_IN => GND_net_1, MGPIO4B_IN => 
        GND_net_1, MGPIO5B_IN => GND_net_1, MGPIO6B_IN => 
        GND_net_1, MGPIO7B_IN => GND_net_1, MGPIO8B_IN => 
        GND_net_1, MGPIO9B_IN => GND_net_1, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => GND_net_1, 
        MMUART0_DCD_MGPIO22B_IN => GND_net_1, 
        MMUART0_DSR_MGPIO20B_IN => GND_net_1, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => GND_net_1, 
        MMUART0_RI_MGPIO21B_IN => GND_net_1, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => GND_net_1, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => GND_net_1, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => GND_net_1, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => GND_net_1, 
        MMUART1_CTS_MGPIO13B_IN => GND_net_1, 
        MMUART1_DCD_MGPIO16B_IN => GND_net_1, 
        MMUART1_DSR_MGPIO14B_IN => GND_net_1, 
        MMUART1_DTR_MGPIO12B_IN => GND_net_1, 
        MMUART1_RI_MGPIO15B_IN => GND_net_1, 
        MMUART1_RTS_MGPIO11B_IN => GND_net_1, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => GND_net_1, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => GND_net_1, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => GND_net_1, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => GND_net_1, 
        RGMII_MDC_RMII_MDC_IN => GND_net_1, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => GND_net_1, 
        RGMII_RX_CLK_IN => GND_net_1, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => GND_net_1, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => GND_net_1, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => GND_net_1, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => GND_net_1, 
        RGMII_RXD3_USBB_DATA4_IN => GND_net_1, RGMII_TX_CLK_IN
         => GND_net_1, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => 
        GND_net_1, RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => GND_net_1, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => GND_net_1, 
        RGMII_TXD2_USBB_DATA5_IN => GND_net_1, 
        RGMII_TXD3_USBB_DATA6_IN => GND_net_1, 
        SPI0_SCK_USBA_XCLK_IN => GND_net_1, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => GND_net_1, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => GND_net_1, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => GND_net_1, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => GND_net_1, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => GND_net_1, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => GND_net_1, 
        SPI0_SS4_MGPIO19A_IN => GND_net_1, SPI0_SS5_MGPIO20A_IN
         => GND_net_1, SPI0_SS6_MGPIO21A_IN => GND_net_1, 
        SPI0_SS7_MGPIO22A_IN => GND_net_1, SPI1_SCK_IN => 
        GND_net_1, SPI1_SDI_MGPIO11A_IN => GND_net_1, 
        SPI1_SDO_MGPIO12A_IN => GND_net_1, SPI1_SS0_MGPIO13A_IN
         => GND_net_1, SPI1_SS1_MGPIO14A_IN => GND_net_1, 
        SPI1_SS2_MGPIO15A_IN => GND_net_1, SPI1_SS3_MGPIO16A_IN
         => GND_net_1, SPI1_SS4_MGPIO17A_IN => GND_net_1, 
        SPI1_SS5_MGPIO18A_IN => GND_net_1, SPI1_SS6_MGPIO23A_IN
         => GND_net_1, SPI1_SS7_MGPIO24A_IN => GND_net_1, 
        USBC_XCLK_IN => GND_net_1, USBD_DATA0_IN => GND_net_1, 
        USBD_DATA1_IN => GND_net_1, USBD_DATA2_IN => GND_net_1, 
        USBD_DATA3_IN => GND_net_1, USBD_DATA4_IN => GND_net_1, 
        USBD_DATA5_IN => GND_net_1, USBD_DATA6_IN => GND_net_1, 
        USBD_DATA7_MGPIO23B_IN => GND_net_1, USBD_DIR_IN => 
        GND_net_1, USBD_NXT_IN => GND_net_1, USBD_STP_IN => 
        GND_net_1, USBD_XCLK_IN => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => OPEN, DRAM_ADDR(15)
         => nc206, DRAM_ADDR(14) => nc174, DRAM_ADDR(13) => nc38, 
        DRAM_ADDR(12) => nc113, DRAM_ADDR(11) => nc218, 
        DRAM_ADDR(10) => nc106, DRAM_ADDR(9) => nc261, 
        DRAM_ADDR(8) => nc25, DRAM_ADDR(7) => nc1, DRAM_ADDR(6)
         => nc322, DRAM_ADDR(5) => nc299, DRAM_ADDR(4) => nc37, 
        DRAM_ADDR(3) => nc202, DRAM_ADDR(2) => nc144, 
        DRAM_ADDR(1) => nc153, DRAM_ADDR(0) => nc46, DRAM_BA(2)
         => nc258, DRAM_BA(1) => nc71, DRAM_BA(0) => nc124, 
        DRAM_CASN => OPEN, DRAM_CKE => OPEN, DRAM_CLK => OPEN, 
        DRAM_CSN => OPEN, DRAM_DM_RDQS_OUT(2) => nc332, 
        DRAM_DM_RDQS_OUT(1) => nc81, DRAM_DM_RDQS_OUT(0) => nc201, 
        DRAM_DQ_OUT(17) => nc168, DRAM_DQ_OUT(16) => nc323, 
        DRAM_DQ_OUT(15) => nc34, DRAM_DQ_OUT(14) => nc28, 
        DRAM_DQ_OUT(13) => nc115, DRAM_DQ_OUT(12) => nc264, 
        DRAM_DQ_OUT(11) => nc192, DRAM_DQ_OUT(10) => nc319, 
        DRAM_DQ_OUT(9) => nc134, DRAM_DQ_OUT(8) => nc32, 
        DRAM_DQ_OUT(7) => nc40, DRAM_DQ_OUT(6) => nc297, 
        DRAM_DQ_OUT(5) => nc99, DRAM_DQ_OUT(4) => nc75, 
        DRAM_DQ_OUT(3) => nc183, DRAM_DQ_OUT(2) => nc333, 
        DRAM_DQ_OUT(1) => nc288, DRAM_DQ_OUT(0) => nc85, 
        DRAM_DQS_OUT(2) => nc27, DRAM_DQS_OUT(1) => nc108, 
        DRAM_DQS_OUT(0) => nc325, DRAM_FIFO_WE_OUT(1) => nc16, 
        DRAM_FIFO_WE_OUT(0) => nc155, DRAM_ODT => OPEN, DRAM_RASN
         => OPEN, DRAM_RSTN => OPEN, DRAM_WEN => OPEN, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OUT => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => OPEN, MGPIO0B_OUT => 
        OPEN, MGPIO10B_OUT => OPEN, MGPIO1B_OUT => OPEN, 
        MGPIO25A_OUT => OPEN, MGPIO26A_OUT => OPEN, MGPIO27A_OUT
         => OPEN, MGPIO28A_OUT => OPEN, MGPIO29A_OUT => OPEN, 
        MGPIO2B_OUT => OPEN, MGPIO30A_OUT => OPEN, MGPIO31A_OUT
         => OPEN, MGPIO3B_OUT => OPEN, MGPIO4B_OUT => OPEN, 
        MGPIO5B_OUT => OPEN, MGPIO6B_OUT => OPEN, MGPIO7B_OUT => 
        OPEN, MGPIO8B_OUT => OPEN, MGPIO9B_OUT => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT => OPEN, 
        MMUART0_DCD_MGPIO22B_OUT => OPEN, 
        MMUART0_DSR_MGPIO20B_OUT => OPEN, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => OPEN, 
        MMUART1_CTS_MGPIO13B_OUT => OPEN, 
        MMUART1_DCD_MGPIO16B_OUT => OPEN, 
        MMUART1_DSR_MGPIO14B_OUT => OPEN, 
        MMUART1_DTR_MGPIO12B_OUT => OPEN, MMUART1_RI_MGPIO15B_OUT
         => OPEN, MMUART1_RTS_MGPIO11B_OUT => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => OPEN, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => OPEN, 
        RGMII_RXD3_USBB_DATA4_OUT => OPEN, RGMII_TX_CLK_OUT => 
        OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => OPEN, 
        RGMII_TXD2_USBB_DATA5_OUT => OPEN, 
        RGMII_TXD3_USBB_DATA6_OUT => OPEN, SPI0_SCK_USBA_XCLK_OUT
         => OPEN, SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => OPEN, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => OPEN, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => OPEN, 
        SPI0_SS4_MGPIO19A_OUT => OPEN, SPI0_SS5_MGPIO20A_OUT => 
        OPEN, SPI0_SS6_MGPIO21A_OUT => OPEN, 
        SPI0_SS7_MGPIO22A_OUT => OPEN, SPI1_SCK_OUT => OPEN, 
        SPI1_SDI_MGPIO11A_OUT => OPEN, SPI1_SDO_MGPIO12A_OUT => 
        OPEN, SPI1_SS0_MGPIO13A_OUT => OPEN, 
        SPI1_SS1_MGPIO14A_OUT => OPEN, SPI1_SS2_MGPIO15A_OUT => 
        OPEN, SPI1_SS3_MGPIO16A_OUT => OPEN, 
        SPI1_SS4_MGPIO17A_OUT => OPEN, SPI1_SS5_MGPIO18A_OUT => 
        OPEN, SPI1_SS6_MGPIO23A_OUT => OPEN, 
        SPI1_SS7_MGPIO24A_OUT => OPEN, USBC_XCLK_OUT => OPEN, 
        USBD_DATA0_OUT => OPEN, USBD_DATA1_OUT => OPEN, 
        USBD_DATA2_OUT => OPEN, USBD_DATA3_OUT => OPEN, 
        USBD_DATA4_OUT => OPEN, USBD_DATA5_OUT => OPEN, 
        USBD_DATA6_OUT => OPEN, USBD_DATA7_MGPIO23B_OUT => OPEN, 
        USBD_DIR_OUT => OPEN, USBD_NXT_OUT => OPEN, USBD_STP_OUT
         => OPEN, USBD_XCLK_OUT => OPEN, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => OPEN, DM_OE(2) => nc51, 
        DM_OE(1) => nc301, DM_OE(0) => nc33, DRAM_DQ_OE(17) => 
        nc204, DRAM_DQ_OE(16) => nc173, DRAM_DQ_OE(15) => nc278, 
        DRAM_DQ_OE(14) => nc169, DRAM_DQ_OE(13) => nc78, 
        DRAM_DQ_OE(12) => nc263, DRAM_DQ_OE(11) => nc24, 
        DRAM_DQ_OE(10) => nc88, DRAM_DQ_OE(9) => nc111, 
        DRAM_DQ_OE(8) => nc55, DRAM_DQ_OE(7) => nc10, 
        DRAM_DQ_OE(6) => nc22, DRAM_DQ_OE(5) => nc210, 
        DRAM_DQ_OE(4) => nc185, DRAM_DQ_OE(3) => nc143, 
        DRAM_DQ_OE(2) => nc248, DRAM_DQ_OE(1) => nc77, 
        DRAM_DQ_OE(0) => nc6, DRAM_DQS_OE(2) => nc109, 
        DRAM_DQS_OE(1) => nc87, DRAM_DQS_OE(0) => nc123, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => OPEN, MGPIO0B_OE => 
        OPEN, MGPIO10B_OE => OPEN, MGPIO1B_OE => OPEN, 
        MGPIO25A_OE => OPEN, MGPIO26A_OE => OPEN, MGPIO27A_OE => 
        OPEN, MGPIO28A_OE => OPEN, MGPIO29A_OE => OPEN, 
        MGPIO2B_OE => OPEN, MGPIO30A_OE => OPEN, MGPIO31A_OE => 
        OPEN, MGPIO3B_OE => OPEN, MGPIO4B_OE => OPEN, MGPIO5B_OE
         => OPEN, MGPIO6B_OE => OPEN, MGPIO7B_OE => OPEN, 
        MGPIO8B_OE => OPEN, MGPIO9B_OE => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => OPEN, 
        MMUART0_DCD_MGPIO22B_OE => OPEN, MMUART0_DSR_MGPIO20B_OE
         => OPEN, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => OPEN, 
        MMUART1_CTS_MGPIO13B_OE => OPEN, MMUART1_DCD_MGPIO16B_OE
         => OPEN, MMUART1_DSR_MGPIO14B_OE => OPEN, 
        MMUART1_DTR_MGPIO12B_OE => OPEN, MMUART1_RI_MGPIO15B_OE
         => OPEN, MMUART1_RTS_MGPIO11B_OE => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => OPEN, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => OPEN, 
        RGMII_RXD3_USBB_DATA4_OE => OPEN, RGMII_TX_CLK_OE => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => OPEN, 
        RGMII_TXD2_USBB_DATA5_OE => OPEN, 
        RGMII_TXD3_USBB_DATA6_OE => OPEN, SPI0_SCK_USBA_XCLK_OE
         => OPEN, SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => OPEN, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => OPEN, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => OPEN, 
        SPI0_SS4_MGPIO19A_OE => OPEN, SPI0_SS5_MGPIO20A_OE => 
        OPEN, SPI0_SS6_MGPIO21A_OE => OPEN, SPI0_SS7_MGPIO22A_OE
         => OPEN, SPI1_SCK_OE => OPEN, SPI1_SDI_MGPIO11A_OE => 
        OPEN, SPI1_SDO_MGPIO12A_OE => OPEN, SPI1_SS0_MGPIO13A_OE
         => OPEN, SPI1_SS1_MGPIO14A_OE => OPEN, 
        SPI1_SS2_MGPIO15A_OE => OPEN, SPI1_SS3_MGPIO16A_OE => 
        OPEN, SPI1_SS4_MGPIO17A_OE => OPEN, SPI1_SS5_MGPIO18A_OE
         => OPEN, SPI1_SS6_MGPIO23A_OE => OPEN, 
        SPI1_SS7_MGPIO24A_OE => OPEN, USBC_XCLK_OE => OPEN, 
        USBD_DATA0_OE => OPEN, USBD_DATA1_OE => OPEN, 
        USBD_DATA2_OE => OPEN, USBD_DATA3_OE => OPEN, 
        USBD_DATA4_OE => OPEN, USBD_DATA5_OE => OPEN, 
        USBD_DATA6_OE => OPEN, USBD_DATA7_MGPIO23B_OE => OPEN, 
        USBD_DIR_OE => OPEN, USBD_NXT_OE => OPEN, USBD_STP_OE => 
        OPEN, USBD_XCLK_OE => OPEN);
    
    MSS_ADLIB_INST_RNO_5 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_505, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_571, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[6]\);
    
    MSS_ADLIB_INST_RNO_25 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_525, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_591, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[26]\);
    
    MSS_ADLIB_INST_RNO_24 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_524, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_590, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[25]\);
    
    MSS_ADLIB_INST_RNO_45 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_3_4, B => line_4_4, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[11]\, D => 
        result_addr_net_0(1), Y => N_246);
    
    MSS_ADLIB_INST_RNO_1 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_501, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_567, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[2]\);
    
    MSS_ADLIB_INST_RNO_30 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_273, B => N_59, C => N_208, D => N_205, Y
         => \AMBA_SLAVE_0_HRDATA_S0_m[31]\);
    
    MSS_ADLIB_INST_RNO_44 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_3_3, B => line_4_3, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[10]\, D => 
        result_addr_net_0(1), Y => N_196);
    
    MSS_ADLIB_INST_RNO_33 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_274, B => N_273, C => line_7_4, D => N_246, 
        Y => \AMBA_SLAVE_0_HRDATA_S0_m_0_0[11]\);
    
    MSS_ADLIB_INST_RNO_26 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_526, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_592, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[27]\);
    
    MSS_ADLIB_INST_RNO_39 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_13, B => line_0_13, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[20]\, D => 
        result_addr_net_0(1), Y => N_199);
    
    MSS_ADLIB_INST_RNO_8 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_508, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_574, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[9]\);
    
    MSS_ADLIB_INST_RNO_6 : CFG3
      generic map(INIT => x"EC")

      port map(A => N_59, B => \AMBA_SLAVE_0_HRDATA_S0_m_0_0[7]\, 
        C => N_237, Y => \AMBA_SLAVE_0_HRDATA_S0_m[7]\);
    
    MSS_ADLIB_INST_RNO_46 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_3_13, B => line_4_13, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[20]\, D => 
        result_addr_net_0(1), Y => N_202);
    
    MSS_ADLIB_INST_RNO_31 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_274, B => N_273, C => line_7_0, D => N_240, 
        Y => \AMBA_SLAVE_0_HRDATA_S0_m_0_0[7]\);
    
    MSS_ADLIB_INST_RNO_55 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_0, B => line_2_0, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[7]\);
    
    MSS_ADLIB_INST_RNO_28 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_528, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_594, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[29]\);
    
    MSS_ADLIB_INST_RNO_54 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_24, B => line_6_24, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[31]\);
    
    MSS_ADLIB_INST_RNO_32 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_274, B => N_273, C => line_7_3, D => N_196, 
        Y => \AMBA_SLAVE_0_HRDATA_S0_m_0_0[10]\);
    
    MSS_ADLIB_INST_RNO_9 : CFG3
      generic map(INIT => x"EC")

      port map(A => N_59, B => \AMBA_SLAVE_0_HRDATA_S0_m_0_0[10]\, 
        C => N_188, Y => \AMBA_SLAVE_0_HRDATA_S0_m[10]\);
    
    MSS_ADLIB_INST_RNO_48 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_0, B => line_6_0, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[7]\);
    
    MSS_ADLIB_INST_RNO_15 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_515, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_581, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[16]\);
    
    MSS_ADLIB_INST_RNO_0 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_500, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_566, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[1]\);
    
    MSS_ADLIB_INST_RNO_14 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_514, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_580, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[15]\);
    
    MSS_ADLIB_INST_RNO_37 : CFG4
      generic map(INIT => x"AC0F")

      port map(A => line_3_d0, B => line_0_3, C => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_1_1[10]\, D => 
        result_addr_net_0(1), Y => N_188);
    
    MSS_ADLIB_INST_RNO_56 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_3, B => line_6_3, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[10]\);
    
    MSS_ADLIB_INST_RNO_16 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_516, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_582, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[17]\);
    
    MSS_ADLIB_INST_RNO_58 : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_13, B => line_6_13, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m_0_m3_0_2[20]\);
    
    MSS_ADLIB_INST_RNO_18 : CFG4
      generic map(INIT => x"80B0")

      port map(A => N_74, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_228, Y => N_34_i_0);
    
    MSS_ADLIB_INST_RNO_3 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_503, B => result_addr_net_0(0), C => 
        hready_m_xhdl339, D => N_569, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[4]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_system_sb_FABOSC_0_OSC is

    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );

end sha256_system_sb_FABOSC_0_OSC;

architecture DEF_ARCH of sha256_system_sb_FABOSC_0_OSC is 

  component RCOSC_25_50MHZ
    generic (FREQUENCY:real := 50.0);

    port( CLKOUT : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    I_RCOSC_25_50MHZ : RCOSC_25_50MHZ
      generic map(FREQUENCY => 50.0)

      port map(CLKOUT => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreResetP is

    port( MSS_READY                                       : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK                    : in    std_logic;
          sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic;
          sha256_system_sb_0_POWER_ON_RESET_N             : in    std_logic
        );

end CoreResetP;

architecture DEF_ARCH of CoreResetP is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \MSS_HPMS_READY_int\, \mss_ready_select\, VCC_net_1, 
        \POWER_ON_RESET_N_clk_base\, 
        \un6_fic_2_apb_m_preset_n_clk_base\, GND_net_1, 
        \mss_ready_state\, \RESET_N_M2F_clk_base\, 
        \RESET_N_M2F_q1\, \FIC_2_APB_M_PRESET_N_clk_base\, 
        \FIC_2_APB_M_PRESET_N_q1\, \MSS_HPMS_READY_int_3\, 
        \POWER_ON_RESET_N_q1\ : std_logic;

begin 


    RESET_N_M2F_clk_base : SLE
      port map(D => \RESET_N_M2F_q1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RESET_N_M2F_clk_base\);
    
    POWER_ON_RESET_N_clk_base : SLE
      port map(D => \POWER_ON_RESET_N_q1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \POWER_ON_RESET_N_clk_base\);
    
    mss_ready_select : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => 
        \un6_fic_2_apb_m_preset_n_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_select\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    mss_ready_state : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => 
        \RESET_N_M2F_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_state\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    un6_fic_2_apb_m_preset_n_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \FIC_2_APB_M_PRESET_N_clk_base\, B => 
        \mss_ready_state\, Y => 
        \un6_fic_2_apb_m_preset_n_clk_base\);
    
    RESET_N_M2F_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RESET_N_M2F_q1\);
    
    FIC_2_APB_M_PRESET_N_clk_base : SLE
      port map(D => \FIC_2_APB_M_PRESET_N_q1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FIC_2_APB_M_PRESET_N_clk_base\);
    
    POWER_ON_RESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \POWER_ON_RESET_N_q1\);
    
    MSS_HPMS_READY_int_RNIFQTF : CLKINT
      port map(A => \MSS_HPMS_READY_int\, Y => MSS_READY);
    
    FIC_2_APB_M_PRESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FIC_2_APB_M_PRESET_N_q1\);
    
    MSS_HPMS_READY_int_3 : CFG3
      generic map(INIT => x"E0")

      port map(A => \RESET_N_M2F_clk_base\, B => 
        \mss_ready_select\, C => \FIC_2_APB_M_PRESET_N_clk_base\, 
        Y => \MSS_HPMS_READY_int_3\);
    
    MSS_HPMS_READY_int : SLE
      port map(D => \MSS_HPMS_READY_int_3\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \MSS_HPMS_READY_int\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVEARBITER_0 is

    port( arbRegSMCurrentState                   : out   std_logic_vector(15 downto 14);
          MSS_READY                              : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK           : in    std_logic;
          N_14_i                                 : out   std_logic;
          N_19                                   : in    std_logic;
          N_165                                  : in    std_logic;
          m6                                     : out   std_logic;
          N_164                                  : in    std_logic;
          N_166                                  : in    std_logic;
          N_8                                    : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY : in    std_logic;
          N_158_i_0                              : out   std_logic
        );

end COREAHBLITE_SLAVEARBITER_0;

architecture DEF_ARCH of COREAHBLITE_SLAVEARBITER_0 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \arbRegSMCurrentState[15]_net_1\, VCC_net_1, 
        N_104_i_0, GND_net_1, \arbRegSMCurrentState[14]_net_1\, 
        N_106_i_0, \N_14_i\, \m6\, N_141, \N_8\ : std_logic;

begin 

    arbRegSMCurrentState(15) <= \arbRegSMCurrentState[15]_net_1\;
    arbRegSMCurrentState(14) <= \arbRegSMCurrentState[14]_net_1\;
    N_14_i <= \N_14_i\;
    m6 <= \m6\;
    N_8 <= \N_8\;

    \arbRegSMCurrentState_RNIUAEK[14]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => N_19, B => \arbRegSMCurrentState[14]_net_1\, 
        C => \N_14_i\, Y => \N_8\);
    
    \arbRegSMCurrentState[15]\ : SLE
      port map(D => N_104_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[15]_net_1\);
    
    \arbRegSMCurrentState_RNO_0[14]\ : CFG4
      generic map(INIT => x"7F00")

      port map(A => N_164, B => N_166, C => \N_14_i\, D => \m6\, 
        Y => N_141);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \arbRegSMCurrentState_RNIBN4P[14]\ : CFG4
      generic map(INIT => x"0111")

      port map(A => \arbRegSMCurrentState[14]_net_1\, B => 
        \arbRegSMCurrentState[15]_net_1\, C => N_165, D => 
        \N_14_i\, Y => \m6\);
    
    \arbRegSMCurrentState_RNO[15]\ : CFG3
      generic map(INIT => x"54")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \N_8\, C => \arbRegSMCurrentState[15]_net_1\, Y => 
        N_104_i_0);
    
    \arbRegSMCurrentState[14]\ : SLE
      port map(D => N_106_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[14]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \arbRegSMCurrentState_RNIJN5M[14]\ : CFG4
      generic map(INIT => x"FCEC")

      port map(A => \arbRegSMCurrentState[14]_net_1\, B => 
        \arbRegSMCurrentState[15]_net_1\, C => N_19, D => 
        \N_14_i\, Y => N_158_i_0);
    
    \arbRegSMCurrentState[2]\ : SLE
      port map(D => GND_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_19, ALn => 
        MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \N_14_i\);
    
    \arbRegSMCurrentState_RNO[14]\ : CFG4
      generic map(INIT => x"00AE")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \arbRegSMCurrentState[14]_net_1\, C => N_19, D => N_141, 
        Y => N_106_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVESTAGE_1 is

    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA : in    std_logic_vector(31 downto 0);
          AHB_slave_dummy_0_mem_wdata                        : out   std_logic_vector(31 downto 0);
          arbRegSMCurrentState                               : out   std_logic_vector(15 downto 14);
          hwdata10                                           : out   std_logic;
          MSS_READY                                          : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                       : in    std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY             : in    std_logic;
          N_14_i                                             : out   std_logic;
          N_19                                               : in    std_logic;
          N_165                                              : in    std_logic;
          m6                                                 : out   std_logic;
          N_164                                              : in    std_logic;
          N_166                                              : in    std_logic;
          N_8                                                : out   std_logic
        );

end COREAHBLITE_SLAVESTAGE_1;

architecture DEF_ARCH of COREAHBLITE_SLAVESTAGE_1 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVEARBITER_0
    port( arbRegSMCurrentState                   : out   std_logic_vector(15 downto 14);
          MSS_READY                              : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK           : in    std_logic := 'U';
          N_14_i                                 : out   std_logic;
          N_19                                   : in    std_logic := 'U';
          N_165                                  : in    std_logic := 'U';
          m6                                     : out   std_logic;
          N_164                                  : in    std_logic := 'U';
          N_166                                  : in    std_logic := 'U';
          N_8                                    : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY : in    std_logic := 'U';
          N_158_i_0                              : out   std_logic
        );
  end component;

    signal \hwdata10\, VCC_net_1, N_158_i_0, GND_net_1
         : std_logic;

    for all : COREAHBLITE_SLAVEARBITER_0
	Use entity work.COREAHBLITE_SLAVEARBITER_0(DEF_ARCH);
begin 

    hwdata10 <= \hwdata10\;

    \masterDataInProg_RNI5BHU_25[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(15));
    
    \masterDataInProg_RNI5BHU_30[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(10));
    
    \masterDataInProg_RNI5BHU_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(6));
    
    \masterDataInProg_RNI5BHU_2[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(8));
    
    \masterDataInProg_RNI5BHU_23[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(17));
    
    \masterDataInProg_RNI5BHU_1[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(9));
    
    \masterDataInProg_RNI5BHU_28[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(12));
    
    \masterDataInProg_RNI5BHU_24[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(16));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \masterDataInProg_RNI5BHU_22[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(18));
    
    \masterDataInProg_RNI5BHU_6[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(4));
    
    \masterDataInProg_RNI5BHU_7[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(3));
    
    \masterDataInProg_RNI5BHU_16[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(24));
    
    \masterDataInProg_RNI5BHU_5[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(5));
    
    \masterDataInProg_RNI5BHU_27[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(13));
    
    \masterDataInProg_RNI5BHU_10[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(30));
    
    \masterDataInProg_RNI5BHU_0[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(0));
    
    \masterDataInProg_RNI5BHU_29[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(11));
    
    \masterDataInProg_RNI5BHU_15[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(25));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \masterDataInProg_RNI5BHU_21[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(19));
    
    \masterDataInProg[0]\ : SLE
      port map(D => N_158_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \hwdata10\);
    
    \masterDataInProg_RNI5BHU_13[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(27));
    
    \masterDataInProg_RNI5BHU[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(1));
    
    \masterDataInProg_RNI5BHU_18[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(22));
    
    \masterDataInProg_RNI5BHU_14[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(26));
    
    \masterDataInProg_RNI5BHU_12[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(28));
    
    \masterDataInProg_RNI5BHU_8[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(2));
    
    \masterDataInProg_RNI5BHU_17[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(23));
    
    slave_arbiter : COREAHBLITE_SLAVEARBITER_0
      port map(arbRegSMCurrentState(15) => 
        arbRegSMCurrentState(15), arbRegSMCurrentState(14) => 
        arbRegSMCurrentState(14), MSS_READY => MSS_READY, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, N_14_i => N_14_i, N_19 => 
        N_19, N_165 => N_165, m6 => m6, N_164 => N_164, N_166 => 
        N_166, N_8 => N_8, sha256_system_sb_0_AMBA_SLAVE_0_HREADY
         => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, N_158_i_0 => 
        N_158_i_0);
    
    \masterDataInProg_RNI5BHU_9[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(31));
    
    \masterDataInProg_RNI5BHU_3[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(7));
    
    \masterDataInProg_RNI5BHU_19[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(21));
    
    \masterDataInProg_RNI5BHU_26[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(14));
    
    \masterDataInProg_RNI5BHU_11[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(29));
    
    \masterDataInProg_RNI5BHU_20[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(20));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_DEFAULTSLAVESM_0 is

    port( SDATASELInt                  : in    std_logic_vector(1 to 1);
          defSlaveSMCurrentState       : out   std_logic;
          MSS_READY                    : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK : in    std_logic;
          N_135                        : in    std_logic
        );

end COREAHBLITE_DEFAULTSLAVESM_0;

architecture DEF_ARCH of COREAHBLITE_DEFAULTSLAVESM_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal defSlaveSMCurrentState_net_1, VCC_net_1, N_17_i_0, 
        GND_net_1 : std_logic;

begin 

    defSlaveSMCurrentState <= defSlaveSMCurrentState_net_1;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    defSlaveSMCurrentState_RNO : CFG3
      generic map(INIT => x"45")

      port map(A => defSlaveSMCurrentState_net_1, B => 
        SDATASELInt(1), C => N_135, Y => N_17_i_0);
    
    \defSlaveSMCurrentState\ : SLE
      port map(D => N_17_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        defSlaveSMCurrentState_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MASTERSTAGE_2_1_0_1_0 is

    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1);
          arbRegSMCurrentState                                 : in    std_logic_vector(15 downto 14);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic;
          result_addr_net_0_0                                  : in    std_logic;
          result_addr_net_0_3                                  : in    std_logic;
          MSS_READY                                            : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic;
          N_19                                                 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic;
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_165                                                : out   std_logic;
          N_166                                                : out   std_logic;
          N_164                                                : out   std_logic;
          N_114                                                : out   std_logic;
          N_115                                                : out   std_logic;
          N_116                                                : out   std_logic;
          N_117                                                : out   std_logic;
          N_118                                                : out   std_logic;
          N_119                                                : out   std_logic;
          N_14_i                                               : in    std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic;
          hwdata10                                             : in    std_logic;
          ren_pos                                              : in    std_logic;
          N_273                                                : out   std_logic;
          m6                                                   : in    std_logic;
          N_274                                                : out   std_logic;
          N_59                                                 : out   std_logic;
          N_8                                                  : in    std_logic;
          N_31                                                 : out   std_logic;
          defSlaveSMCurrentState                               : out   std_logic;
          N_23_i_0                                             : out   std_logic
        );

end COREAHBLITE_MASTERSTAGE_2_1_0_1_0;

architecture DEF_ARCH of COREAHBLITE_MASTERSTAGE_2_1_0_1_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_DEFAULTSLAVESM_0
    port( SDATASELInt                  : in    std_logic_vector(1 to 1) := (others => 'U');
          defSlaveSMCurrentState       : out   std_logic;
          MSS_READY                    : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK : in    std_logic := 'U';
          N_135                        : in    std_logic := 'U'
        );
  end component;

    signal \SDATASELInt[1]_net_1\, VCC_net_1, \SADDRSEL[1]\, 
        N_21_i_0, GND_net_1, \SDATASELInt[2]_net_1\, 
        \SADDRSEL[2]\, \SDATASELInt[3]_net_1\, \SADDRSEL[3]\, 
        \SDATASELInt[4]_net_1\, \SADDRSEL[4]\, 
        \SDATASELInt[5]_net_1\, \SADDRSEL[5]\, 
        \SDATASELInt[6]_net_1\, \SADDRSEL[6]\, 
        \SDATASELInt[7]_net_1\, \SADDRSEL[7]\, 
        \SDATASELInt[8]_net_1\, \SADDRSEL[8]\, 
        \SDATASELInt[9]_net_1\, \SADDRSEL[9]\, 
        \SDATASELInt[10]_net_1\, \SADDRSEL[10]\, 
        \SDATASELInt[11]_net_1\, \SADDRSEL[11]\, 
        \SDATASELInt[12]_net_1\, \SADDRSEL[12]\, 
        \SDATASELInt[13]_net_1\, \SADDRSEL[13]\, 
        \SDATASELInt[14]_net_1\, \SADDRSEL[14]\, 
        \SDATASELInt[15]_net_1\, N_137, \regHADDR[2]_net_1\, 
        masterAddrClockEnable, \regHADDR[3]_net_1\, 
        \regHADDR[4]_net_1\, \regHADDR[5]_net_1\, 
        \regHADDR[6]_net_1\, \xhdl1222[0]\, \N_19\, \regHWRITE\, 
        regHTRANS_net_1, masterRegAddrSel_net_1, 
        d_masterRegAddrSel, \N_165\, \N_166\, 
        \masterAddrClockEnable_0_a2_1_0_s_a0_2\, \N_164\, N_131, 
        N_147, N_126, hready_m_xhdl343_10, N_162, HREADY_m1_e_0, 
        \masterAddrClockEnable_0_a2_1_0_s_a0_3\, N_53, N_54, N_55, 
        N_190, N_135, hready_m_xhdl347_2_0, 
        \un1_hready_m_xhdl339_2_i_a2_2_0\, 
        un1_hready_m_xhdl339_2_i_a2_out, \hready_m_xhdl339\, 
        \masterAddrClockEnable_0_a2_1_c_0\, N_148, 
        \un1_hready_m_xhdl339_2_i_0_0\, N_128, 
        \masterAddrClockEnable_0_a2_1_c\, N_43, N_90, 
        masterAddrClockEnable_0_a2_1_0_out, N_154, 
        \un1_hready_m_xhdl339_2_i_0_2\, \N_31\, 
        \defSlaveSMCurrentState\, \masterAddrClockEnable_0_a2_0\
         : std_logic;

    for all : COREAHBLITE_DEFAULTSLAVESM_0
	Use entity work.COREAHBLITE_DEFAULTSLAVESM_0(DEF_ARCH);
begin 

    N_19 <= \N_19\;
    regHTRANS <= regHTRANS_net_1;
    masterRegAddrSel <= masterRegAddrSel_net_1;
    N_165 <= \N_165\;
    N_166 <= \N_166\;
    N_164 <= \N_164\;
    hready_m_xhdl339 <= \hready_m_xhdl339\;
    N_31 <= \N_31\;
    defSlaveSMCurrentState <= \defSlaveSMCurrentState\;

    un1_hready_m_xhdl339_2_i_0_2_RNIJDRL3 : CFG4
      generic map(INIT => x"00CD")

      port map(A => N_43, B => \defSlaveSMCurrentState\, C => 
        \un1_hready_m_xhdl339_2_i_0_2\, D => N_128, Y => N_23_i_0);
    
    \PREGATEDHADDR_i_m2[6]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, C
         => \regHADDR[6]_net_1\, Y => N_114);
    
    d_masterRegAddrSel_0_o2_0 : CFG4
      generic map(INIT => x"5700")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        arbRegSMCurrentState(15), C => N_8, D => \N_165\, Y => 
        N_154);
    
    un1_hready_m_xhdl339_2_i_o2 : CFG4
      generic map(INIT => x"0112")

      port map(A => \SDATASELInt[11]_net_1\, B => \xhdl1222[0]\, 
        C => \SDATASELInt[15]_net_1\, D => 
        \SDATASELInt[14]_net_1\, Y => N_53);
    
    \PREGATEDHADDR_i_m2[3]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, C
         => \regHADDR[3]_net_1\, Y => N_117);
    
    un1_hready_m_xhdl339_2_i_a2_14 : CFG4
      generic map(INIT => x"1300")

      port map(A => \xhdl1222[0]\, B => \SDATASELInt[1]_net_1\, C
         => N_135, D => hready_m_xhdl343_10, Y => N_148);
    
    \SADDRSEL_0_a2[6]\ : CFG4
      generic map(INIT => x"0040")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => N_162, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, D
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        Y => \SADDRSEL[6]\);
    
    masterAddrClockEnable_0_a2_0 : CFG4
      generic map(INIT => x"8088")

      port map(A => \N_164\, B => \N_166\, C => 
        \defSlaveSMCurrentState\, D => \N_31\, Y => 
        \masterAddrClockEnable_0_a2_0\);
    
    hready_m_xhdl339_0_a2_RNI6IGQ : CFG3
      generic map(INIT => x"70")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        hwdata10, C => \hready_m_xhdl339\, Y => N_128);
    
    un1_hready_m_xhdl339_2_i_a2_13 : CFG3
      generic map(INIT => x"01")

      port map(A => \SDATASELInt[4]_net_1\, B => 
        \SDATASELInt[3]_net_1\, C => \SDATASELInt[2]_net_1\, Y
         => N_147);
    
    masterAddrClockEnable_0_a2_1_c_0 : CFG4
      generic map(INIT => x"5155")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        N_135, C => \SDATASELInt[1]_net_1\, D => \xhdl1222[0]\, Y
         => \masterAddrClockEnable_0_a2_1_c_0\);
    
    hready_m_xhdl339_0_a2_RNII7CF : CFG3
      generic map(INIT => x"80")

      port map(A => ren_pos, B => \hready_m_xhdl339\, C => 
        result_addr_net_0_0, Y => N_273);
    
    \SADDRSEL_0_a2[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, B
         => \N_164\, C => N_162, Y => \SADDRSEL[3]\);
    
    \masterRegAddrSel\ : SLE
      port map(D => d_masterRegAddrSel, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => masterRegAddrSel_net_1);
    
    \regHTRANS\ : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => masterAddrClockEnable, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => regHTRANS_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \SADDRSEL_0_a2[12]\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => \N_166\, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, Y
         => \SADDRSEL[12]\);
    
    \SADDRSEL_0_a2[4]\ : CFG3
      generic map(INIT => x"40")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => \N_166\, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, Y
         => \SADDRSEL[4]\);
    
    masterAddrClockEnable_0_a2_1_0_s_a0_2 : CFG2
      generic map(INIT => x"1")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        Y => \masterAddrClockEnable_0_a2_1_0_s_a0_2\);
    
    \SADDRSEL_0_a2[14]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => N_162, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, D
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        Y => \SADDRSEL[14]\);
    
    \SADDRSEL_0_a2[10]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => N_162, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, D
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        Y => \SADDRSEL[10]\);
    
    \PREGATEDHADDR_i_m2[5]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, C
         => \regHADDR[5]_net_1\, Y => N_115);
    
    un1_hready_m_xhdl339_2_i_a2_2_0 : CFG4
      generic map(INIT => x"0448")

      port map(A => \SDATASELInt[2]_net_1\, B => 
        hready_m_xhdl347_2_0, C => \SDATASELInt[4]_net_1\, D => 
        \SDATASELInt[3]_net_1\, Y => 
        \un1_hready_m_xhdl339_2_i_a2_2_0\);
    
    \SADDRSEL_0_a2[8]\ : CFG3
      generic map(INIT => x"08")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => \N_166\, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, Y
         => \SADDRSEL[8]\);
    
    un1_hready_m_xhdl339_2_i_0_0 : CFG4
      generic map(INIT => x"BF20")

      port map(A => \SDATASELInt[1]_net_1\, B => \xhdl1222[0]\, C
         => N_135, D => un1_hready_m_xhdl339_2_i_a2_out, Y => 
        \un1_hready_m_xhdl339_2_i_0_0\);
    
    \regHADDR[5]\ : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => 
        masterAddrClockEnable, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \regHADDR[5]_net_1\);
    
    \SDATASELInt[4]\ : SLE
      port map(D => \SADDRSEL[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[4]_net_1\);
    
    \SADDRSEL_0_a2_1[10]\ : CFG3
      generic map(INIT => x"20")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, B
         => masterRegAddrSel_net_1, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), Y
         => N_162);
    
    \regHADDR[2]\ : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => 
        masterAddrClockEnable, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \regHADDR[2]_net_1\);
    
    \SDATASELInt[15]\ : SLE
      port map(D => N_137, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_21_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[15]_net_1\);
    
    \SDATASELInt[14]\ : SLE
      port map(D => \SADDRSEL[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[14]_net_1\);
    
    GATEDHWRITE_i_m2 : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, C => 
        \regHWRITE\, Y => N_119);
    
    \SDATASELInt[2]\ : SLE
      port map(D => \SADDRSEL[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[2]_net_1\);
    
    \PREGATEDHADDR_i_m2[4]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, C
         => \regHADDR[4]_net_1\, Y => N_116);
    
    hready_m_xhdl339_0_a2 : CFG3
      generic map(INIT => x"08")

      port map(A => \xhdl1222[0]\, B => N_135, C => 
        \SDATASELInt[1]_net_1\, Y => \hready_m_xhdl339\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    hready_m_xhdl339_10_0_a2_0_a2 : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt[8]_net_1\, B => 
        \SDATASELInt[7]_net_1\, C => \SDATASELInt[6]_net_1\, D
         => \SDATASELInt[5]_net_1\, Y => hready_m_xhdl343_10);
    
    hready_m_xhdl339_0_a2_RNILTVP : CFG4
      generic map(INIT => x"0080")

      port map(A => ren_pos, B => \hready_m_xhdl339\, C => 
        result_addr_net_0_3, D => result_addr_net_0_0, Y => N_274);
    
    un1_hready_m_xhdl339_2_i_0_RNI6NON : CFG4
      generic map(INIT => x"8ACF")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \defSlaveSMCurrentState\, C => \N_31\, D => 
        \hready_m_xhdl339\, Y => N_21_i_0);
    
    un1_hready_m_xhdl339_2_i_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \un1_hready_m_xhdl339_2_i_0_2\, B => N_43, Y
         => \N_31\);
    
    \SADDRSEL_0_a2_1[15]\ : CFG2
      generic map(INIT => x"8")

      port map(A => masterRegAddrSel_net_1, B => regHTRANS_net_1, 
        Y => \N_165\);
    
    \SADDRSEL_0_a2[7]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => N_162, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, D
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        Y => \SADDRSEL[7]\);
    
    masterAddrClockEnable_0_a2_1_c : CFG3
      generic map(INIT => x"C4")

      port map(A => arbRegSMCurrentState(14), B => 
        \masterAddrClockEnable_0_a2_1_c_0\, C => \N_19\, Y => 
        \masterAddrClockEnable_0_a2_1_c\);
    
    \regHADDR[6]\ : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => 
        masterAddrClockEnable, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \regHADDR[6]_net_1\);
    
    \SDATASELInt[13]\ : SLE
      port map(D => \SADDRSEL[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[13]_net_1\);
    
    \SADDRSEL_0_a2_0[15]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => N_162, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, D
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        Y => N_137);
    
    \SADDRSEL_0_a2[11]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => N_162, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, D
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        Y => \SADDRSEL[11]\);
    
    regHWRITE : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => 
        masterAddrClockEnable, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \regHWRITE\);
    
    hready_m_xhdl340_2_0_0_a2_0_a2 : CFG3
      generic map(INIT => x"40")

      port map(A => \xhdl1222[0]\, B => N_131, C => N_126, Y => 
        hready_m_xhdl347_2_0);
    
    \SDATASELInt[9]\ : SLE
      port map(D => \SADDRSEL[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[9]_net_1\);
    
    \SDATASELInt[1]\ : SLE
      port map(D => \SADDRSEL[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[1]_net_1\);
    
    \SDATASELInt[12]\ : SLE
      port map(D => \SADDRSEL[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[12]_net_1\);
    
    \SDATASELInt[0]\ : SLE
      port map(D => \N_19\, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_21_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \xhdl1222[0]\);
    
    \SADDRSEL_0_a2_0[9]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, B
         => masterRegAddrSel_net_1, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, D
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        Y => N_190);
    
    masterAddrClockEnable_0_a2_1_0_s_a0_3 : CFG4
      generic map(INIT => x"4000")

      port map(A => masterRegAddrSel_net_1, B => N_14_i, C => 
        \masterAddrClockEnable_0_a2_1_0_s_a0_2\, D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), Y
         => \masterAddrClockEnable_0_a2_1_0_s_a0_3\);
    
    \SDATASELInt[5]\ : SLE
      port map(D => \SADDRSEL[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[5]_net_1\);
    
    d_masterRegAddrSel_0 : CFG4
      generic map(INIT => x"FCEC")

      port map(A => \masterAddrClockEnable_0_a2_1_c\, B => N_154, 
        C => \masterAddrClockEnable_0_a2_0\, D => 
        masterAddrClockEnable_0_a2_1_0_out, Y => 
        d_masterRegAddrSel);
    
    \regHADDR[3]\ : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => 
        masterAddrClockEnable, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \regHADDR[3]_net_1\);
    
    \SADDRSEL_0_a2[5]\ : CFG3
      generic map(INIT => x"40")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => N_190, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, Y
         => \SADDRSEL[5]\);
    
    \SDATASELInt_RNIDU2C1[11]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt[11]_net_1\, B => \xhdl1222[0]\, 
        C => \SDATASELInt[15]_net_1\, D => 
        \SDATASELInt[14]_net_1\, Y => HREADY_m1_e_0);
    
    \SADDRSEL_0_a2_0[1]\ : CFG2
      generic map(INIT => x"1")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        Y => \N_164\);
    
    un1_hready_m_xhdl339_1_1_0_a2_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => hready_m_xhdl343_10, B => N_126, C => N_131, 
        D => N_147, Y => N_135);
    
    \SDATASELInt[3]\ : SLE
      port map(D => \SADDRSEL[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[3]_net_1\);
    
    un1_hready_m_xhdl339_2_i_o2_0_RNIGAAE2 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_147, B => N_148, C => N_54, D => 
        HREADY_m1_e_0, Y => N_43);
    
    \PREGATEDHADDR_i_m2[2]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, C
         => \regHADDR[2]_net_1\, Y => N_118);
    
    \SADDRSEL_0_a2_0[8]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, B
         => masterRegAddrSel_net_1, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, D
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        Y => \N_166\);
    
    un1_hready_m_xhdl339_2_i_0_2 : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \un1_hready_m_xhdl339_2_i_a2_2_0\, B => N_148, 
        C => \un1_hready_m_xhdl339_2_i_0_0\, D => N_90, Y => 
        \un1_hready_m_xhdl339_2_i_0_2\);
    
    \SDATASELInt[7]\ : SLE
      port map(D => \SADDRSEL[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[7]_net_1\);
    
    un1_hready_m_xhdl339_2_i_a2_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_53, B => N_147, C => N_148, D => N_126, Y
         => N_90);
    
    \SADDRSEL_0_a2[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_190, B => \N_164\, Y => \SADDRSEL[1]\);
    
    \SADDRSEL_0_a2[13]\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => N_190, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, Y
         => \SADDRSEL[13]\);
    
    masterAddrClockEnable_0_a2_1_0_s_0 : CFG4
      generic map(INIT => x"0070")

      port map(A => \N_164\, B => 
        \masterAddrClockEnable_0_a2_1_0_s_a0_3\, C => m6, D => 
        N_128, Y => masterAddrClockEnable_0_a2_1_0_out);
    
    \SDATASELInt[6]\ : SLE
      port map(D => \SADDRSEL[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[6]_net_1\);
    
    \SADDRSEL_0_a2[2]\ : CFG3
      generic map(INIT => x"40")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, B
         => \N_164\, C => N_162, Y => \SADDRSEL[2]\);
    
    hready_m_xhdl339_0_a2_RNILTVP_0 : CFG4
      generic map(INIT => x"0008")

      port map(A => ren_pos, B => \hready_m_xhdl339\, C => 
        result_addr_net_0_3, D => result_addr_net_0_0, Y => N_59);
    
    un1_hready_m_xhdl339_2_i_a2_10_0_a2_0 : CFG3
      generic map(INIT => x"01")

      port map(A => \SDATASELInt[15]_net_1\, B => 
        \SDATASELInt[14]_net_1\, C => \SDATASELInt[11]_net_1\, Y
         => N_131);
    
    \SDATASELInt[11]\ : SLE
      port map(D => \SADDRSEL[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[11]_net_1\);
    
    un1_hready_m_xhdl339_2_i_o2_0 : CFG4
      generic map(INIT => x"0116")

      port map(A => \SDATASELInt[13]_net_1\, B => 
        \SDATASELInt[12]_net_1\, C => \SDATASELInt[10]_net_1\, D
         => \SDATASELInt[9]_net_1\, Y => N_54);
    
    \SDATASELInt[8]\ : SLE
      port map(D => \SADDRSEL[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[8]_net_1\);
    
    un1_hready_m_xhdl339_2_i_a2_s : CFG4
      generic map(INIT => x"2000")

      port map(A => N_55, B => \SDATASELInt[1]_net_1\, C => 
        hready_m_xhdl347_2_0, D => N_147, Y => 
        un1_hready_m_xhdl339_2_i_a2_out);
    
    \SADDRSEL_0[0]\ : CFG4
      generic map(INIT => x"CCDC")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, B
         => \N_165\, C => \N_166\, D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, Y
         => \N_19\);
    
    \regHADDR[4]\ : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => 
        masterAddrClockEnable, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \regHADDR[4]_net_1\);
    
    un1_hready_m_xhdl339_2_i_o2_1 : CFG4
      generic map(INIT => x"0116")

      port map(A => \SDATASELInt[8]_net_1\, B => 
        \SDATASELInt[7]_net_1\, C => \SDATASELInt[6]_net_1\, D
         => \SDATASELInt[5]_net_1\, Y => N_55);
    
    un1_hready_m_xhdl339_2_i_a2_11_0_a2 : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt[13]_net_1\, B => 
        \SDATASELInt[12]_net_1\, C => \SDATASELInt[10]_net_1\, D
         => \SDATASELInt[9]_net_1\, Y => N_126);
    
    \SDATASELInt[10]\ : SLE
      port map(D => \SADDRSEL[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[10]_net_1\);
    
    masterAddrClockEnable_0_a2 : CFG3
      generic map(INIT => x"A8")

      port map(A => \masterAddrClockEnable_0_a2_0\, B => 
        masterAddrClockEnable_0_a2_1_0_out, C => 
        \masterAddrClockEnable_0_a2_1_c\, Y => 
        masterAddrClockEnable);
    
    \SADDRSEL_0_a2[9]\ : CFG3
      generic map(INIT => x"08")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => N_190, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, Y
         => \SADDRSEL[9]\);
    
    default_slave_sm : COREAHBLITE_DEFAULTSLAVESM_0
      port map(SDATASELInt(1) => \SDATASELInt[1]_net_1\, 
        defSlaveSMCurrentState => \defSlaveSMCurrentState\, 
        MSS_READY => MSS_READY, sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, N_135 => N_135);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MATRIX4X16 is

    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1);
          arbRegSMCurrentState                                 : out   std_logic_vector(15 downto 14);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0);
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic;
          result_addr_net_0_0                                  : in    std_logic;
          result_addr_net_0_3                                  : in    std_logic;
          MSS_READY                                            : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic;
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_165                                                : out   std_logic;
          N_164                                                : out   std_logic;
          N_114                                                : out   std_logic;
          N_115                                                : out   std_logic;
          N_116                                                : out   std_logic;
          N_117                                                : out   std_logic;
          N_118                                                : out   std_logic;
          N_119                                                : out   std_logic;
          N_14_i                                               : out   std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic;
          ren_pos                                              : in    std_logic;
          N_273                                                : out   std_logic;
          N_274                                                : out   std_logic;
          N_59                                                 : out   std_logic;
          N_31                                                 : out   std_logic;
          defSlaveSMCurrentState                               : out   std_logic;
          N_23_i_0                                             : out   std_logic
        );

end COREAHBLITE_MATRIX4X16;

architecture DEF_ARCH of COREAHBLITE_MATRIX4X16 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVESTAGE_1
    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA : in    std_logic_vector(31 downto 0) := (others => 'U');
          AHB_slave_dummy_0_mem_wdata                        : out   std_logic_vector(31 downto 0);
          arbRegSMCurrentState                               : out   std_logic_vector(15 downto 14);
          hwdata10                                           : out   std_logic;
          MSS_READY                                          : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                       : in    std_logic := 'U';
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY             : in    std_logic := 'U';
          N_14_i                                             : out   std_logic;
          N_19                                               : in    std_logic := 'U';
          N_165                                              : in    std_logic := 'U';
          m6                                                 : out   std_logic;
          N_164                                              : in    std_logic := 'U';
          N_166                                              : in    std_logic := 'U';
          N_8                                                : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MASTERSTAGE_2_1_0_1_0
    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1) := (others => 'U');
          arbRegSMCurrentState                                 : in    std_logic_vector(15 downto 14) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic := 'U';
          result_addr_net_0_0                                  : in    std_logic := 'U';
          result_addr_net_0_3                                  : in    std_logic := 'U';
          MSS_READY                                            : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic := 'U';
          N_19                                                 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_165                                                : out   std_logic;
          N_166                                                : out   std_logic;
          N_164                                                : out   std_logic;
          N_114                                                : out   std_logic;
          N_115                                                : out   std_logic;
          N_116                                                : out   std_logic;
          N_117                                                : out   std_logic;
          N_118                                                : out   std_logic;
          N_119                                                : out   std_logic;
          N_14_i                                               : in    std_logic := 'U';
          hready_m_xhdl339                                     : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic := 'U';
          hwdata10                                             : in    std_logic := 'U';
          ren_pos                                              : in    std_logic := 'U';
          N_273                                                : out   std_logic;
          m6                                                   : in    std_logic := 'U';
          N_274                                                : out   std_logic;
          N_59                                                 : out   std_logic;
          N_8                                                  : in    std_logic := 'U';
          N_31                                                 : out   std_logic;
          defSlaveSMCurrentState                               : out   std_logic;
          N_23_i_0                                             : out   std_logic
        );
  end component;

    signal \arbRegSMCurrentState[14]\, 
        \arbRegSMCurrentState[15]\, N_19, \N_165\, N_166, \N_164\, 
        \N_14_i\, hwdata10, m6, N_8, GND_net_1, VCC_net_1
         : std_logic;

    for all : COREAHBLITE_SLAVESTAGE_1
	Use entity work.COREAHBLITE_SLAVESTAGE_1(DEF_ARCH);
    for all : COREAHBLITE_MASTERSTAGE_2_1_0_1_0
	Use entity work.COREAHBLITE_MASTERSTAGE_2_1_0_1_0(DEF_ARCH);
begin 

    arbRegSMCurrentState(15) <= \arbRegSMCurrentState[15]\;
    arbRegSMCurrentState(14) <= \arbRegSMCurrentState[14]\;
    N_165 <= \N_165\;
    N_164 <= \N_164\;
    N_14_i <= \N_14_i\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    slavestage_0 : COREAHBLITE_SLAVESTAGE_1
      port map(
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        AHB_slave_dummy_0_mem_wdata(31) => 
        AHB_slave_dummy_0_mem_wdata(31), 
        AHB_slave_dummy_0_mem_wdata(30) => 
        AHB_slave_dummy_0_mem_wdata(30), 
        AHB_slave_dummy_0_mem_wdata(29) => 
        AHB_slave_dummy_0_mem_wdata(29), 
        AHB_slave_dummy_0_mem_wdata(28) => 
        AHB_slave_dummy_0_mem_wdata(28), 
        AHB_slave_dummy_0_mem_wdata(27) => 
        AHB_slave_dummy_0_mem_wdata(27), 
        AHB_slave_dummy_0_mem_wdata(26) => 
        AHB_slave_dummy_0_mem_wdata(26), 
        AHB_slave_dummy_0_mem_wdata(25) => 
        AHB_slave_dummy_0_mem_wdata(25), 
        AHB_slave_dummy_0_mem_wdata(24) => 
        AHB_slave_dummy_0_mem_wdata(24), 
        AHB_slave_dummy_0_mem_wdata(23) => 
        AHB_slave_dummy_0_mem_wdata(23), 
        AHB_slave_dummy_0_mem_wdata(22) => 
        AHB_slave_dummy_0_mem_wdata(22), 
        AHB_slave_dummy_0_mem_wdata(21) => 
        AHB_slave_dummy_0_mem_wdata(21), 
        AHB_slave_dummy_0_mem_wdata(20) => 
        AHB_slave_dummy_0_mem_wdata(20), 
        AHB_slave_dummy_0_mem_wdata(19) => 
        AHB_slave_dummy_0_mem_wdata(19), 
        AHB_slave_dummy_0_mem_wdata(18) => 
        AHB_slave_dummy_0_mem_wdata(18), 
        AHB_slave_dummy_0_mem_wdata(17) => 
        AHB_slave_dummy_0_mem_wdata(17), 
        AHB_slave_dummy_0_mem_wdata(16) => 
        AHB_slave_dummy_0_mem_wdata(16), 
        AHB_slave_dummy_0_mem_wdata(15) => 
        AHB_slave_dummy_0_mem_wdata(15), 
        AHB_slave_dummy_0_mem_wdata(14) => 
        AHB_slave_dummy_0_mem_wdata(14), 
        AHB_slave_dummy_0_mem_wdata(13) => 
        AHB_slave_dummy_0_mem_wdata(13), 
        AHB_slave_dummy_0_mem_wdata(12) => 
        AHB_slave_dummy_0_mem_wdata(12), 
        AHB_slave_dummy_0_mem_wdata(11) => 
        AHB_slave_dummy_0_mem_wdata(11), 
        AHB_slave_dummy_0_mem_wdata(10) => 
        AHB_slave_dummy_0_mem_wdata(10), 
        AHB_slave_dummy_0_mem_wdata(9) => 
        AHB_slave_dummy_0_mem_wdata(9), 
        AHB_slave_dummy_0_mem_wdata(8) => 
        AHB_slave_dummy_0_mem_wdata(8), 
        AHB_slave_dummy_0_mem_wdata(7) => 
        AHB_slave_dummy_0_mem_wdata(7), 
        AHB_slave_dummy_0_mem_wdata(6) => 
        AHB_slave_dummy_0_mem_wdata(6), 
        AHB_slave_dummy_0_mem_wdata(5) => 
        AHB_slave_dummy_0_mem_wdata(5), 
        AHB_slave_dummy_0_mem_wdata(4) => 
        AHB_slave_dummy_0_mem_wdata(4), 
        AHB_slave_dummy_0_mem_wdata(3) => 
        AHB_slave_dummy_0_mem_wdata(3), 
        AHB_slave_dummy_0_mem_wdata(2) => 
        AHB_slave_dummy_0_mem_wdata(2), 
        AHB_slave_dummy_0_mem_wdata(1) => 
        AHB_slave_dummy_0_mem_wdata(1), 
        AHB_slave_dummy_0_mem_wdata(0) => 
        AHB_slave_dummy_0_mem_wdata(0), arbRegSMCurrentState(15)
         => \arbRegSMCurrentState[15]\, arbRegSMCurrentState(14)
         => \arbRegSMCurrentState[14]\, hwdata10 => hwdata10, 
        MSS_READY => MSS_READY, sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, N_14_i => 
        \N_14_i\, N_19 => N_19, N_165 => \N_165\, m6 => m6, N_164
         => \N_164\, N_166 => N_166, N_8 => N_8);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    masterstage_0 : COREAHBLITE_MASTERSTAGE_2_1_0_1_0
      port map(
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        arbRegSMCurrentState(15) => \arbRegSMCurrentState[15]\, 
        arbRegSMCurrentState(14) => \arbRegSMCurrentState[14]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        result_addr_net_0_0 => result_addr_net_0_0, 
        result_addr_net_0_3 => result_addr_net_0_3, MSS_READY => 
        MSS_READY, sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, N_19 => N_19, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        regHTRANS => regHTRANS, masterRegAddrSel => 
        masterRegAddrSel, N_165 => \N_165\, N_166 => N_166, N_164
         => \N_164\, N_114 => N_114, N_115 => N_115, N_116 => 
        N_116, N_117 => N_117, N_118 => N_118, N_119 => N_119, 
        N_14_i => \N_14_i\, hready_m_xhdl339 => hready_m_xhdl339, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, hwdata10 => 
        hwdata10, ren_pos => ren_pos, N_273 => N_273, m6 => m6, 
        N_274 => N_274, N_59 => N_59, N_8 => N_8, N_31 => N_31, 
        defSlaveSMCurrentState => defSlaveSMCurrentState, 
        N_23_i_0 => N_23_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLite is

    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1);
          arbRegSMCurrentState                                 : out   std_logic_vector(15 downto 14);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0);
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic;
          result_addr_net_0_0                                  : in    std_logic;
          result_addr_net_0_3                                  : in    std_logic;
          MSS_READY                                            : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic;
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_165                                                : out   std_logic;
          N_164                                                : out   std_logic;
          N_114                                                : out   std_logic;
          N_115                                                : out   std_logic;
          N_116                                                : out   std_logic;
          N_117                                                : out   std_logic;
          N_118                                                : out   std_logic;
          N_119                                                : out   std_logic;
          N_14_i                                               : out   std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic;
          ren_pos                                              : in    std_logic;
          N_273                                                : out   std_logic;
          N_274                                                : out   std_logic;
          N_59                                                 : out   std_logic;
          N_31                                                 : out   std_logic;
          defSlaveSMCurrentState                               : out   std_logic;
          N_23_i_0                                             : out   std_logic
        );

end CoreAHBLite;

architecture DEF_ARCH of CoreAHBLite is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MATRIX4X16
    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1) := (others => 'U');
          arbRegSMCurrentState                                 : out   std_logic_vector(15 downto 14);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0) := (others => 'U');
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic := 'U';
          result_addr_net_0_0                                  : in    std_logic := 'U';
          result_addr_net_0_3                                  : in    std_logic := 'U';
          MSS_READY                                            : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_165                                                : out   std_logic;
          N_164                                                : out   std_logic;
          N_114                                                : out   std_logic;
          N_115                                                : out   std_logic;
          N_116                                                : out   std_logic;
          N_117                                                : out   std_logic;
          N_118                                                : out   std_logic;
          N_119                                                : out   std_logic;
          N_14_i                                               : out   std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic := 'U';
          ren_pos                                              : in    std_logic := 'U';
          N_273                                                : out   std_logic;
          N_274                                                : out   std_logic;
          N_59                                                 : out   std_logic;
          N_31                                                 : out   std_logic;
          defSlaveSMCurrentState                               : out   std_logic;
          N_23_i_0                                             : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : COREAHBLITE_MATRIX4X16
	Use entity work.COREAHBLITE_MATRIX4X16(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    matrix4x16 : COREAHBLITE_MATRIX4X16
      port map(
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        arbRegSMCurrentState(15) => arbRegSMCurrentState(15), 
        arbRegSMCurrentState(14) => arbRegSMCurrentState(14), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        AHB_slave_dummy_0_mem_wdata(31) => 
        AHB_slave_dummy_0_mem_wdata(31), 
        AHB_slave_dummy_0_mem_wdata(30) => 
        AHB_slave_dummy_0_mem_wdata(30), 
        AHB_slave_dummy_0_mem_wdata(29) => 
        AHB_slave_dummy_0_mem_wdata(29), 
        AHB_slave_dummy_0_mem_wdata(28) => 
        AHB_slave_dummy_0_mem_wdata(28), 
        AHB_slave_dummy_0_mem_wdata(27) => 
        AHB_slave_dummy_0_mem_wdata(27), 
        AHB_slave_dummy_0_mem_wdata(26) => 
        AHB_slave_dummy_0_mem_wdata(26), 
        AHB_slave_dummy_0_mem_wdata(25) => 
        AHB_slave_dummy_0_mem_wdata(25), 
        AHB_slave_dummy_0_mem_wdata(24) => 
        AHB_slave_dummy_0_mem_wdata(24), 
        AHB_slave_dummy_0_mem_wdata(23) => 
        AHB_slave_dummy_0_mem_wdata(23), 
        AHB_slave_dummy_0_mem_wdata(22) => 
        AHB_slave_dummy_0_mem_wdata(22), 
        AHB_slave_dummy_0_mem_wdata(21) => 
        AHB_slave_dummy_0_mem_wdata(21), 
        AHB_slave_dummy_0_mem_wdata(20) => 
        AHB_slave_dummy_0_mem_wdata(20), 
        AHB_slave_dummy_0_mem_wdata(19) => 
        AHB_slave_dummy_0_mem_wdata(19), 
        AHB_slave_dummy_0_mem_wdata(18) => 
        AHB_slave_dummy_0_mem_wdata(18), 
        AHB_slave_dummy_0_mem_wdata(17) => 
        AHB_slave_dummy_0_mem_wdata(17), 
        AHB_slave_dummy_0_mem_wdata(16) => 
        AHB_slave_dummy_0_mem_wdata(16), 
        AHB_slave_dummy_0_mem_wdata(15) => 
        AHB_slave_dummy_0_mem_wdata(15), 
        AHB_slave_dummy_0_mem_wdata(14) => 
        AHB_slave_dummy_0_mem_wdata(14), 
        AHB_slave_dummy_0_mem_wdata(13) => 
        AHB_slave_dummy_0_mem_wdata(13), 
        AHB_slave_dummy_0_mem_wdata(12) => 
        AHB_slave_dummy_0_mem_wdata(12), 
        AHB_slave_dummy_0_mem_wdata(11) => 
        AHB_slave_dummy_0_mem_wdata(11), 
        AHB_slave_dummy_0_mem_wdata(10) => 
        AHB_slave_dummy_0_mem_wdata(10), 
        AHB_slave_dummy_0_mem_wdata(9) => 
        AHB_slave_dummy_0_mem_wdata(9), 
        AHB_slave_dummy_0_mem_wdata(8) => 
        AHB_slave_dummy_0_mem_wdata(8), 
        AHB_slave_dummy_0_mem_wdata(7) => 
        AHB_slave_dummy_0_mem_wdata(7), 
        AHB_slave_dummy_0_mem_wdata(6) => 
        AHB_slave_dummy_0_mem_wdata(6), 
        AHB_slave_dummy_0_mem_wdata(5) => 
        AHB_slave_dummy_0_mem_wdata(5), 
        AHB_slave_dummy_0_mem_wdata(4) => 
        AHB_slave_dummy_0_mem_wdata(4), 
        AHB_slave_dummy_0_mem_wdata(3) => 
        AHB_slave_dummy_0_mem_wdata(3), 
        AHB_slave_dummy_0_mem_wdata(2) => 
        AHB_slave_dummy_0_mem_wdata(2), 
        AHB_slave_dummy_0_mem_wdata(1) => 
        AHB_slave_dummy_0_mem_wdata(1), 
        AHB_slave_dummy_0_mem_wdata(0) => 
        AHB_slave_dummy_0_mem_wdata(0), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        result_addr_net_0_0 => result_addr_net_0_0, 
        result_addr_net_0_3 => result_addr_net_0_3, MSS_READY => 
        MSS_READY, sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        regHTRANS => regHTRANS, masterRegAddrSel => 
        masterRegAddrSel, N_165 => N_165, N_164 => N_164, N_114
         => N_114, N_115 => N_115, N_116 => N_116, N_117 => N_117, 
        N_118 => N_118, N_119 => N_119, N_14_i => N_14_i, 
        hready_m_xhdl339 => hready_m_xhdl339, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, ren_pos => 
        ren_pos, N_273 => N_273, N_274 => N_274, N_59 => N_59, 
        N_31 => N_31, defSlaveSMCurrentState => 
        defSlaveSMCurrentState, N_23_i_0 => N_23_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_system_sb_CCC_0_FCCC is

    port( sha256_system_sb_0_FIC_0_CLK                       : out   std_logic;
          FIC_0_LOCK                                         : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic
        );

end sha256_system_sb_CCC_0_FCCC;

architecture DEF_ARCH of sha256_system_sb_CCC_0_FCCC is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => sha256_system_sb_0_FIC_0_CLK);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007FB8000044D74000318C6318C1F18C61EC0404040400301",
         VCOFREQUENCY => 800.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => FIC_0_LOCK, 
        BUSY => OPEN, CLK0 => VCC_net_1, CLK1 => VCC_net_1, CLK2
         => VCC_net_1, CLK3 => VCC_net_1, NGMUX0_SEL => GND_net_1, 
        NGMUX1_SEL => GND_net_1, NGMUX2_SEL => GND_net_1, 
        NGMUX3_SEL => GND_net_1, NGMUX0_HOLD_N => VCC_net_1, 
        NGMUX1_HOLD_N => VCC_net_1, NGMUX2_HOLD_N => VCC_net_1, 
        NGMUX3_HOLD_N => VCC_net_1, NGMUX0_ARST_N => VCC_net_1, 
        NGMUX1_ARST_N => VCC_net_1, NGMUX2_ARST_N => VCC_net_1, 
        NGMUX3_ARST_N => VCC_net_1, PLL_BYPASS_N => VCC_net_1, 
        PLL_ARST_N => VCC_net_1, PLL_POWERDOWN_N => VCC_net_1, 
        GPD0_ARST_N => VCC_net_1, GPD1_ARST_N => VCC_net_1, 
        GPD2_ARST_N => VCC_net_1, GPD3_ARST_N => VCC_net_1, 
        PRESET_N => GND_net_1, PCLK => VCC_net_1, PSEL => 
        VCC_net_1, PENABLE => VCC_net_1, PWRITE => VCC_net_1, 
        PADDR(7) => VCC_net_1, PADDR(6) => VCC_net_1, PADDR(5)
         => VCC_net_1, PADDR(4) => VCC_net_1, PADDR(3) => 
        VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7) => VCC_net_1, 
        PWDATA(6) => VCC_net_1, PWDATA(5) => VCC_net_1, PWDATA(4)
         => VCC_net_1, PWDATA(3) => VCC_net_1, PWDATA(2) => 
        VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0) => VCC_net_1, 
        CLK0_PAD => GND_net_1, CLK1_PAD => GND_net_1, CLK2_PAD
         => GND_net_1, CLK3_PAD => GND_net_1, GL0 => GL0_net, GL1
         => OPEN, GL2 => OPEN, GL3 => OPEN, RCOSC_25_50MHZ => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        RCOSC_1MHZ => GND_net_1, XTLOSC => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_system_sb is

    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : inout std_logic_vector(1 to 1) := (others => 'Z');
          arbRegSMCurrentState                                 : out   std_logic_vector(15 downto 14);
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          result_addr_net_0                                    : in    std_logic_vector(3 downto 0);
          state_out_net_0                                      : in    std_logic_vector(0 to 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : inout std_logic := 'Z';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : inout std_logic := 'Z';
          line_4_d0                                            : in    std_logic;
          line_21                                              : in    std_logic;
          line_3_d0                                            : in    std_logic;
          line_13                                              : in    std_logic;
          line_0_d0                                            : in    std_logic;
          line_24                                              : in    std_logic;
          line_0_4                                             : in    std_logic;
          line_0_21                                            : in    std_logic;
          line_0_3                                             : in    std_logic;
          line_0_13                                            : in    std_logic;
          line_0_0                                             : in    std_logic;
          line_0_24                                            : in    std_logic;
          line_1_4                                             : in    std_logic;
          line_1_21                                            : in    std_logic;
          line_1_3                                             : in    std_logic;
          line_1_13                                            : in    std_logic;
          line_1_0                                             : in    std_logic;
          line_1_24                                            : in    std_logic;
          line_2_4                                             : in    std_logic;
          line_2_21                                            : in    std_logic;
          line_2_3                                             : in    std_logic;
          line_2_13                                            : in    std_logic;
          line_2_0                                             : in    std_logic;
          line_2_24                                            : in    std_logic;
          line_3_3                                             : in    std_logic;
          line_3_21                                            : in    std_logic;
          line_3_0                                             : in    std_logic;
          line_3_4                                             : in    std_logic;
          line_3_24                                            : in    std_logic;
          line_3_13                                            : in    std_logic;
          line_4_3                                             : in    std_logic;
          line_4_21                                            : in    std_logic;
          line_4_0                                             : in    std_logic;
          line_4_4                                             : in    std_logic;
          line_4_24                                            : in    std_logic;
          line_4_13                                            : in    std_logic;
          line_5_3                                             : in    std_logic;
          line_5_21                                            : in    std_logic;
          line_5_0                                             : in    std_logic;
          line_5_4                                             : in    std_logic;
          line_5_24                                            : in    std_logic;
          line_5_13                                            : in    std_logic;
          line_6_3                                             : in    std_logic;
          line_6_21                                            : in    std_logic;
          line_6_0                                             : in    std_logic;
          line_6_4                                             : in    std_logic;
          line_6_24                                            : in    std_logic;
          line_6_13                                            : in    std_logic;
          line_7_3                                             : in    std_logic;
          line_7_0                                             : in    std_logic;
          line_7_13                                            : in    std_logic;
          line_7_4                                             : in    std_logic;
          line_7_21                                            : in    std_logic;
          sha256_system_sb_0_POWER_ON_RESET_N                  : out   std_logic;
          DEVRST_N                                             : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : out   std_logic;
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_165                                                : out   std_logic;
          N_164                                                : out   std_logic;
          N_114                                                : out   std_logic;
          N_115                                                : out   std_logic;
          N_116                                                : out   std_logic;
          N_117                                                : out   std_logic;
          N_118                                                : out   std_logic;
          N_119                                                : out   std_logic;
          N_14_i                                               : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic;
          ren_pos                                              : in    std_logic;
          N_31                                                 : out   std_logic;
          defSlaveSMCurrentState                               : out   std_logic;
          N_96                                                 : in    std_logic;
          N_516                                                : in    std_logic;
          N_582                                                : in    std_logic;
          N_520                                                : in    std_logic;
          N_586                                                : in    std_logic;
          N_504                                                : in    std_logic;
          N_570                                                : in    std_logic;
          N_508                                                : in    std_logic;
          N_574                                                : in    std_logic;
          N_512                                                : in    std_logic;
          N_578                                                : in    std_logic;
          N_503                                                : in    std_logic;
          N_569                                                : in    std_logic;
          N_505                                                : in    std_logic;
          N_571                                                : in    std_logic;
          N_517                                                : in    std_logic;
          N_583                                                : in    std_logic;
          N_523                                                : in    std_logic;
          N_589                                                : in    std_logic;
          N_528                                                : in    std_logic;
          N_594                                                : in    std_logic;
          N_529                                                : in    std_logic;
          N_595                                                : in    std_logic;
          N_526                                                : in    std_logic;
          N_592                                                : in    std_logic;
          N_524                                                : in    std_logic;
          N_590                                                : in    std_logic;
          N_515                                                : in    std_logic;
          N_581                                                : in    std_logic;
          N_514                                                : in    std_logic;
          N_580                                                : in    std_logic;
          N_522                                                : in    std_logic;
          N_588                                                : in    std_logic;
          N_502                                                : in    std_logic;
          N_568                                                : in    std_logic;
          N_513                                                : in    std_logic;
          N_579                                                : in    std_logic;
          N_525                                                : in    std_logic;
          N_591                                                : in    std_logic;
          N_500                                                : in    std_logic;
          N_566                                                : in    std_logic;
          N_501                                                : in    std_logic;
          N_567                                                : in    std_logic;
          N_499                                                : in    std_logic;
          N_565                                                : in    std_logic;
          N_74                                                 : in    std_logic;
          N_228                                                : in    std_logic;
          N_81                                                 : in    std_logic;
          N_7                                                  : in    std_logic;
          N_75                                                 : in    std_logic;
          sha256_system_sb_0_GPIO_1_M2F                        : out   std_logic;
          GPIO_0_M2F_c                                         : out   std_logic;
          sha256_system_sb_0_GPIO_9_M2F                        : out   std_logic;
          N_87_i_0                                             : in    std_logic;
          N_88_i_0                                             : in    std_logic;
          ce_i_i_2_i_0                                         : in    std_logic;
          SHA256_Module_0_data_available_lastbank_8            : in    std_logic;
          SHA256_Module_0_di_req_o                             : in    std_logic;
          SHA256_Module_0_data_out_ready                       : in    std_logic;
          SHA256_Module_0_do_valid_o                           : in    std_logic;
          SHA256_Module_0_data_available                       : in    std_logic;
          SHA256_Module_0_error_o                              : in    std_logic
        );

end sha256_system_sb;

architecture DEF_ARCH of sha256_system_sb is 

  component sha256_system_sb_MSS
    port( result_addr_net_0                                    : in    std_logic_vector(2 downto 0) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : out   std_logic_vector(1 to 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : out   std_logic_vector(31 downto 0);
          state_out_net_0                                      : in    std_logic_vector(0 to 0) := (others => 'U');
          line_4_d0                                            : in    std_logic := 'U';
          line_21                                              : in    std_logic := 'U';
          line_3_d0                                            : in    std_logic := 'U';
          line_13                                              : in    std_logic := 'U';
          line_0_d0                                            : in    std_logic := 'U';
          line_24                                              : in    std_logic := 'U';
          line_0_4                                             : in    std_logic := 'U';
          line_0_21                                            : in    std_logic := 'U';
          line_0_3                                             : in    std_logic := 'U';
          line_0_13                                            : in    std_logic := 'U';
          line_0_0                                             : in    std_logic := 'U';
          line_0_24                                            : in    std_logic := 'U';
          line_1_4                                             : in    std_logic := 'U';
          line_1_21                                            : in    std_logic := 'U';
          line_1_3                                             : in    std_logic := 'U';
          line_1_13                                            : in    std_logic := 'U';
          line_1_0                                             : in    std_logic := 'U';
          line_1_24                                            : in    std_logic := 'U';
          line_2_4                                             : in    std_logic := 'U';
          line_2_21                                            : in    std_logic := 'U';
          line_2_3                                             : in    std_logic := 'U';
          line_2_13                                            : in    std_logic := 'U';
          line_2_0                                             : in    std_logic := 'U';
          line_2_24                                            : in    std_logic := 'U';
          line_3_3                                             : in    std_logic := 'U';
          line_3_21                                            : in    std_logic := 'U';
          line_3_0                                             : in    std_logic := 'U';
          line_3_4                                             : in    std_logic := 'U';
          line_3_24                                            : in    std_logic := 'U';
          line_3_13                                            : in    std_logic := 'U';
          line_4_3                                             : in    std_logic := 'U';
          line_4_21                                            : in    std_logic := 'U';
          line_4_0                                             : in    std_logic := 'U';
          line_4_4                                             : in    std_logic := 'U';
          line_4_24                                            : in    std_logic := 'U';
          line_4_13                                            : in    std_logic := 'U';
          line_5_3                                             : in    std_logic := 'U';
          line_5_21                                            : in    std_logic := 'U';
          line_5_0                                             : in    std_logic := 'U';
          line_5_4                                             : in    std_logic := 'U';
          line_5_24                                            : in    std_logic := 'U';
          line_5_13                                            : in    std_logic := 'U';
          line_6_3                                             : in    std_logic := 'U';
          line_6_21                                            : in    std_logic := 'U';
          line_6_0                                             : in    std_logic := 'U';
          line_6_4                                             : in    std_logic := 'U';
          line_6_24                                            : in    std_logic := 'U';
          line_6_13                                            : in    std_logic := 'U';
          line_7_3                                             : in    std_logic := 'U';
          line_7_0                                             : in    std_logic := 'U';
          line_7_13                                            : in    std_logic := 'U';
          line_7_4                                             : in    std_logic := 'U';
          line_7_21                                            : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_26 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_27 : out   std_logic;
          N_96                                                 : in    std_logic := 'U';
          hready_m_xhdl339                                     : in    std_logic := 'U';
          ren_pos                                              : in    std_logic := 'U';
          N_516                                                : in    std_logic := 'U';
          N_582                                                : in    std_logic := 'U';
          N_520                                                : in    std_logic := 'U';
          N_586                                                : in    std_logic := 'U';
          N_504                                                : in    std_logic := 'U';
          N_570                                                : in    std_logic := 'U';
          N_508                                                : in    std_logic := 'U';
          N_574                                                : in    std_logic := 'U';
          N_512                                                : in    std_logic := 'U';
          N_578                                                : in    std_logic := 'U';
          N_503                                                : in    std_logic := 'U';
          N_569                                                : in    std_logic := 'U';
          N_505                                                : in    std_logic := 'U';
          N_571                                                : in    std_logic := 'U';
          N_517                                                : in    std_logic := 'U';
          N_583                                                : in    std_logic := 'U';
          N_523                                                : in    std_logic := 'U';
          N_589                                                : in    std_logic := 'U';
          N_528                                                : in    std_logic := 'U';
          N_594                                                : in    std_logic := 'U';
          N_529                                                : in    std_logic := 'U';
          N_595                                                : in    std_logic := 'U';
          N_526                                                : in    std_logic := 'U';
          N_592                                                : in    std_logic := 'U';
          N_524                                                : in    std_logic := 'U';
          N_590                                                : in    std_logic := 'U';
          N_515                                                : in    std_logic := 'U';
          N_581                                                : in    std_logic := 'U';
          N_514                                                : in    std_logic := 'U';
          N_580                                                : in    std_logic := 'U';
          N_522                                                : in    std_logic := 'U';
          N_588                                                : in    std_logic := 'U';
          N_502                                                : in    std_logic := 'U';
          N_568                                                : in    std_logic := 'U';
          N_513                                                : in    std_logic := 'U';
          N_579                                                : in    std_logic := 'U';
          N_525                                                : in    std_logic := 'U';
          N_591                                                : in    std_logic := 'U';
          N_500                                                : in    std_logic := 'U';
          N_566                                                : in    std_logic := 'U';
          N_501                                                : in    std_logic := 'U';
          N_567                                                : in    std_logic := 'U';
          N_499                                                : in    std_logic := 'U';
          N_565                                                : in    std_logic := 'U';
          N_74                                                 : in    std_logic := 'U';
          N_228                                                : in    std_logic := 'U';
          N_81                                                 : in    std_logic := 'U';
          N_7                                                  : in    std_logic := 'U';
          N_75                                                 : in    std_logic := 'U';
          N_274                                                : in    std_logic := 'U';
          N_273                                                : in    std_logic := 'U';
          N_59                                                 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N      : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : out   std_logic;
          sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F           : out   std_logic;
          sha256_system_sb_0_GPIO_1_M2F                        : out   std_logic;
          GPIO_0_M2F_c                                         : out   std_logic;
          sha256_system_sb_0_GPIO_9_M2F                        : out   std_logic;
          N_23_i_0                                             : in    std_logic := 'U';
          N_31                                                 : in    std_logic := 'U';
          FIC_0_LOCK                                           : in    std_logic := 'U';
          N_87_i_0                                             : in    std_logic := 'U';
          N_88_i_0                                             : in    std_logic := 'U';
          ce_i_i_2_i_0                                         : in    std_logic := 'U';
          SHA256_Module_0_data_available_lastbank_8            : in    std_logic := 'U';
          SHA256_Module_0_di_req_o                             : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready                       : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o                           : in    std_logic := 'U';
          SHA256_Module_0_data_available                       : in    std_logic := 'U';
          SHA256_Module_0_error_o                              : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic := 'U'
        );
  end component;

  component sha256_system_sb_FABOSC_0_OSC
    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );
  end component;

  component CoreResetP
    port( MSS_READY                                       : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK                    : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic := 'U';
          sha256_system_sb_0_POWER_ON_RESET_N             : in    std_logic := 'U'
        );
  end component;

  component CoreAHBLite
    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1) := (others => 'U');
          arbRegSMCurrentState                                 : out   std_logic_vector(15 downto 14);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0) := (others => 'U');
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic := 'U';
          result_addr_net_0_0                                  : in    std_logic := 'U';
          result_addr_net_0_3                                  : in    std_logic := 'U';
          MSS_READY                                            : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_165                                                : out   std_logic;
          N_164                                                : out   std_logic;
          N_114                                                : out   std_logic;
          N_115                                                : out   std_logic;
          N_116                                                : out   std_logic;
          N_117                                                : out   std_logic;
          N_118                                                : out   std_logic;
          N_119                                                : out   std_logic;
          N_14_i                                               : out   std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic := 'U';
          ren_pos                                              : in    std_logic := 'U';
          N_273                                                : out   std_logic;
          N_274                                                : out   std_logic;
          N_59                                                 : out   std_logic;
          N_31                                                 : out   std_logic;
          defSlaveSMCurrentState                               : out   std_logic;
          N_23_i_0                                             : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component sha256_system_sb_CCC_0_FCCC
    port( sha256_system_sb_0_FIC_0_CLK                       : out   std_logic;
          FIC_0_LOCK                                         : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

    signal \sha256_system_sb_0_POWER_ON_RESET_N\, \SYSRESET_POR\, 
        \sha256_system_sb_0_FIC_0_CLK\, FIC_0_LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[6]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[26]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[27]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        MSS_READY, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        hready_m_xhdl339, N_273, N_274, N_59, \N_31\, N_23_i_0, 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        GND_net_1, VCC_net_1 : std_logic;

    for all : sha256_system_sb_MSS
	Use entity work.sha256_system_sb_MSS(DEF_ARCH);
    for all : sha256_system_sb_FABOSC_0_OSC
	Use entity work.sha256_system_sb_FABOSC_0_OSC(DEF_ARCH);
    for all : CoreResetP
	Use entity work.CoreResetP(DEF_ARCH);
    for all : CoreAHBLite
	Use entity work.CoreAHBLite(DEF_ARCH);
    for all : sha256_system_sb_CCC_0_FCCC
	Use entity work.sha256_system_sb_CCC_0_FCCC(DEF_ARCH);
begin 

    sha256_system_sb_0_POWER_ON_RESET_N <= 
        \sha256_system_sb_0_POWER_ON_RESET_N\;
    sha256_system_sb_0_FIC_0_CLK <= 
        \sha256_system_sb_0_FIC_0_CLK\;
    N_31 <= \N_31\;

    sha256_system_sb_MSS_0 : sha256_system_sb_MSS
      port map(result_addr_net_0(2) => result_addr_net_0(2), 
        result_addr_net_0(1) => result_addr_net_0(1), 
        result_addr_net_0(0) => result_addr_net_0(0), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        state_out_net_0(0) => state_out_net_0(0), line_4_d0 => 
        line_4_d0, line_21 => line_21, line_3_d0 => line_3_d0, 
        line_13 => line_13, line_0_d0 => line_0_d0, line_24 => 
        line_24, line_0_4 => line_0_4, line_0_21 => line_0_21, 
        line_0_3 => line_0_3, line_0_13 => line_0_13, line_0_0
         => line_0_0, line_0_24 => line_0_24, line_1_4 => 
        line_1_4, line_1_21 => line_1_21, line_1_3 => line_1_3, 
        line_1_13 => line_1_13, line_1_0 => line_1_0, line_1_24
         => line_1_24, line_2_4 => line_2_4, line_2_21 => 
        line_2_21, line_2_3 => line_2_3, line_2_13 => line_2_13, 
        line_2_0 => line_2_0, line_2_24 => line_2_24, line_3_3
         => line_3_3, line_3_21 => line_3_21, line_3_0 => 
        line_3_0, line_3_4 => line_3_4, line_3_24 => line_3_24, 
        line_3_13 => line_3_13, line_4_3 => line_4_3, line_4_21
         => line_4_21, line_4_0 => line_4_0, line_4_4 => line_4_4, 
        line_4_24 => line_4_24, line_4_13 => line_4_13, line_5_3
         => line_5_3, line_5_21 => line_5_21, line_5_0 => 
        line_5_0, line_5_4 => line_5_4, line_5_24 => line_5_24, 
        line_5_13 => line_5_13, line_6_3 => line_6_3, line_6_21
         => line_6_21, line_6_0 => line_6_0, line_6_4 => line_6_4, 
        line_6_24 => line_6_24, line_6_13 => line_6_13, line_7_3
         => line_7_3, line_7_0 => line_7_0, line_7_13 => 
        line_7_13, line_7_4 => line_7_4, line_7_21 => line_7_21, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[6]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_26 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[26]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_27 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[27]\, 
        N_96 => N_96, hready_m_xhdl339 => hready_m_xhdl339, 
        ren_pos => ren_pos, N_516 => N_516, N_582 => N_582, N_520
         => N_520, N_586 => N_586, N_504 => N_504, N_570 => N_570, 
        N_508 => N_508, N_574 => N_574, N_512 => N_512, N_578 => 
        N_578, N_503 => N_503, N_569 => N_569, N_505 => N_505, 
        N_571 => N_571, N_517 => N_517, N_583 => N_583, N_523 => 
        N_523, N_589 => N_589, N_528 => N_528, N_594 => N_594, 
        N_529 => N_529, N_595 => N_595, N_526 => N_526, N_592 => 
        N_592, N_524 => N_524, N_590 => N_590, N_515 => N_515, 
        N_581 => N_581, N_514 => N_514, N_580 => N_580, N_522 => 
        N_522, N_588 => N_588, N_502 => N_502, N_568 => N_568, 
        N_513 => N_513, N_579 => N_579, N_525 => N_525, N_591 => 
        N_591, N_500 => N_500, N_566 => N_566, N_501 => N_501, 
        N_567 => N_567, N_499 => N_499, N_565 => N_565, N_74 => 
        N_74, N_228 => N_228, N_81 => N_81, N_7 => N_7, N_75 => 
        N_75, N_274 => N_274, N_273 => N_273, N_59 => N_59, 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        sha256_system_sb_0_GPIO_1_M2F => 
        sha256_system_sb_0_GPIO_1_M2F, GPIO_0_M2F_c => 
        GPIO_0_M2F_c, sha256_system_sb_0_GPIO_9_M2F => 
        sha256_system_sb_0_GPIO_9_M2F, N_23_i_0 => N_23_i_0, N_31
         => \N_31\, FIC_0_LOCK => FIC_0_LOCK, N_87_i_0 => 
        N_87_i_0, N_88_i_0 => N_88_i_0, ce_i_i_2_i_0 => 
        ce_i_i_2_i_0, SHA256_Module_0_data_available_lastbank_8
         => SHA256_Module_0_data_available_lastbank_8, 
        SHA256_Module_0_di_req_o => SHA256_Module_0_di_req_o, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready, 
        SHA256_Module_0_do_valid_o => SHA256_Module_0_do_valid_o, 
        SHA256_Module_0_data_available => 
        SHA256_Module_0_data_available, SHA256_Module_0_error_o
         => SHA256_Module_0_error_o, sha256_system_sb_0_FIC_0_CLK
         => \sha256_system_sb_0_FIC_0_CLK\);
    
    FABOSC_0 : sha256_system_sb_FABOSC_0_OSC
      port map(FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
         => FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    CORERESETP_0 : CoreResetP
      port map(MSS_READY => MSS_READY, 
        sha256_system_sb_0_FIC_0_CLK => 
        \sha256_system_sb_0_FIC_0_CLK\, 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        sha256_system_sb_0_POWER_ON_RESET_N => 
        \sha256_system_sb_0_POWER_ON_RESET_N\);
    
    CoreAHBLite_0 : CoreAHBLite
      port map(
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        arbRegSMCurrentState(15) => arbRegSMCurrentState(15), 
        arbRegSMCurrentState(14) => arbRegSMCurrentState(14), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        AHB_slave_dummy_0_mem_wdata(31) => 
        AHB_slave_dummy_0_mem_wdata(31), 
        AHB_slave_dummy_0_mem_wdata(30) => 
        AHB_slave_dummy_0_mem_wdata(30), 
        AHB_slave_dummy_0_mem_wdata(29) => 
        AHB_slave_dummy_0_mem_wdata(29), 
        AHB_slave_dummy_0_mem_wdata(28) => 
        AHB_slave_dummy_0_mem_wdata(28), 
        AHB_slave_dummy_0_mem_wdata(27) => 
        AHB_slave_dummy_0_mem_wdata(27), 
        AHB_slave_dummy_0_mem_wdata(26) => 
        AHB_slave_dummy_0_mem_wdata(26), 
        AHB_slave_dummy_0_mem_wdata(25) => 
        AHB_slave_dummy_0_mem_wdata(25), 
        AHB_slave_dummy_0_mem_wdata(24) => 
        AHB_slave_dummy_0_mem_wdata(24), 
        AHB_slave_dummy_0_mem_wdata(23) => 
        AHB_slave_dummy_0_mem_wdata(23), 
        AHB_slave_dummy_0_mem_wdata(22) => 
        AHB_slave_dummy_0_mem_wdata(22), 
        AHB_slave_dummy_0_mem_wdata(21) => 
        AHB_slave_dummy_0_mem_wdata(21), 
        AHB_slave_dummy_0_mem_wdata(20) => 
        AHB_slave_dummy_0_mem_wdata(20), 
        AHB_slave_dummy_0_mem_wdata(19) => 
        AHB_slave_dummy_0_mem_wdata(19), 
        AHB_slave_dummy_0_mem_wdata(18) => 
        AHB_slave_dummy_0_mem_wdata(18), 
        AHB_slave_dummy_0_mem_wdata(17) => 
        AHB_slave_dummy_0_mem_wdata(17), 
        AHB_slave_dummy_0_mem_wdata(16) => 
        AHB_slave_dummy_0_mem_wdata(16), 
        AHB_slave_dummy_0_mem_wdata(15) => 
        AHB_slave_dummy_0_mem_wdata(15), 
        AHB_slave_dummy_0_mem_wdata(14) => 
        AHB_slave_dummy_0_mem_wdata(14), 
        AHB_slave_dummy_0_mem_wdata(13) => 
        AHB_slave_dummy_0_mem_wdata(13), 
        AHB_slave_dummy_0_mem_wdata(12) => 
        AHB_slave_dummy_0_mem_wdata(12), 
        AHB_slave_dummy_0_mem_wdata(11) => 
        AHB_slave_dummy_0_mem_wdata(11), 
        AHB_slave_dummy_0_mem_wdata(10) => 
        AHB_slave_dummy_0_mem_wdata(10), 
        AHB_slave_dummy_0_mem_wdata(9) => 
        AHB_slave_dummy_0_mem_wdata(9), 
        AHB_slave_dummy_0_mem_wdata(8) => 
        AHB_slave_dummy_0_mem_wdata(8), 
        AHB_slave_dummy_0_mem_wdata(7) => 
        AHB_slave_dummy_0_mem_wdata(7), 
        AHB_slave_dummy_0_mem_wdata(6) => 
        AHB_slave_dummy_0_mem_wdata(6), 
        AHB_slave_dummy_0_mem_wdata(5) => 
        AHB_slave_dummy_0_mem_wdata(5), 
        AHB_slave_dummy_0_mem_wdata(4) => 
        AHB_slave_dummy_0_mem_wdata(4), 
        AHB_slave_dummy_0_mem_wdata(3) => 
        AHB_slave_dummy_0_mem_wdata(3), 
        AHB_slave_dummy_0_mem_wdata(2) => 
        AHB_slave_dummy_0_mem_wdata(2), 
        AHB_slave_dummy_0_mem_wdata(1) => 
        AHB_slave_dummy_0_mem_wdata(1), 
        AHB_slave_dummy_0_mem_wdata(0) => 
        AHB_slave_dummy_0_mem_wdata(0), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[6]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[26]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[27]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        result_addr_net_0_0 => result_addr_net_0(0), 
        result_addr_net_0_3 => result_addr_net_0(3), MSS_READY
         => MSS_READY, sha256_system_sb_0_FIC_0_CLK => 
        \sha256_system_sb_0_FIC_0_CLK\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        regHTRANS => regHTRANS, masterRegAddrSel => 
        masterRegAddrSel, N_165 => N_165, N_164 => N_164, N_114
         => N_114, N_115 => N_115, N_116 => N_116, N_117 => N_117, 
        N_118 => N_118, N_119 => N_119, N_14_i => N_14_i, 
        hready_m_xhdl339 => hready_m_xhdl339, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, ren_pos => 
        ren_pos, N_273 => N_273, N_274 => N_274, N_59 => N_59, 
        N_31 => \N_31\, defSlaveSMCurrentState => 
        defSlaveSMCurrentState, N_23_i_0 => N_23_i_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    SYSRESET_POR_RNI03O8 : CLKINT
      port map(A => \SYSRESET_POR\, Y => 
        \sha256_system_sb_0_POWER_ON_RESET_N\);
    
    CCC_0 : sha256_system_sb_CCC_0_FCCC
      port map(sha256_system_sb_0_FIC_0_CLK => 
        \sha256_system_sb_0_FIC_0_CLK\, FIC_0_LOCK => FIC_0_LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => \SYSRESET_POR\, DEVRST_N => 
        DEVRST_N);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_system is

    port( DEVRST_N   : in    std_logic;
          GPIO_0_M2F : out   std_logic
        );

end sha256_system;

architecture DEF_ARCH of sha256_system is 

  component SHA256_Module
    port( result_addr_net_0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          AHB_slave_dummy_0_mem_wdata               : in    std_logic_vector(31 downto 0) := (others => 'U');
          waddr_in_net_0                            : in    std_logic_vector(4 downto 0) := (others => 'U');
          state_out_net_0                           : out   std_logic_vector(0 to 0);
          line_0_d0                                 : out   std_logic;
          line_3_d0                                 : out   std_logic;
          line_4_d0                                 : out   std_logic;
          line_13                                   : out   std_logic;
          line_21                                   : out   std_logic;
          line_24                                   : out   std_logic;
          line_0_0                                  : out   std_logic;
          line_0_3                                  : out   std_logic;
          line_0_4                                  : out   std_logic;
          line_0_13                                 : out   std_logic;
          line_0_21                                 : out   std_logic;
          line_0_24                                 : out   std_logic;
          line_1_0                                  : out   std_logic;
          line_1_3                                  : out   std_logic;
          line_1_4                                  : out   std_logic;
          line_1_13                                 : out   std_logic;
          line_1_21                                 : out   std_logic;
          line_1_24                                 : out   std_logic;
          line_2_0                                  : out   std_logic;
          line_2_3                                  : out   std_logic;
          line_2_4                                  : out   std_logic;
          line_2_13                                 : out   std_logic;
          line_2_21                                 : out   std_logic;
          line_2_24                                 : out   std_logic;
          line_3_0                                  : out   std_logic;
          line_3_3                                  : out   std_logic;
          line_3_4                                  : out   std_logic;
          line_3_13                                 : out   std_logic;
          line_3_21                                 : out   std_logic;
          line_3_24                                 : out   std_logic;
          line_4_0                                  : out   std_logic;
          line_4_3                                  : out   std_logic;
          line_4_4                                  : out   std_logic;
          line_4_13                                 : out   std_logic;
          line_4_21                                 : out   std_logic;
          line_4_24                                 : out   std_logic;
          line_5_0                                  : out   std_logic;
          line_5_3                                  : out   std_logic;
          line_5_4                                  : out   std_logic;
          line_5_13                                 : out   std_logic;
          line_5_21                                 : out   std_logic;
          line_5_24                                 : out   std_logic;
          line_6_0                                  : out   std_logic;
          line_6_3                                  : out   std_logic;
          line_6_4                                  : out   std_logic;
          line_6_13                                 : out   std_logic;
          line_6_21                                 : out   std_logic;
          line_6_24                                 : out   std_logic;
          line_7_21                                 : out   std_logic;
          line_7_13                                 : out   std_logic;
          line_7_4                                  : out   std_logic;
          line_7_3                                  : out   std_logic;
          line_7_0                                  : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK              : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o                : out   std_logic;
          N_568                                     : out   std_logic;
          N_579                                     : out   std_logic;
          N_580                                     : out   std_logic;
          N_581                                     : out   std_logic;
          N_583                                     : out   std_logic;
          N_588                                     : out   std_logic;
          N_589                                     : out   std_logic;
          N_590                                     : out   std_logic;
          N_591                                     : out   std_logic;
          N_592                                     : out   std_logic;
          N_595                                     : out   std_logic;
          N_594                                     : out   std_logic;
          N_586                                     : out   std_logic;
          N_582                                     : out   std_logic;
          N_578                                     : out   std_logic;
          N_574                                     : out   std_logic;
          N_571                                     : out   std_logic;
          N_570                                     : out   std_logic;
          N_569                                     : out   std_logic;
          N_96                                      : out   std_logic;
          N_81                                      : out   std_logic;
          N_74                                      : out   std_logic;
          N_75                                      : out   std_logic;
          N_499                                     : out   std_logic;
          N_501                                     : out   std_logic;
          N_525                                     : out   std_logic;
          N_513                                     : out   std_logic;
          N_502                                     : out   std_logic;
          N_522                                     : out   std_logic;
          N_500                                     : out   std_logic;
          N_514                                     : out   std_logic;
          N_515                                     : out   std_logic;
          N_524                                     : out   std_logic;
          N_526                                     : out   std_logic;
          N_529                                     : out   std_logic;
          N_528                                     : out   std_logic;
          N_523                                     : out   std_logic;
          N_517                                     : out   std_logic;
          N_505                                     : out   std_logic;
          N_503                                     : out   std_logic;
          N_512                                     : out   std_logic;
          N_508                                     : out   std_logic;
          N_504                                     : out   std_logic;
          N_520                                     : out   std_logic;
          N_516                                     : out   std_logic;
          ren_pos                                   : out   std_logic;
          N_228                                     : out   std_logic;
          N_7                                       : out   std_logic;
          N_566                                     : out   std_logic;
          N_567                                     : out   std_logic;
          N_565                                     : out   std_logic;
          SHA256_Module_0_data_out_ready            : out   std_logic;
          AHB_slave_dummy_0_read_en                 : in    std_logic := 'U';
          SHA256_Module_0_error_o                   : out   std_logic;
          SHA256_Module_0_di_req_o                  : out   std_logic;
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic;
          sha256_system_sb_0_GPIO_9_M2F             : in    std_logic := 'U';
          SHA256_Module_0_data_available            : out   std_logic;
          sha256_system_sb_0_GPIO_1_M2F             : in    std_logic := 'U';
          AHB_slave_dummy_0_write_en                : in    std_logic := 'U';
          ce_i_i_2_i_0                              : out   std_logic;
          N_88_i_0                                  : out   std_logic;
          N_87_i_0                                  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AHB_slave_dummy
    port( waddr_in_net_0                                     : out   std_logic_vector(4 downto 0);
          result_addr_net_0                                  : out   std_logic_vector(3 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS : in    std_logic_vector(1 to 1) := (others => 'U');
          arbRegSMCurrentState                               : in    std_logic_vector(15 downto 14) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR  : in    std_logic_vector(25 downto 24) := (others => 'U');
          sha256_system_sb_0_POWER_ON_RESET_N                : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                       : in    std_logic := 'U';
          N_118                                              : in    std_logic := 'U';
          N_117                                              : in    std_logic := 'U';
          N_116                                              : in    std_logic := 'U';
          N_115                                              : in    std_logic := 'U';
          N_114                                              : in    std_logic := 'U';
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY             : out   std_logic;
          AHB_slave_dummy_0_write_en                         : out   std_logic;
          AHB_slave_dummy_0_read_en                          : out   std_logic;
          N_119                                              : in    std_logic := 'U';
          masterRegAddrSel                                   : in    std_logic := 'U';
          regHTRANS                                          : in    std_logic := 'U';
          N_165                                              : in    std_logic := 'U';
          N_14_i                                             : in    std_logic := 'U';
          N_164                                              : in    std_logic := 'U';
          defSlaveSMCurrentState                             : in    std_logic := 'U';
          N_31                                               : in    std_logic := 'U'
        );
  end component;

  component sha256_system_sb
    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : inout   std_logic_vector(1 to 1);
          arbRegSMCurrentState                                 : out   std_logic_vector(15 downto 14);
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          result_addr_net_0                                    : in    std_logic_vector(3 downto 0) := (others => 'U');
          state_out_net_0                                      : in    std_logic_vector(0 to 0) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : inout   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : inout   std_logic;
          line_4_d0                                            : in    std_logic := 'U';
          line_21                                              : in    std_logic := 'U';
          line_3_d0                                            : in    std_logic := 'U';
          line_13                                              : in    std_logic := 'U';
          line_0_d0                                            : in    std_logic := 'U';
          line_24                                              : in    std_logic := 'U';
          line_0_4                                             : in    std_logic := 'U';
          line_0_21                                            : in    std_logic := 'U';
          line_0_3                                             : in    std_logic := 'U';
          line_0_13                                            : in    std_logic := 'U';
          line_0_0                                             : in    std_logic := 'U';
          line_0_24                                            : in    std_logic := 'U';
          line_1_4                                             : in    std_logic := 'U';
          line_1_21                                            : in    std_logic := 'U';
          line_1_3                                             : in    std_logic := 'U';
          line_1_13                                            : in    std_logic := 'U';
          line_1_0                                             : in    std_logic := 'U';
          line_1_24                                            : in    std_logic := 'U';
          line_2_4                                             : in    std_logic := 'U';
          line_2_21                                            : in    std_logic := 'U';
          line_2_3                                             : in    std_logic := 'U';
          line_2_13                                            : in    std_logic := 'U';
          line_2_0                                             : in    std_logic := 'U';
          line_2_24                                            : in    std_logic := 'U';
          line_3_3                                             : in    std_logic := 'U';
          line_3_21                                            : in    std_logic := 'U';
          line_3_0                                             : in    std_logic := 'U';
          line_3_4                                             : in    std_logic := 'U';
          line_3_24                                            : in    std_logic := 'U';
          line_3_13                                            : in    std_logic := 'U';
          line_4_3                                             : in    std_logic := 'U';
          line_4_21                                            : in    std_logic := 'U';
          line_4_0                                             : in    std_logic := 'U';
          line_4_4                                             : in    std_logic := 'U';
          line_4_24                                            : in    std_logic := 'U';
          line_4_13                                            : in    std_logic := 'U';
          line_5_3                                             : in    std_logic := 'U';
          line_5_21                                            : in    std_logic := 'U';
          line_5_0                                             : in    std_logic := 'U';
          line_5_4                                             : in    std_logic := 'U';
          line_5_24                                            : in    std_logic := 'U';
          line_5_13                                            : in    std_logic := 'U';
          line_6_3                                             : in    std_logic := 'U';
          line_6_21                                            : in    std_logic := 'U';
          line_6_0                                             : in    std_logic := 'U';
          line_6_4                                             : in    std_logic := 'U';
          line_6_24                                            : in    std_logic := 'U';
          line_6_13                                            : in    std_logic := 'U';
          line_7_3                                             : in    std_logic := 'U';
          line_7_0                                             : in    std_logic := 'U';
          line_7_13                                            : in    std_logic := 'U';
          line_7_4                                             : in    std_logic := 'U';
          line_7_21                                            : in    std_logic := 'U';
          sha256_system_sb_0_POWER_ON_RESET_N                  : out   std_logic;
          DEVRST_N                                             : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : out   std_logic;
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_165                                                : out   std_logic;
          N_164                                                : out   std_logic;
          N_114                                                : out   std_logic;
          N_115                                                : out   std_logic;
          N_116                                                : out   std_logic;
          N_117                                                : out   std_logic;
          N_118                                                : out   std_logic;
          N_119                                                : out   std_logic;
          N_14_i                                               : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic := 'U';
          ren_pos                                              : in    std_logic := 'U';
          N_31                                                 : out   std_logic;
          defSlaveSMCurrentState                               : out   std_logic;
          N_96                                                 : in    std_logic := 'U';
          N_516                                                : in    std_logic := 'U';
          N_582                                                : in    std_logic := 'U';
          N_520                                                : in    std_logic := 'U';
          N_586                                                : in    std_logic := 'U';
          N_504                                                : in    std_logic := 'U';
          N_570                                                : in    std_logic := 'U';
          N_508                                                : in    std_logic := 'U';
          N_574                                                : in    std_logic := 'U';
          N_512                                                : in    std_logic := 'U';
          N_578                                                : in    std_logic := 'U';
          N_503                                                : in    std_logic := 'U';
          N_569                                                : in    std_logic := 'U';
          N_505                                                : in    std_logic := 'U';
          N_571                                                : in    std_logic := 'U';
          N_517                                                : in    std_logic := 'U';
          N_583                                                : in    std_logic := 'U';
          N_523                                                : in    std_logic := 'U';
          N_589                                                : in    std_logic := 'U';
          N_528                                                : in    std_logic := 'U';
          N_594                                                : in    std_logic := 'U';
          N_529                                                : in    std_logic := 'U';
          N_595                                                : in    std_logic := 'U';
          N_526                                                : in    std_logic := 'U';
          N_592                                                : in    std_logic := 'U';
          N_524                                                : in    std_logic := 'U';
          N_590                                                : in    std_logic := 'U';
          N_515                                                : in    std_logic := 'U';
          N_581                                                : in    std_logic := 'U';
          N_514                                                : in    std_logic := 'U';
          N_580                                                : in    std_logic := 'U';
          N_522                                                : in    std_logic := 'U';
          N_588                                                : in    std_logic := 'U';
          N_502                                                : in    std_logic := 'U';
          N_568                                                : in    std_logic := 'U';
          N_513                                                : in    std_logic := 'U';
          N_579                                                : in    std_logic := 'U';
          N_525                                                : in    std_logic := 'U';
          N_591                                                : in    std_logic := 'U';
          N_500                                                : in    std_logic := 'U';
          N_566                                                : in    std_logic := 'U';
          N_501                                                : in    std_logic := 'U';
          N_567                                                : in    std_logic := 'U';
          N_499                                                : in    std_logic := 'U';
          N_565                                                : in    std_logic := 'U';
          N_74                                                 : in    std_logic := 'U';
          N_228                                                : in    std_logic := 'U';
          N_81                                                 : in    std_logic := 'U';
          N_7                                                  : in    std_logic := 'U';
          N_75                                                 : in    std_logic := 'U';
          sha256_system_sb_0_GPIO_1_M2F                        : out   std_logic;
          GPIO_0_M2F_c                                         : out   std_logic;
          sha256_system_sb_0_GPIO_9_M2F                        : out   std_logic;
          N_87_i_0                                             : in    std_logic := 'U';
          N_88_i_0                                             : in    std_logic := 'U';
          ce_i_i_2_i_0                                         : in    std_logic := 'U';
          SHA256_Module_0_data_available_lastbank_8            : in    std_logic := 'U';
          SHA256_Module_0_di_req_o                             : in    std_logic := 'U';
          SHA256_Module_0_data_out_ready                       : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o                           : in    std_logic := 'U';
          SHA256_Module_0_data_available                       : in    std_logic := 'U';
          SHA256_Module_0_error_o                              : in    std_logic := 'U'
        );
  end component;

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

    signal sha256_system_sb_0_FIC_0_CLK, 
        sha256_system_sb_0_POWER_ON_RESET_N, 
        \AHB_slave_dummy_0_mem_wdata[0]\, 
        \AHB_slave_dummy_0_mem_wdata[1]\, 
        \AHB_slave_dummy_0_mem_wdata[2]\, 
        \AHB_slave_dummy_0_mem_wdata[3]\, 
        \AHB_slave_dummy_0_mem_wdata[4]\, 
        \AHB_slave_dummy_0_mem_wdata[5]\, 
        \AHB_slave_dummy_0_mem_wdata[6]\, 
        \AHB_slave_dummy_0_mem_wdata[7]\, 
        \AHB_slave_dummy_0_mem_wdata[8]\, 
        \AHB_slave_dummy_0_mem_wdata[9]\, 
        \AHB_slave_dummy_0_mem_wdata[10]\, 
        \AHB_slave_dummy_0_mem_wdata[11]\, 
        \AHB_slave_dummy_0_mem_wdata[12]\, 
        \AHB_slave_dummy_0_mem_wdata[13]\, 
        \AHB_slave_dummy_0_mem_wdata[14]\, 
        \AHB_slave_dummy_0_mem_wdata[15]\, 
        \AHB_slave_dummy_0_mem_wdata[16]\, 
        \AHB_slave_dummy_0_mem_wdata[17]\, 
        \AHB_slave_dummy_0_mem_wdata[18]\, 
        \AHB_slave_dummy_0_mem_wdata[19]\, 
        \AHB_slave_dummy_0_mem_wdata[20]\, 
        \AHB_slave_dummy_0_mem_wdata[21]\, 
        \AHB_slave_dummy_0_mem_wdata[22]\, 
        \AHB_slave_dummy_0_mem_wdata[23]\, 
        \AHB_slave_dummy_0_mem_wdata[24]\, 
        \AHB_slave_dummy_0_mem_wdata[25]\, 
        \AHB_slave_dummy_0_mem_wdata[26]\, 
        \AHB_slave_dummy_0_mem_wdata[27]\, 
        \AHB_slave_dummy_0_mem_wdata[28]\, 
        \AHB_slave_dummy_0_mem_wdata[29]\, 
        \AHB_slave_dummy_0_mem_wdata[30]\, 
        \AHB_slave_dummy_0_mem_wdata[31]\, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, 
        \waddr_in_net_0[0]\, \waddr_in_net_0[1]\, 
        \waddr_in_net_0[2]\, \waddr_in_net_0[3]\, 
        \waddr_in_net_0[4]\, \result_addr_net_0[0]\, 
        \result_addr_net_0[1]\, \result_addr_net_0[2]\, 
        \result_addr_net_0[3]\, AHB_slave_dummy_0_write_en, 
        AHB_slave_dummy_0_read_en, sha256_system_sb_0_GPIO_9_M2F, 
        sha256_system_sb_0_GPIO_1_M2F, 
        SHA256_Module_0_data_available, 
        SHA256_Module_0_data_available_lastbank_8, 
        SHA256_Module_0_data_out_ready, 
        SHA256_Module_0_do_valid_o, SHA256_Module_0_error_o, 
        \state_out_net_0[0]\, GND_net_1, VCC_net_1, 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[24]\, 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[25]\, 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.masterRegAddrSel\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.regHTRANS\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.default_slave_sm.defSlaveSMCurrentState\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.slave_arbiter.arbRegSMCurrentState[15]\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.slave_arbiter.arbRegSMCurrentState[14]\, 
        N_14_i, \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.ren_pos\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[31]\, N_31, 
        N_96, N_7, N_228, N_81, N_74, N_75, 
        \SHA256_Module_0.reg9_1x32_0.N_565\, 
        \SHA256_Module_0.reg9_1x32_0.N_499\, 
        \SHA256_Module_0.reg9_1x32_0.N_567\, 
        \SHA256_Module_0.reg9_1x32_0.N_501\, 
        \SHA256_Module_0.reg9_1x32_0.N_591\, 
        \SHA256_Module_0.reg9_1x32_0.N_525\, 
        \SHA256_Module_0.reg9_1x32_0.N_579\, 
        \SHA256_Module_0.reg9_1x32_0.N_513\, 
        \SHA256_Module_0.reg9_1x32_0.N_568\, 
        \SHA256_Module_0.reg9_1x32_0.N_502\, 
        \SHA256_Module_0.reg9_1x32_0.N_522\, 
        \SHA256_Module_0.reg9_1x32_0.N_588\, 
        \SHA256_Module_0.reg9_1x32_0.N_583\, 
        \SHA256_Module_0.reg9_1x32_0.N_500\, 
        \SHA256_Module_0.reg9_1x32_0.N_514\, 
        \SHA256_Module_0.reg9_1x32_0.N_515\, 
        \SHA256_Module_0.reg9_1x32_0.N_524\, 
        \SHA256_Module_0.reg9_1x32_0.N_526\, 
        \SHA256_Module_0.reg9_1x32_0.N_529\, 
        \SHA256_Module_0.reg9_1x32_0.N_566\, 
        \SHA256_Module_0.reg9_1x32_0.N_580\, 
        \SHA256_Module_0.reg9_1x32_0.N_581\, 
        \SHA256_Module_0.reg9_1x32_0.N_590\, 
        \SHA256_Module_0.reg9_1x32_0.N_592\, 
        \SHA256_Module_0.reg9_1x32_0.N_595\, 
        \SHA256_Module_0.reg9_1x32_0.N_589\, 
        SHA256_Module_0_di_req_o, GPIO_0_M2F_c, N_164, N_165, 
        N_119, N_114, N_115, N_116, N_117, N_118, 
        \SHA256_Module_0.reg9_1x32_0.N_594\, 
        \SHA256_Module_0.reg9_1x32_0.N_586\, 
        \SHA256_Module_0.reg9_1x32_0.N_582\, 
        \SHA256_Module_0.reg9_1x32_0.N_578\, 
        \SHA256_Module_0.reg9_1x32_0.N_574\, 
        \SHA256_Module_0.reg9_1x32_0.N_571\, 
        \SHA256_Module_0.reg9_1x32_0.N_570\, 
        \SHA256_Module_0.reg9_1x32_0.N_569\, 
        \SHA256_Module_0.reg9_1x32_0.N_528\, 
        \SHA256_Module_0.reg9_1x32_0.N_523\, 
        \SHA256_Module_0.reg9_1x32_0.N_517\, 
        \SHA256_Module_0.reg9_1x32_0.N_505\, 
        \SHA256_Module_0.reg9_1x32_0.N_503\, 
        \SHA256_Module_0.reg9_1x32_0.N_512\, 
        \SHA256_Module_0.reg9_1x32_0.N_508\, 
        \SHA256_Module_0.reg9_1x32_0.N_504\, 
        \SHA256_Module_0.reg9_1x32_0.N_520\, 
        \SHA256_Module_0.reg9_1x32_0.N_516\, 
        \SHA256_Module_0.SHA256_BLOCK_0.gv_sha256_0.ce_i_i_2_i_0\, 
        \SHA256_Module_0.SHA256_BLOCK_0.sha256_controller_0.N_87_i_0\, 
        \SHA256_Module_0.SHA256_BLOCK_0.sha256_controller_0.N_88_i_0\
         : std_logic;

    for all : SHA256_Module
	Use entity work.SHA256_Module(DEF_ARCH);
    for all : AHB_slave_dummy
	Use entity work.AHB_slave_dummy(DEF_ARCH);
    for all : sha256_system_sb
	Use entity work.sha256_system_sb(DEF_ARCH);
begin 


    SHA256_Module_0 : SHA256_Module
      port map(result_addr_net_0(3) => \result_addr_net_0[3]\, 
        result_addr_net_0(2) => \result_addr_net_0[2]\, 
        result_addr_net_0(1) => \result_addr_net_0[1]\, 
        result_addr_net_0(0) => \result_addr_net_0[0]\, 
        AHB_slave_dummy_0_mem_wdata(31) => 
        \AHB_slave_dummy_0_mem_wdata[31]\, 
        AHB_slave_dummy_0_mem_wdata(30) => 
        \AHB_slave_dummy_0_mem_wdata[30]\, 
        AHB_slave_dummy_0_mem_wdata(29) => 
        \AHB_slave_dummy_0_mem_wdata[29]\, 
        AHB_slave_dummy_0_mem_wdata(28) => 
        \AHB_slave_dummy_0_mem_wdata[28]\, 
        AHB_slave_dummy_0_mem_wdata(27) => 
        \AHB_slave_dummy_0_mem_wdata[27]\, 
        AHB_slave_dummy_0_mem_wdata(26) => 
        \AHB_slave_dummy_0_mem_wdata[26]\, 
        AHB_slave_dummy_0_mem_wdata(25) => 
        \AHB_slave_dummy_0_mem_wdata[25]\, 
        AHB_slave_dummy_0_mem_wdata(24) => 
        \AHB_slave_dummy_0_mem_wdata[24]\, 
        AHB_slave_dummy_0_mem_wdata(23) => 
        \AHB_slave_dummy_0_mem_wdata[23]\, 
        AHB_slave_dummy_0_mem_wdata(22) => 
        \AHB_slave_dummy_0_mem_wdata[22]\, 
        AHB_slave_dummy_0_mem_wdata(21) => 
        \AHB_slave_dummy_0_mem_wdata[21]\, 
        AHB_slave_dummy_0_mem_wdata(20) => 
        \AHB_slave_dummy_0_mem_wdata[20]\, 
        AHB_slave_dummy_0_mem_wdata(19) => 
        \AHB_slave_dummy_0_mem_wdata[19]\, 
        AHB_slave_dummy_0_mem_wdata(18) => 
        \AHB_slave_dummy_0_mem_wdata[18]\, 
        AHB_slave_dummy_0_mem_wdata(17) => 
        \AHB_slave_dummy_0_mem_wdata[17]\, 
        AHB_slave_dummy_0_mem_wdata(16) => 
        \AHB_slave_dummy_0_mem_wdata[16]\, 
        AHB_slave_dummy_0_mem_wdata(15) => 
        \AHB_slave_dummy_0_mem_wdata[15]\, 
        AHB_slave_dummy_0_mem_wdata(14) => 
        \AHB_slave_dummy_0_mem_wdata[14]\, 
        AHB_slave_dummy_0_mem_wdata(13) => 
        \AHB_slave_dummy_0_mem_wdata[13]\, 
        AHB_slave_dummy_0_mem_wdata(12) => 
        \AHB_slave_dummy_0_mem_wdata[12]\, 
        AHB_slave_dummy_0_mem_wdata(11) => 
        \AHB_slave_dummy_0_mem_wdata[11]\, 
        AHB_slave_dummy_0_mem_wdata(10) => 
        \AHB_slave_dummy_0_mem_wdata[10]\, 
        AHB_slave_dummy_0_mem_wdata(9) => 
        \AHB_slave_dummy_0_mem_wdata[9]\, 
        AHB_slave_dummy_0_mem_wdata(8) => 
        \AHB_slave_dummy_0_mem_wdata[8]\, 
        AHB_slave_dummy_0_mem_wdata(7) => 
        \AHB_slave_dummy_0_mem_wdata[7]\, 
        AHB_slave_dummy_0_mem_wdata(6) => 
        \AHB_slave_dummy_0_mem_wdata[6]\, 
        AHB_slave_dummy_0_mem_wdata(5) => 
        \AHB_slave_dummy_0_mem_wdata[5]\, 
        AHB_slave_dummy_0_mem_wdata(4) => 
        \AHB_slave_dummy_0_mem_wdata[4]\, 
        AHB_slave_dummy_0_mem_wdata(3) => 
        \AHB_slave_dummy_0_mem_wdata[3]\, 
        AHB_slave_dummy_0_mem_wdata(2) => 
        \AHB_slave_dummy_0_mem_wdata[2]\, 
        AHB_slave_dummy_0_mem_wdata(1) => 
        \AHB_slave_dummy_0_mem_wdata[1]\, 
        AHB_slave_dummy_0_mem_wdata(0) => 
        \AHB_slave_dummy_0_mem_wdata[0]\, waddr_in_net_0(4) => 
        \waddr_in_net_0[4]\, waddr_in_net_0(3) => 
        \waddr_in_net_0[3]\, waddr_in_net_0(2) => 
        \waddr_in_net_0[2]\, waddr_in_net_0(1) => 
        \waddr_in_net_0[1]\, waddr_in_net_0(0) => 
        \waddr_in_net_0[0]\, state_out_net_0(0) => 
        \state_out_net_0[0]\, line_0_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[7]\, 
        line_3_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[10]\, 
        line_4_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[11]\, 
        line_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[20]\, 
        line_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[28]\, 
        line_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[31]\, 
        line_0_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[7]\, 
        line_0_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[10]\, 
        line_0_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[11]\, 
        line_0_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[20]\, 
        line_0_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[28]\, 
        line_0_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[31]\, 
        line_1_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[7]\, 
        line_1_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[10]\, 
        line_1_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[11]\, 
        line_1_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[20]\, 
        line_1_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[28]\, 
        line_1_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[31]\, 
        line_2_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[7]\, 
        line_2_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[10]\, 
        line_2_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[11]\, 
        line_2_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[20]\, 
        line_2_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[28]\, 
        line_2_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[31]\, 
        line_3_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[7]\, 
        line_3_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[10]\, 
        line_3_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[11]\, 
        line_3_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[20]\, 
        line_3_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[28]\, 
        line_3_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[31]\, 
        line_4_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[7]\, 
        line_4_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[10]\, 
        line_4_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[11]\, 
        line_4_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[20]\, 
        line_4_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[28]\, 
        line_4_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[31]\, 
        line_5_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[7]\, 
        line_5_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[10]\, 
        line_5_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[11]\, 
        line_5_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[20]\, 
        line_5_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[28]\, 
        line_5_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[31]\, 
        line_6_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[7]\, 
        line_6_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[10]\, 
        line_6_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[11]\, 
        line_6_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[20]\, 
        line_6_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[28]\, 
        line_6_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[31]\, 
        line_7_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[28]\, 
        line_7_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[20]\, 
        line_7_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[11]\, 
        line_7_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[10]\, 
        line_7_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[7]\, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, SHA256_Module_0_do_valid_o
         => SHA256_Module_0_do_valid_o, N_568 => 
        \SHA256_Module_0.reg9_1x32_0.N_568\, N_579 => 
        \SHA256_Module_0.reg9_1x32_0.N_579\, N_580 => 
        \SHA256_Module_0.reg9_1x32_0.N_580\, N_581 => 
        \SHA256_Module_0.reg9_1x32_0.N_581\, N_583 => 
        \SHA256_Module_0.reg9_1x32_0.N_583\, N_588 => 
        \SHA256_Module_0.reg9_1x32_0.N_588\, N_589 => 
        \SHA256_Module_0.reg9_1x32_0.N_589\, N_590 => 
        \SHA256_Module_0.reg9_1x32_0.N_590\, N_591 => 
        \SHA256_Module_0.reg9_1x32_0.N_591\, N_592 => 
        \SHA256_Module_0.reg9_1x32_0.N_592\, N_595 => 
        \SHA256_Module_0.reg9_1x32_0.N_595\, N_594 => 
        \SHA256_Module_0.reg9_1x32_0.N_594\, N_586 => 
        \SHA256_Module_0.reg9_1x32_0.N_586\, N_582 => 
        \SHA256_Module_0.reg9_1x32_0.N_582\, N_578 => 
        \SHA256_Module_0.reg9_1x32_0.N_578\, N_574 => 
        \SHA256_Module_0.reg9_1x32_0.N_574\, N_571 => 
        \SHA256_Module_0.reg9_1x32_0.N_571\, N_570 => 
        \SHA256_Module_0.reg9_1x32_0.N_570\, N_569 => 
        \SHA256_Module_0.reg9_1x32_0.N_569\, N_96 => N_96, N_81
         => N_81, N_74 => N_74, N_75 => N_75, N_499 => 
        \SHA256_Module_0.reg9_1x32_0.N_499\, N_501 => 
        \SHA256_Module_0.reg9_1x32_0.N_501\, N_525 => 
        \SHA256_Module_0.reg9_1x32_0.N_525\, N_513 => 
        \SHA256_Module_0.reg9_1x32_0.N_513\, N_502 => 
        \SHA256_Module_0.reg9_1x32_0.N_502\, N_522 => 
        \SHA256_Module_0.reg9_1x32_0.N_522\, N_500 => 
        \SHA256_Module_0.reg9_1x32_0.N_500\, N_514 => 
        \SHA256_Module_0.reg9_1x32_0.N_514\, N_515 => 
        \SHA256_Module_0.reg9_1x32_0.N_515\, N_524 => 
        \SHA256_Module_0.reg9_1x32_0.N_524\, N_526 => 
        \SHA256_Module_0.reg9_1x32_0.N_526\, N_529 => 
        \SHA256_Module_0.reg9_1x32_0.N_529\, N_528 => 
        \SHA256_Module_0.reg9_1x32_0.N_528\, N_523 => 
        \SHA256_Module_0.reg9_1x32_0.N_523\, N_517 => 
        \SHA256_Module_0.reg9_1x32_0.N_517\, N_505 => 
        \SHA256_Module_0.reg9_1x32_0.N_505\, N_503 => 
        \SHA256_Module_0.reg9_1x32_0.N_503\, N_512 => 
        \SHA256_Module_0.reg9_1x32_0.N_512\, N_508 => 
        \SHA256_Module_0.reg9_1x32_0.N_508\, N_504 => 
        \SHA256_Module_0.reg9_1x32_0.N_504\, N_520 => 
        \SHA256_Module_0.reg9_1x32_0.N_520\, N_516 => 
        \SHA256_Module_0.reg9_1x32_0.N_516\, ren_pos => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.ren_pos\, N_228
         => N_228, N_7 => N_7, N_566 => 
        \SHA256_Module_0.reg9_1x32_0.N_566\, N_567 => 
        \SHA256_Module_0.reg9_1x32_0.N_567\, N_565 => 
        \SHA256_Module_0.reg9_1x32_0.N_565\, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready, AHB_slave_dummy_0_read_en
         => AHB_slave_dummy_0_read_en, SHA256_Module_0_error_o
         => SHA256_Module_0_error_o, SHA256_Module_0_di_req_o => 
        SHA256_Module_0_di_req_o, 
        SHA256_Module_0_data_available_lastbank_8 => 
        SHA256_Module_0_data_available_lastbank_8, 
        sha256_system_sb_0_GPIO_9_M2F => 
        sha256_system_sb_0_GPIO_9_M2F, 
        SHA256_Module_0_data_available => 
        SHA256_Module_0_data_available, 
        sha256_system_sb_0_GPIO_1_M2F => 
        sha256_system_sb_0_GPIO_1_M2F, AHB_slave_dummy_0_write_en
         => AHB_slave_dummy_0_write_en, ce_i_i_2_i_0 => 
        \SHA256_Module_0.SHA256_BLOCK_0.gv_sha256_0.ce_i_i_2_i_0\, 
        N_88_i_0 => 
        \SHA256_Module_0.SHA256_BLOCK_0.sha256_controller_0.N_88_i_0\, 
        N_87_i_0 => 
        \SHA256_Module_0.SHA256_BLOCK_0.sha256_controller_0.N_87_i_0\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    AHB_slave_dummy_0 : AHB_slave_dummy
      port map(waddr_in_net_0(4) => \waddr_in_net_0[4]\, 
        waddr_in_net_0(3) => \waddr_in_net_0[3]\, 
        waddr_in_net_0(2) => \waddr_in_net_0[2]\, 
        waddr_in_net_0(1) => \waddr_in_net_0[1]\, 
        waddr_in_net_0(0) => \waddr_in_net_0[0]\, 
        result_addr_net_0(3) => \result_addr_net_0[3]\, 
        result_addr_net_0(2) => \result_addr_net_0[2]\, 
        result_addr_net_0(1) => \result_addr_net_0[1]\, 
        result_addr_net_0(0) => \result_addr_net_0[0]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        arbRegSMCurrentState(15) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.slave_arbiter.arbRegSMCurrentState[15]\, 
        arbRegSMCurrentState(14) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.slave_arbiter.arbRegSMCurrentState[14]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(25) => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[25]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(24) => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[24]\, 
        sha256_system_sb_0_POWER_ON_RESET_N => 
        sha256_system_sb_0_POWER_ON_RESET_N, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, N_118 => N_118, N_117 => 
        N_117, N_116 => N_116, N_115 => N_115, N_114 => N_114, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, 
        AHB_slave_dummy_0_write_en => AHB_slave_dummy_0_write_en, 
        AHB_slave_dummy_0_read_en => AHB_slave_dummy_0_read_en, 
        N_119 => N_119, masterRegAddrSel => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.masterRegAddrSel\, 
        regHTRANS => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.regHTRANS\, 
        N_165 => N_165, N_14_i => N_14_i, N_164 => N_164, 
        defSlaveSMCurrentState => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.default_slave_sm.defSlaveSMCurrentState\, 
        N_31 => N_31);
    
    sha256_system_sb_0 : sha256_system_sb
      port map(
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        arbRegSMCurrentState(15) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.slave_arbiter.arbRegSMCurrentState[15]\, 
        arbRegSMCurrentState(14) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.slave_arbiter.arbRegSMCurrentState[14]\, 
        AHB_slave_dummy_0_mem_wdata(31) => 
        \AHB_slave_dummy_0_mem_wdata[31]\, 
        AHB_slave_dummy_0_mem_wdata(30) => 
        \AHB_slave_dummy_0_mem_wdata[30]\, 
        AHB_slave_dummy_0_mem_wdata(29) => 
        \AHB_slave_dummy_0_mem_wdata[29]\, 
        AHB_slave_dummy_0_mem_wdata(28) => 
        \AHB_slave_dummy_0_mem_wdata[28]\, 
        AHB_slave_dummy_0_mem_wdata(27) => 
        \AHB_slave_dummy_0_mem_wdata[27]\, 
        AHB_slave_dummy_0_mem_wdata(26) => 
        \AHB_slave_dummy_0_mem_wdata[26]\, 
        AHB_slave_dummy_0_mem_wdata(25) => 
        \AHB_slave_dummy_0_mem_wdata[25]\, 
        AHB_slave_dummy_0_mem_wdata(24) => 
        \AHB_slave_dummy_0_mem_wdata[24]\, 
        AHB_slave_dummy_0_mem_wdata(23) => 
        \AHB_slave_dummy_0_mem_wdata[23]\, 
        AHB_slave_dummy_0_mem_wdata(22) => 
        \AHB_slave_dummy_0_mem_wdata[22]\, 
        AHB_slave_dummy_0_mem_wdata(21) => 
        \AHB_slave_dummy_0_mem_wdata[21]\, 
        AHB_slave_dummy_0_mem_wdata(20) => 
        \AHB_slave_dummy_0_mem_wdata[20]\, 
        AHB_slave_dummy_0_mem_wdata(19) => 
        \AHB_slave_dummy_0_mem_wdata[19]\, 
        AHB_slave_dummy_0_mem_wdata(18) => 
        \AHB_slave_dummy_0_mem_wdata[18]\, 
        AHB_slave_dummy_0_mem_wdata(17) => 
        \AHB_slave_dummy_0_mem_wdata[17]\, 
        AHB_slave_dummy_0_mem_wdata(16) => 
        \AHB_slave_dummy_0_mem_wdata[16]\, 
        AHB_slave_dummy_0_mem_wdata(15) => 
        \AHB_slave_dummy_0_mem_wdata[15]\, 
        AHB_slave_dummy_0_mem_wdata(14) => 
        \AHB_slave_dummy_0_mem_wdata[14]\, 
        AHB_slave_dummy_0_mem_wdata(13) => 
        \AHB_slave_dummy_0_mem_wdata[13]\, 
        AHB_slave_dummy_0_mem_wdata(12) => 
        \AHB_slave_dummy_0_mem_wdata[12]\, 
        AHB_slave_dummy_0_mem_wdata(11) => 
        \AHB_slave_dummy_0_mem_wdata[11]\, 
        AHB_slave_dummy_0_mem_wdata(10) => 
        \AHB_slave_dummy_0_mem_wdata[10]\, 
        AHB_slave_dummy_0_mem_wdata(9) => 
        \AHB_slave_dummy_0_mem_wdata[9]\, 
        AHB_slave_dummy_0_mem_wdata(8) => 
        \AHB_slave_dummy_0_mem_wdata[8]\, 
        AHB_slave_dummy_0_mem_wdata(7) => 
        \AHB_slave_dummy_0_mem_wdata[7]\, 
        AHB_slave_dummy_0_mem_wdata(6) => 
        \AHB_slave_dummy_0_mem_wdata[6]\, 
        AHB_slave_dummy_0_mem_wdata(5) => 
        \AHB_slave_dummy_0_mem_wdata[5]\, 
        AHB_slave_dummy_0_mem_wdata(4) => 
        \AHB_slave_dummy_0_mem_wdata[4]\, 
        AHB_slave_dummy_0_mem_wdata(3) => 
        \AHB_slave_dummy_0_mem_wdata[3]\, 
        AHB_slave_dummy_0_mem_wdata(2) => 
        \AHB_slave_dummy_0_mem_wdata[2]\, 
        AHB_slave_dummy_0_mem_wdata(1) => 
        \AHB_slave_dummy_0_mem_wdata[1]\, 
        AHB_slave_dummy_0_mem_wdata(0) => 
        \AHB_slave_dummy_0_mem_wdata[0]\, result_addr_net_0(3)
         => \result_addr_net_0[3]\, result_addr_net_0(2) => 
        \result_addr_net_0[2]\, result_addr_net_0(1) => 
        \result_addr_net_0[1]\, result_addr_net_0(0) => 
        \result_addr_net_0[0]\, state_out_net_0(0) => 
        \state_out_net_0[0]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[25]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[24]\, 
        line_4_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[11]\, 
        line_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[28]\, 
        line_3_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[10]\, 
        line_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[20]\, 
        line_0_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[7]\, line_24
         => \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[31]\, 
        line_0_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[11]\, 
        line_0_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[28]\, 
        line_0_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[10]\, 
        line_0_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[20]\, 
        line_0_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[7]\, 
        line_0_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[31]\, 
        line_1_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[11]\, 
        line_1_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[28]\, 
        line_1_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[10]\, 
        line_1_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[20]\, 
        line_1_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[7]\, 
        line_1_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[31]\, 
        line_2_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[11]\, 
        line_2_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[28]\, 
        line_2_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[10]\, 
        line_2_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[20]\, 
        line_2_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[7]\, 
        line_2_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[31]\, 
        line_3_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[10]\, 
        line_3_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[28]\, 
        line_3_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[7]\, 
        line_3_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[11]\, 
        line_3_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[31]\, 
        line_3_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[20]\, 
        line_4_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[10]\, 
        line_4_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[28]\, 
        line_4_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[7]\, 
        line_4_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[11]\, 
        line_4_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[31]\, 
        line_4_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[20]\, 
        line_5_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[10]\, 
        line_5_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[28]\, 
        line_5_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[7]\, 
        line_5_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[11]\, 
        line_5_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[31]\, 
        line_5_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[20]\, 
        line_6_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[10]\, 
        line_6_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[28]\, 
        line_6_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[7]\, 
        line_6_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[11]\, 
        line_6_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[31]\, 
        line_6_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[20]\, 
        line_7_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[10]\, 
        line_7_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[7]\, 
        line_7_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[20]\, 
        line_7_4 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[11]\, 
        line_7_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[28]\, 
        sha256_system_sb_0_POWER_ON_RESET_N => 
        sha256_system_sb_0_POWER_ON_RESET_N, DEVRST_N => DEVRST_N, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, regHTRANS => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.regHTRANS\, 
        masterRegAddrSel => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.masterRegAddrSel\, 
        N_165 => N_165, N_164 => N_164, N_114 => N_114, N_115 => 
        N_115, N_116 => N_116, N_117 => N_117, N_118 => N_118, 
        N_119 => N_119, N_14_i => N_14_i, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, ren_pos => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.ren_pos\, N_31
         => N_31, defSlaveSMCurrentState => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.default_slave_sm.defSlaveSMCurrentState\, 
        N_96 => N_96, N_516 => 
        \SHA256_Module_0.reg9_1x32_0.N_516\, N_582 => 
        \SHA256_Module_0.reg9_1x32_0.N_582\, N_520 => 
        \SHA256_Module_0.reg9_1x32_0.N_520\, N_586 => 
        \SHA256_Module_0.reg9_1x32_0.N_586\, N_504 => 
        \SHA256_Module_0.reg9_1x32_0.N_504\, N_570 => 
        \SHA256_Module_0.reg9_1x32_0.N_570\, N_508 => 
        \SHA256_Module_0.reg9_1x32_0.N_508\, N_574 => 
        \SHA256_Module_0.reg9_1x32_0.N_574\, N_512 => 
        \SHA256_Module_0.reg9_1x32_0.N_512\, N_578 => 
        \SHA256_Module_0.reg9_1x32_0.N_578\, N_503 => 
        \SHA256_Module_0.reg9_1x32_0.N_503\, N_569 => 
        \SHA256_Module_0.reg9_1x32_0.N_569\, N_505 => 
        \SHA256_Module_0.reg9_1x32_0.N_505\, N_571 => 
        \SHA256_Module_0.reg9_1x32_0.N_571\, N_517 => 
        \SHA256_Module_0.reg9_1x32_0.N_517\, N_583 => 
        \SHA256_Module_0.reg9_1x32_0.N_583\, N_523 => 
        \SHA256_Module_0.reg9_1x32_0.N_523\, N_589 => 
        \SHA256_Module_0.reg9_1x32_0.N_589\, N_528 => 
        \SHA256_Module_0.reg9_1x32_0.N_528\, N_594 => 
        \SHA256_Module_0.reg9_1x32_0.N_594\, N_529 => 
        \SHA256_Module_0.reg9_1x32_0.N_529\, N_595 => 
        \SHA256_Module_0.reg9_1x32_0.N_595\, N_526 => 
        \SHA256_Module_0.reg9_1x32_0.N_526\, N_592 => 
        \SHA256_Module_0.reg9_1x32_0.N_592\, N_524 => 
        \SHA256_Module_0.reg9_1x32_0.N_524\, N_590 => 
        \SHA256_Module_0.reg9_1x32_0.N_590\, N_515 => 
        \SHA256_Module_0.reg9_1x32_0.N_515\, N_581 => 
        \SHA256_Module_0.reg9_1x32_0.N_581\, N_514 => 
        \SHA256_Module_0.reg9_1x32_0.N_514\, N_580 => 
        \SHA256_Module_0.reg9_1x32_0.N_580\, N_522 => 
        \SHA256_Module_0.reg9_1x32_0.N_522\, N_588 => 
        \SHA256_Module_0.reg9_1x32_0.N_588\, N_502 => 
        \SHA256_Module_0.reg9_1x32_0.N_502\, N_568 => 
        \SHA256_Module_0.reg9_1x32_0.N_568\, N_513 => 
        \SHA256_Module_0.reg9_1x32_0.N_513\, N_579 => 
        \SHA256_Module_0.reg9_1x32_0.N_579\, N_525 => 
        \SHA256_Module_0.reg9_1x32_0.N_525\, N_591 => 
        \SHA256_Module_0.reg9_1x32_0.N_591\, N_500 => 
        \SHA256_Module_0.reg9_1x32_0.N_500\, N_566 => 
        \SHA256_Module_0.reg9_1x32_0.N_566\, N_501 => 
        \SHA256_Module_0.reg9_1x32_0.N_501\, N_567 => 
        \SHA256_Module_0.reg9_1x32_0.N_567\, N_499 => 
        \SHA256_Module_0.reg9_1x32_0.N_499\, N_565 => 
        \SHA256_Module_0.reg9_1x32_0.N_565\, N_74 => N_74, N_228
         => N_228, N_81 => N_81, N_7 => N_7, N_75 => N_75, 
        sha256_system_sb_0_GPIO_1_M2F => 
        sha256_system_sb_0_GPIO_1_M2F, GPIO_0_M2F_c => 
        GPIO_0_M2F_c, sha256_system_sb_0_GPIO_9_M2F => 
        sha256_system_sb_0_GPIO_9_M2F, N_87_i_0 => 
        \SHA256_Module_0.SHA256_BLOCK_0.sha256_controller_0.N_87_i_0\, 
        N_88_i_0 => 
        \SHA256_Module_0.SHA256_BLOCK_0.sha256_controller_0.N_88_i_0\, 
        ce_i_i_2_i_0 => 
        \SHA256_Module_0.SHA256_BLOCK_0.gv_sha256_0.ce_i_i_2_i_0\, 
        SHA256_Module_0_data_available_lastbank_8 => 
        SHA256_Module_0_data_available_lastbank_8, 
        SHA256_Module_0_di_req_o => SHA256_Module_0_di_req_o, 
        SHA256_Module_0_data_out_ready => 
        SHA256_Module_0_data_out_ready, 
        SHA256_Module_0_do_valid_o => SHA256_Module_0_do_valid_o, 
        SHA256_Module_0_data_available => 
        SHA256_Module_0_data_available, SHA256_Module_0_error_o
         => SHA256_Module_0_error_o);
    
    GPIO_0_M2F_obuf : OUTBUF
      port map(D => GPIO_0_M2F_c, PAD => GPIO_0_M2F);
    

end DEF_ARCH; 
