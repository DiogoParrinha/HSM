----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Tue Apr 18 22:36:06 2017
-- Parameters for CORESMIP
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant HDL_license : string( 1 to 1 ) := "O";
    constant ZEROIZATION_LEVEL : integer := 3;
end coreparameters;
