-- Version: v11.7 SP1 11.7.1.14

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_8x32 is

    port( raddr_in_net_0                      : in    std_logic_vector(3 downto 0);
          waddr_in_net_0                      : in    std_logic_vector(3 downto 0);
          AHB_slave_dummy_0_mem_wdata         : in    std_logic_vector(31 downto 0);
          data_out_9_0_29                     : out   std_logic;
          data_out_9_0_1                      : out   std_logic;
          data_out_9_0_0                      : out   std_logic;
          data_out_9_0_31                     : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK        : in    std_logic;
          sha256_system_sb_0_POWER_ON_RESET_N : in    std_logic;
          N_1323                              : out   std_logic;
          N_1328                              : out   std_logic;
          N_1330                              : out   std_logic;
          N_1331                              : out   std_logic;
          N_1332                              : out   std_logic;
          N_1324                              : out   std_logic;
          N_1325                              : out   std_logic;
          N_1326                              : out   std_logic;
          N_1329                              : out   std_logic;
          N_1333                              : out   std_logic;
          N_1334                              : out   std_logic;
          N_1335                              : out   std_logic;
          N_1336                              : out   std_logic;
          N_1337                              : out   std_logic;
          N_1338                              : out   std_logic;
          N_1339                              : out   std_logic;
          N_1340                              : out   std_logic;
          N_1341                              : out   std_logic;
          N_1342                              : out   std_logic;
          N_1343                              : out   std_logic;
          N_1344                              : out   std_logic;
          N_1345                              : out   std_logic;
          N_1327                              : out   std_logic;
          N_1346                              : out   std_logic;
          N_1347                              : out   std_logic;
          N_1348                              : out   std_logic;
          N_1349                              : out   std_logic;
          N_1351                              : out   std_logic;
          N_1270                              : out   std_logic;
          N_1256                              : out   std_logic;
          N_1261                              : out   std_logic;
          N_1263                              : out   std_logic;
          N_1265                              : out   std_logic;
          N_1257                              : out   std_logic;
          N_1258                              : out   std_logic;
          N_1259                              : out   std_logic;
          N_1262                              : out   std_logic;
          N_1264                              : out   std_logic;
          N_1266                              : out   std_logic;
          N_1267                              : out   std_logic;
          N_1268                              : out   std_logic;
          N_1269                              : out   std_logic;
          N_1271                              : out   std_logic;
          N_1272                              : out   std_logic;
          N_1273                              : out   std_logic;
          N_1274                              : out   std_logic;
          N_1275                              : out   std_logic;
          N_1276                              : out   std_logic;
          N_1277                              : out   std_logic;
          N_1278                              : out   std_logic;
          N_1260                              : out   std_logic;
          N_1279                              : out   std_logic;
          N_1280                              : out   std_logic;
          N_1281                              : out   std_logic;
          N_1282                              : out   std_logic;
          N_1284                              : out   std_logic;
          AHB_slave_dummy_0_read_en           : in    std_logic;
          AHB_slave_dummy_0_write_en          : in    std_logic;
          N_1446                              : out   std_logic;
          N_53                                : out   std_logic;
          N_1458                              : out   std_logic;
          N_1457                              : out   std_logic;
          data_out_sn_N_12_mux                : out   std_logic;
          N_1423_3                            : out   std_logic
        );

end reg_8x32;

architecture DEF_ARCH of reg_8x32 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \ren_pos\, VCC_net_1, N_35_i_0, GND_net_1, 
        \line3[63]_net_1\, N_18_i_0, \line3_or[0]_net_1\, 
        \line3[62]_net_1\, \line3_5[62]_net_1\, \line3[61]_net_1\, 
        N_1439_i_0, \line3[60]_net_1\, \line3_5[60]_net_1\, 
        \line3[59]_net_1\, \line3_5[59]_net_1\, \line3[58]_net_1\, 
        \line3_5[58]_net_1\, \line3[57]_net_1\, 
        \line3_5[57]_net_1\, \line3[56]_net_1\, 
        \line3_5[56]_net_1\, \line3[55]_net_1\, 
        \line3_5[55]_net_1\, \line3[54]_net_1\, 
        \line3_5[54]_net_1\, \line3[53]_net_1\, 
        \line3_5[53]_net_1\, \line3[52]_net_1\, 
        \line3_5[52]_net_1\, \line3[51]_net_1\, 
        \line3_5[51]_net_1\, \line3[50]_net_1\, 
        \line3_5[50]_net_1\, \line3[49]_net_1\, 
        \line3_5[49]_net_1\, \line3[48]_net_1\, 
        \line3_5[48]_net_1\, \line3[47]_net_1\, 
        \line3_5[47]_net_1\, \line3[46]_net_1\, 
        \line3_5[46]_net_1\, \line3[45]_net_1\, 
        \line3_5[45]_net_1\, \line3[44]_net_1\, 
        \line3_5[44]_net_1\, \line3[43]_net_1\, 
        \line3_5[43]_net_1\, \line3[42]_net_1\, 
        \line3_5[42]_net_1\, \line3[41]_net_1\, 
        \line3_5[41]_net_1\, \line3[40]_net_1\, 
        \line3_5[40]_net_1\, \line3[39]_net_1\, 
        \line3_5[39]_net_1\, \line3[38]_net_1\, 
        \line3_5[38]_net_1\, \line3[37]_net_1\, 
        \line3_5[37]_net_1\, \line3[36]_net_1\, 
        \line3_5[36]_net_1\, \line3[35]_net_1\, 
        \line3_5[35]_net_1\, \line3[34]_net_1\, 
        \line3_5[34]_net_1\, \line3[33]_net_1\, 
        \line3_5[33]_net_1\, \line3[32]_net_1\, 
        \line3_5[32]_net_1\, \line3[31]_net_1\, N_20_i_0, 
        \line3[30]_net_1\, \line3_5[30]_net_1\, \line3[29]_net_1\, 
        N_1440_i_0, \line3[28]_net_1\, \line3_5[28]_net_1\, 
        \line3[27]_net_1\, \line3_5[27]_net_1\, \line3[26]_net_1\, 
        \line3_5[26]_net_1\, \line3[25]_net_1\, 
        \line3_5[25]_net_1\, \line3[24]_net_1\, 
        \line3_5[24]_net_1\, \line3[23]_net_1\, 
        \line3_5[23]_net_1\, \line3[22]_net_1\, 
        \line3_5[22]_net_1\, \line3[21]_net_1\, 
        \line3_5[21]_net_1\, \line3[20]_net_1\, 
        \line3_5[20]_net_1\, \line3[19]_net_1\, 
        \line3_5[19]_net_1\, \line3[18]_net_1\, 
        \line3_5[18]_net_1\, \line3[17]_net_1\, 
        \line3_5[17]_net_1\, \line3[16]_net_1\, 
        \line3_5[16]_net_1\, \line3[15]_net_1\, 
        \line3_5[15]_net_1\, \line3[14]_net_1\, 
        \line3_5[14]_net_1\, \line3[13]_net_1\, 
        \line3_5[13]_net_1\, \line3[12]_net_1\, 
        \line3_5[12]_net_1\, \line3[11]_net_1\, 
        \line3_5[11]_net_1\, \line3[10]_net_1\, 
        \line3_5[10]_net_1\, \line3[9]_net_1\, \line3_5[9]_net_1\, 
        \line3[8]_net_1\, \line3_5[8]_net_1\, \line3[7]_net_1\, 
        \line3_5[7]_net_1\, \line3[6]_net_1\, \line3_5[6]_net_1\, 
        \line3[5]_net_1\, \line3_5[5]_net_1\, \line3[4]_net_1\, 
        \line3_5[4]_net_1\, \line3[3]_net_1\, \line3_5[3]_net_1\, 
        \line3[2]_net_1\, \line3_5[2]_net_1\, \line3[1]_net_1\, 
        \line3_5[1]_net_1\, \line3[0]_net_1\, \line3_5[0]_net_1\, 
        un1_wen_18_or, \line2[63]_net_1\, N_22_i_0, un1_wen_19_or, 
        \line2[62]_net_1\, \line2_5[62]_net_1\, \line2[61]_net_1\, 
        N_1441_i_0, \line2[60]_net_1\, \line2_5[60]_net_1\, 
        \line2[59]_net_1\, \line2_5[59]_net_1\, \line2[58]_net_1\, 
        \line2_5[58]_net_1\, \line2[57]_net_1\, 
        \line2_5[57]_net_1\, \line2[56]_net_1\, 
        \line2_5[56]_net_1\, \line2[55]_net_1\, 
        \line2_5[55]_net_1\, \line2[54]_net_1\, 
        \line2_5[54]_net_1\, \line2[53]_net_1\, 
        \line2_5[53]_net_1\, \line2[52]_net_1\, 
        \line2_5[52]_net_1\, \line2[51]_net_1\, 
        \line2_5[51]_net_1\, \line2[50]_net_1\, 
        \line2_5[50]_net_1\, \line2[49]_net_1\, 
        \line2_5[49]_net_1\, \line2[48]_net_1\, 
        \line2_5[48]_net_1\, \line2[47]_net_1\, 
        \line2_5[47]_net_1\, \line2[46]_net_1\, 
        \line2_5[46]_net_1\, \line2[45]_net_1\, 
        \line2_5[45]_net_1\, \line2[44]_net_1\, 
        \line2_5[44]_net_1\, \line2[43]_net_1\, 
        \line2_5[43]_net_1\, \line2[42]_net_1\, 
        \line2_5[42]_net_1\, \line2[41]_net_1\, 
        \line2_5[41]_net_1\, \line2[40]_net_1\, 
        \line2_5[40]_net_1\, \line2[39]_net_1\, 
        \line2_5[39]_net_1\, \line2[38]_net_1\, 
        \line2_5[38]_net_1\, \line2[37]_net_1\, 
        \line2_5[37]_net_1\, \line2[36]_net_1\, 
        \line2_5[36]_net_1\, \line2[35]_net_1\, 
        \line2_5[35]_net_1\, \line2[34]_net_1\, 
        \line2_5[34]_net_1\, \line2[33]_net_1\, 
        \line2_5[33]_net_1\, \line2[32]_net_1\, 
        \line2_5[32]_net_1\, \line2[31]_net_1\, N_24_i_0, 
        \line2[30]_net_1\, \line2_5[30]_net_1\, \line2[29]_net_1\, 
        N_1442_i_0, \line2[28]_net_1\, \line2_5[28]_net_1\, 
        \line2[27]_net_1\, \line2_5[27]_net_1\, \line2[26]_net_1\, 
        \line2_5[26]_net_1\, \line2[25]_net_1\, 
        \line2_5[25]_net_1\, \line2[24]_net_1\, 
        \line2_5[24]_net_1\, \line2[23]_net_1\, 
        \line2_5[23]_net_1\, \line2[22]_net_1\, 
        \line2_5[22]_net_1\, \line2[21]_net_1\, 
        \line2_5[21]_net_1\, \line2[20]_net_1\, 
        \line2_5[20]_net_1\, \line2[19]_net_1\, 
        \line2_5[19]_net_1\, \line2[18]_net_1\, 
        \line2_5[18]_net_1\, \line2[17]_net_1\, 
        \line2_5[17]_net_1\, \line2[16]_net_1\, 
        \line2_5[16]_net_1\, \line2[15]_net_1\, 
        \line2_5[15]_net_1\, \line2[14]_net_1\, 
        \line2_5[14]_net_1\, \line2[13]_net_1\, 
        \line2_5[13]_net_1\, \line2[12]_net_1\, 
        \line2_5[12]_net_1\, \line2[11]_net_1\, 
        \line2_5[11]_net_1\, \line2[10]_net_1\, 
        \line2_5[10]_net_1\, \line2[9]_net_1\, \line2_5[9]_net_1\, 
        \line2[8]_net_1\, \line2_5[8]_net_1\, \line2[7]_net_1\, 
        \line2_5[7]_net_1\, \line2[6]_net_1\, \line2_5[6]_net_1\, 
        \line2[5]_net_1\, \line2_5[5]_net_1\, \line2[4]_net_1\, 
        \line2_5[4]_net_1\, \line2[3]_net_1\, \line2_5[3]_net_1\, 
        \line2[2]_net_1\, \line2_5[2]_net_1\, \line2[1]_net_1\, 
        \line2_5[1]_net_1\, \line2[0]_net_1\, \line2_5[0]_net_1\, 
        \line1[63]_net_1\, N_26_i_0, un1_wen_20_or, 
        \line1[62]_net_1\, \line1_5[62]_net_1\, \line1[61]_net_1\, 
        N_1443_i_0, \line1[60]_net_1\, \line1_5[60]_net_1\, 
        \line1[59]_net_1\, \line1_5[59]_net_1\, \line1[58]_net_1\, 
        \line1_5[58]_net_1\, \line1[57]_net_1\, 
        \line1_5[57]_net_1\, \line1[56]_net_1\, 
        \line1_5[56]_net_1\, \line1[55]_net_1\, 
        \line1_5[55]_net_1\, \line1[54]_net_1\, 
        \line1_5[54]_net_1\, \line1[53]_net_1\, 
        \line1_5[53]_net_1\, \line1[52]_net_1\, 
        \line1_5[52]_net_1\, \line1[51]_net_1\, 
        \line1_5[51]_net_1\, \line1[50]_net_1\, 
        \line1_5[50]_net_1\, \line1[49]_net_1\, 
        \line1_5[49]_net_1\, \line1[48]_net_1\, 
        \line1_5[48]_net_1\, \line1[47]_net_1\, 
        \line1_5[47]_net_1\, \line1[46]_net_1\, 
        \line1_5[46]_net_1\, \line1[45]_net_1\, 
        \line1_5[45]_net_1\, \line1[44]_net_1\, 
        \line1_5[44]_net_1\, \line1[43]_net_1\, 
        \line1_5[43]_net_1\, \line1[42]_net_1\, 
        \line1_5[42]_net_1\, \line1[41]_net_1\, 
        \line1_5[41]_net_1\, \line1[40]_net_1\, 
        \line1_5[40]_net_1\, \line1[39]_net_1\, 
        \line1_5[39]_net_1\, \line1[38]_net_1\, 
        \line1_5[38]_net_1\, \line1[37]_net_1\, 
        \line1_5[37]_net_1\, \line1[36]_net_1\, 
        \line1_5[36]_net_1\, \line1[35]_net_1\, 
        \line1_5[35]_net_1\, \line1[34]_net_1\, 
        \line1_5[34]_net_1\, \line1[33]_net_1\, 
        \line1_5[33]_net_1\, \line1[32]_net_1\, 
        \line1_5[32]_net_1\, \line1[31]_net_1\, N_28_i_0, 
        \line1[30]_net_1\, \line1_5[30]_net_1\, \line1[29]_net_1\, 
        N_34_i_0, \line1[28]_net_1\, \line1_5[28]_net_1\, 
        \line1[27]_net_1\, \line1_5[27]_net_1\, \line1[26]_net_1\, 
        \line1_5[26]_net_1\, \line1[25]_net_1\, 
        \line1_5[25]_net_1\, \line1[24]_net_1\, 
        \line1_5[24]_net_1\, \line1[23]_net_1\, 
        \line1_5[23]_net_1\, \line1[22]_net_1\, 
        \line1_5[22]_net_1\, \line1[21]_net_1\, 
        \line1_5[21]_net_1\, \line1[20]_net_1\, 
        \line1_5[20]_net_1\, \line1[19]_net_1\, 
        \line1_5[19]_net_1\, \line1[18]_net_1\, 
        \line1_5[18]_net_1\, \line1[17]_net_1\, 
        \line1_5[17]_net_1\, \line1[16]_net_1\, 
        \line1_5[16]_net_1\, \line1[15]_net_1\, 
        \line1_5[15]_net_1\, \line1[14]_net_1\, 
        \line1_5[14]_net_1\, \line1[13]_net_1\, 
        \line1_5[13]_net_1\, \line1[12]_net_1\, 
        \line1_5[12]_net_1\, \line1[11]_net_1\, 
        \line1_5[11]_net_1\, \line1[10]_net_1\, 
        \line1_5[10]_net_1\, \line1[9]_net_1\, \line1_5[9]_net_1\, 
        \line1[8]_net_1\, \line1_5[8]_net_1\, \line1[7]_net_1\, 
        \line1_5[7]_net_1\, \line1[6]_net_1\, \line1_5[6]_net_1\, 
        \line1[5]_net_1\, \line1_5[5]_net_1\, \line1[4]_net_1\, 
        \line1_5[4]_net_1\, \line1[3]_net_1\, \line1_5[3]_net_1\, 
        \line1[2]_net_1\, \line1_5[2]_net_1\, \line1[1]_net_1\, 
        \line1_5[1]_net_1\, \line1[0]_net_1\, \line1_5[0]_net_1\, 
        \line4[63]_net_1\, \line4_5[63]\, un1_wen_4_or, 
        \line4[62]_net_1\, \line4_5[62]_net_1\, \line4[61]_net_1\, 
        N_1437_i_0, \line4[60]_net_1\, \line4_5[60]_net_1\, 
        \line4[59]_net_1\, \line4_5[59]_net_1\, \line4[58]_net_1\, 
        \line4_5[58]_net_1\, \line4[57]_net_1\, 
        \line4_5[57]_net_1\, \line4[56]_net_1\, 
        \line4_5[56]_net_1\, \line4[55]_net_1\, 
        \line4_5[55]_net_1\, \line4[54]_net_1\, 
        \line4_5[54]_net_1\, \line4[53]_net_1\, 
        \line4_5[53]_net_1\, \line4[52]_net_1\, 
        \line4_5[52]_net_1\, \line4[51]_net_1\, 
        \line4_5[51]_net_1\, \line4[50]_net_1\, 
        \line4_5[50]_net_1\, \line4[49]_net_1\, 
        \line4_5[49]_net_1\, \line4[48]_net_1\, 
        \line4_5[48]_net_1\, \line4[47]_net_1\, 
        \line4_5[47]_net_1\, \line4[46]_net_1\, 
        \line4_5[46]_net_1\, \line4[45]_net_1\, 
        \line4_5[45]_net_1\, \line4[44]_net_1\, 
        \line4_5[44]_net_1\, \line4[43]_net_1\, 
        \line4_5[43]_net_1\, \line4[42]_net_1\, 
        \line4_5[42]_net_1\, \line4[41]_net_1\, 
        \line4_5[41]_net_1\, \line4[40]_net_1\, 
        \line4_5[40]_net_1\, \line4[39]_net_1\, 
        \line4_5[39]_net_1\, \line4[38]_net_1\, 
        \line4_5[38]_net_1\, \line4[37]_net_1\, 
        \line4_5[37]_net_1\, \line4[36]_net_1\, 
        \line4_5[36]_net_1\, \line4[35]_net_1\, 
        \line4_5[35]_net_1\, \line4[34]_net_1\, 
        \line4_5[34]_net_1\, \line4[33]_net_1\, 
        \line4_5[33]_net_1\, \line4[32]_net_1\, \line4_5[32]\, 
        \line4[31]_net_1\, \line4_5[31]\, \line4[30]_net_1\, 
        \line4_5[30]_net_1\, \line4[29]_net_1\, N_1438_i_0, 
        \line4[28]_net_1\, \line4_5[28]_net_1\, \line4[27]_net_1\, 
        \line4_5[27]_net_1\, \line4[26]_net_1\, 
        \line4_5[26]_net_1\, \line4[25]_net_1\, 
        \line4_5[25]_net_1\, \line4[24]_net_1\, 
        \line4_5[24]_net_1\, \line4[23]_net_1\, 
        \line4_5[23]_net_1\, \line4[22]_net_1\, 
        \line4_5[22]_net_1\, \line4[21]_net_1\, 
        \line4_5[21]_net_1\, \line4[20]_net_1\, 
        \line4_5[20]_net_1\, \line4[19]_net_1\, 
        \line4_5[19]_net_1\, \line4[18]_net_1\, 
        \line4_5[18]_net_1\, \line4[17]_net_1\, 
        \line4_5[17]_net_1\, \line4[16]_net_1\, 
        \line4_5[16]_net_1\, \line4[15]_net_1\, 
        \line4_5[15]_net_1\, \line4[14]_net_1\, 
        \line4_5[14]_net_1\, \line4[13]_net_1\, 
        \line4_5[13]_net_1\, \line4[12]_net_1\, 
        \line4_5[12]_net_1\, \line4[11]_net_1\, 
        \line4_5[11]_net_1\, \line4[10]_net_1\, 
        \line4_5[10]_net_1\, \line4[9]_net_1\, \line4_5[9]_net_1\, 
        \line4[8]_net_1\, \line4_5[8]_net_1\, \line4[7]_net_1\, 
        \line4_5[7]_net_1\, \line4[6]_net_1\, \line4_5[6]_net_1\, 
        \line4[5]_net_1\, \line4_5[5]_net_1\, \line4[4]_net_1\, 
        \line4_5[4]_net_1\, \line4[3]_net_1\, \line4_5[3]_net_1\, 
        \line4[2]_net_1\, \line4_5[2]_net_1\, \line4[1]_net_1\, 
        \line4_5[1]_net_1\, \line4[0]_net_1\, \line4_5[0]_net_1\, 
        \line0[63]_net_1\, N_30_i_0, un1_wen_7_or, 
        \line0[62]_net_1\, \line0_6[62]_net_1\, \line0[61]_net_1\, 
        N_36_i_0, \line0[60]_net_1\, \line0_6[60]_net_1\, 
        \line0[59]_net_1\, \line0_6[59]_net_1\, \line0[58]_net_1\, 
        \line0_6[58]_net_1\, \line0[57]_net_1\, 
        \line0_6[57]_net_1\, \line0[56]_net_1\, 
        \line0_6[56]_net_1\, \line0[55]_net_1\, 
        \line0_6[55]_net_1\, \line0[54]_net_1\, 
        \line0_6[54]_net_1\, \line0[53]_net_1\, 
        \line0_6[53]_net_1\, \line0[52]_net_1\, 
        \line0_6[52]_net_1\, \line0[51]_net_1\, 
        \line0_6[51]_net_1\, \line0[50]_net_1\, 
        \line0_6[50]_net_1\, \line0[49]_net_1\, 
        \line0_6[49]_net_1\, \line0[48]_net_1\, 
        \line0_6[48]_net_1\, \line0[47]_net_1\, 
        \line0_6[47]_net_1\, \line0[46]_net_1\, 
        \line0_6[46]_net_1\, \line0[45]_net_1\, 
        \line0_6[45]_net_1\, \line0[44]_net_1\, 
        \line0_6[44]_net_1\, \line0[43]_net_1\, 
        \line0_6[43]_net_1\, \line0[42]_net_1\, 
        \line0_6[42]_net_1\, \line0[41]_net_1\, 
        \line0_6[41]_net_1\, \line0[40]_net_1\, 
        \line0_6[40]_net_1\, \line0[39]_net_1\, 
        \line0_6[39]_net_1\, \line0[38]_net_1\, 
        \line0_6[38]_net_1\, \line0[37]_net_1\, 
        \line0_6[37]_net_1\, \line0[36]_net_1\, 
        \line0_6[36]_net_1\, \line0[35]_net_1\, 
        \line0_6[35]_net_1\, \line0[34]_net_1\, 
        \line0_6[34]_net_1\, \line0[33]_net_1\, 
        \line0_6[33]_net_1\, \line0[32]_net_1\, 
        \line0_6[32]_net_1\, \line0[31]_net_1\, N_32_i_0, 
        \line0[30]_net_1\, \line0_6[30]_net_1\, \line0[29]_net_1\, 
        N_38_i_0, \line0[28]_net_1\, \line0_6[28]_net_1\, 
        \line0[27]_net_1\, \line0_6[27]_net_1\, \line0[26]_net_1\, 
        \line0_6[26]_net_1\, \line0[25]_net_1\, 
        \line0_6[25]_net_1\, \line0[24]_net_1\, 
        \line0_6[24]_net_1\, \line0[23]_net_1\, 
        \line0_6[23]_net_1\, \line0[22]_net_1\, 
        \line0_6[22]_net_1\, \line0[21]_net_1\, 
        \line0_6[21]_net_1\, \line0[20]_net_1\, 
        \line0_6[20]_net_1\, \line0[19]_net_1\, 
        \line0_6[19]_net_1\, \line0[18]_net_1\, 
        \line0_6[18]_net_1\, \line0[17]_net_1\, 
        \line0_6[17]_net_1\, \line0[16]_net_1\, 
        \line0_6[16]_net_1\, \line0[15]_net_1\, 
        \line0_6[15]_net_1\, \line0[14]_net_1\, 
        \line0_6[14]_net_1\, \line0[13]_net_1\, 
        \line0_6[13]_net_1\, \line0[12]_net_1\, 
        \line0_6[12]_net_1\, \line0[11]_net_1\, 
        \line0_6[11]_net_1\, \line0[10]_net_1\, 
        \line0_6[10]_net_1\, \line0[9]_net_1\, \line0_6[9]_net_1\, 
        \line0[8]_net_1\, \line0_6[8]_net_1\, \line0[7]_net_1\, 
        \line0_6[7]_net_1\, \line0[6]_net_1\, \line0_6[6]_net_1\, 
        \line0[5]_net_1\, \line0_6[5]_net_1\, \line0[4]_net_1\, 
        \line0_6[4]_net_1\, \line0[3]_net_1\, \line0_6[3]_net_1\, 
        \line0[2]_net_1\, \line0_6[2]_net_1\, \line0[1]_net_1\, 
        \line0_6[1]_net_1\, \line0[0]_net_1\, \line0_6[0]_net_1\, 
        \raddr_pos[3]_net_1\, N_1424_i_0, \raddr_pos[2]_net_1\, 
        \raddr_pos[1]_net_1\, \raddr_pos[0]_net_1\, 
        \raddr_pos_fast[3]_net_1\, \raddr_pos_3_rep1\, 
        \raddr_pos_3_rep2\, N_47_i, \data_out_8_bm_1_1[2]_net_1\, 
        \data_out_8_bm[2]_net_1\, \data_out_8_bm_1_1[7]_net_1\, 
        \data_out_8_bm[7]_net_1\, \data_out_8_bm_1_1[9]_net_1\, 
        \data_out_8_bm[9]_net_1\, \data_out_8_bm_1_1[10]_net_1\, 
        \data_out_8_bm[10]_net_1\, \data_out_8_bm_1_1[11]_net_1\, 
        \data_out_8_bm[11]_net_1\, \data_out_8_bm_1_1[3]_net_1\, 
        \data_out_8_bm[3]_net_1\, \data_out_8_bm_1_1[4]_net_1\, 
        \data_out_8_bm[4]_net_1\, \data_out_8_bm_1_1[5]_net_1\, 
        \data_out_8_bm[5]_net_1\, \data_out_8_bm_1_1[8]_net_1\, 
        \data_out_8_bm[8]_net_1\, \data_out_8_bm_1_1[12]_net_1\, 
        \data_out_8_bm[12]_net_1\, \data_out_8_bm_1_1[13]_net_1\, 
        \data_out_8_bm[13]_net_1\, \data_out_8_bm_1_1[14]_net_1\, 
        \data_out_8_bm[14]_net_1\, \data_out_8_bm_1_1[15]_net_1\, 
        \data_out_8_bm[15]_net_1\, \data_out_8_bm_1_1[16]_net_1\, 
        \data_out_8_bm[16]_net_1\, \data_out_8_bm_1_1[17]_net_1\, 
        \data_out_8_bm[17]_net_1\, \data_out_8_bm_1_1[18]_net_1\, 
        \data_out_8_bm[18]_net_1\, \data_out_8_bm_1_1[19]_net_1\, 
        \data_out_8_bm[19]_net_1\, \data_out_8_bm_1_1[20]_net_1\, 
        \data_out_8_bm[20]_net_1\, \data_out_8_bm_1_1[21]_net_1\, 
        \data_out_8_bm[21]_net_1\, \data_out_8_bm_1_1[22]_net_1\, 
        \data_out_8_bm[22]_net_1\, \data_out_8_bm_1_1[23]_net_1\, 
        \data_out_8_bm[23]_net_1\, \data_out_8_bm_1_1[24]_net_1\, 
        \data_out_8_bm[24]_net_1\, \data_out_8_bm_1_1[6]_net_1\, 
        \data_out_8_bm[6]_net_1\, \data_out_8_bm_1_1[25]_net_1\, 
        \data_out_8_bm[25]_net_1\, \data_out_8_bm_1_1[26]_net_1\, 
        \data_out_8_bm[26]_net_1\, \data_out_8_bm_1_1[27]_net_1\, 
        \data_out_8_bm[27]_net_1\, \data_out_8_bm_1_1[28]_net_1\, 
        \data_out_8_bm[28]_net_1\, \data_out_8_bm_1_1[30]_net_1\, 
        \data_out_8_bm[30]_net_1\, \data_out_9_m2_0_1_1[31]\, 
        N_56, \data_out_5_i_m2_1_1[0]\, N_1456, 
        \data_out_9_m2_1_1_1[29]\, N_1468, 
        \data_out_5_i_m2_1_1[1]\, N_1455, data_out_sn_N_11_mux, 
        \data_out_8_am[2]_net_1\, \data_out_8_am[7]_net_1\, 
        \data_out_8_am[9]_net_1\, \data_out_8_am[10]_net_1\, 
        \data_out_8_am[11]_net_1\, \data_out_8_am[3]_net_1\, 
        \data_out_8_am[4]_net_1\, \data_out_8_am[5]_net_1\, 
        \data_out_8_am[8]_net_1\, \data_out_8_am[12]_net_1\, 
        \data_out_8_am[13]_net_1\, \data_out_8_am[14]_net_1\, 
        \data_out_8_am[15]_net_1\, \data_out_8_am[16]_net_1\, 
        \data_out_8_am[17]_net_1\, \data_out_8_am[18]_net_1\, 
        \data_out_8_am[19]_net_1\, \data_out_8_am[20]_net_1\, 
        \data_out_8_am[21]_net_1\, \data_out_8_am[22]_net_1\, 
        \data_out_8_am[23]_net_1\, \data_out_8_am[24]_net_1\, 
        \data_out_8_am[6]_net_1\, \data_out_8_am[25]_net_1\, 
        \data_out_8_am[26]_net_1\, \data_out_8_am[27]_net_1\, 
        \data_out_8_am[28]_net_1\, \data_out_8_am[30]_net_1\, 
        \data_out_6_i_m2_bm[1]_net_1\, 
        \data_out_6_i_m2_am[1]_net_1\, N_1453, 
        \data_out_6_i_m2_bm[0]_net_1\, 
        \data_out_6_i_m2_am[0]_net_1\, N_1454, 
        \data_out_9_m2_1_bm[31]_net_1\, 
        \data_out_9_m2_1_am[31]_net_1\, N_60, 
        \data_out_6_bm[16]_net_1\, \data_out_6_am[16]_net_1\, 
        \data_out_6_bm[2]_net_1\, \data_out_6_am[2]_net_1\, 
        \data_out_6_bm[7]_net_1\, \data_out_6_am[7]_net_1\, 
        \data_out_6_bm[9]_net_1\, \data_out_6_am[9]_net_1\, 
        \data_out_6_bm[11]_net_1\, \data_out_6_am[11]_net_1\, 
        \data_out_6_bm[3]_net_1\, \data_out_6_am[3]_net_1\, 
        \data_out_6_bm[4]_net_1\, \data_out_6_am[4]_net_1\, 
        \data_out_6_bm[5]_net_1\, \data_out_6_am[5]_net_1\, 
        \data_out_6_bm[8]_net_1\, \data_out_6_am[8]_net_1\, 
        \data_out_6_bm[10]_net_1\, \data_out_6_am[10]_net_1\, 
        \data_out_6_bm[12]_net_1\, \data_out_6_am[12]_net_1\, 
        \data_out_6_bm[13]_net_1\, \data_out_6_am[13]_net_1\, 
        \data_out_6_bm[14]_net_1\, \data_out_6_am[14]_net_1\, 
        \data_out_6_bm[15]_net_1\, \data_out_6_am[15]_net_1\, 
        \data_out_6_bm[17]_net_1\, \data_out_6_am[17]_net_1\, 
        \data_out_6_bm[18]_net_1\, \data_out_6_am[18]_net_1\, 
        \data_out_6_bm[19]_net_1\, \data_out_6_am[19]_net_1\, 
        \data_out_6_bm[20]_net_1\, \data_out_6_am[20]_net_1\, 
        \data_out_6_bm[21]_net_1\, \data_out_6_am[21]_net_1\, 
        \data_out_6_bm[22]_net_1\, \data_out_6_am[22]_net_1\, 
        \data_out_6_bm[23]_net_1\, \data_out_6_am[23]_net_1\, 
        \data_out_6_bm[24]_net_1\, \data_out_6_am[24]_net_1\, 
        \data_out_6_bm[6]_net_1\, \data_out_6_am[6]_net_1\, 
        \data_out_6_bm[25]_net_1\, \data_out_6_am[25]_net_1\, 
        \data_out_6_bm[26]_net_1\, \data_out_6_am[26]_net_1\, 
        \data_out_6_bm[27]_net_1\, \data_out_6_am[27]_net_1\, 
        \data_out_6_bm[28]_net_1\, \data_out_6_am[28]_net_1\, 
        \data_out_9_m2_0_bm[29]_net_1\, 
        \data_out_9_m2_0_am[29]_net_1\, N_1467, 
        \data_out_6_bm[30]_net_1\, \data_out_6_am[30]_net_1\, 
        N_1423_1, N_44, N_1434, N_61, N_62, 
        \data_out_sn_N_12_mux\, \un1_wen_18_or_0_0\, un5_wen, 
        N_46 : std_logic;

begin 

    data_out_sn_N_12_mux <= \data_out_sn_N_12_mux\;

    \line3[15]\ : SLE
      port map(D => \line3_5[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[15]_net_1\);
    
    \line2_5[51]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(19), C => \line2[51]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[51]_net_1\);
    
    \line3[41]\ : SLE
      port map(D => \line3_5[41]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[41]_net_1\);
    
    \line0_6[54]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(22), C => \line0[54]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[54]_net_1\);
    
    \line1[30]\ : SLE
      port map(D => \line1_5[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[30]_net_1\);
    
    \line1[16]\ : SLE
      port map(D => \line1_5[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[16]_net_1\);
    
    \line2_RNO[31]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(31), C => \line2[31]_net_1\, 
        D => waddr_in_net_0(0), Y => N_24_i_0);
    
    \data_out_8_am[19]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[51]_net_1\, D => \line1[19]_net_1\, Y => 
        \data_out_8_am[19]_net_1\);
    
    \line1[22]\ : SLE
      port map(D => \line1_5[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[22]_net_1\);
    
    \line3[0]\ : SLE
      port map(D => \line3_5[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[0]_net_1\);
    
    \line1[14]\ : SLE
      port map(D => \line1_5[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[14]_net_1\);
    
    \line0_6[25]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(25), C => \line0[25]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[25]_net_1\);
    
    \line3_5[7]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(7), C => \line3[7]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[7]_net_1\);
    
    \line4_5[57]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(25), 
        C => \line4[57]_net_1\, D => N_47_i, Y => 
        \line4_5[57]_net_1\);
    
    \line3_5[24]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(24), C => \line3[24]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[24]_net_1\);
    
    \data_out_8_ns[27]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[27]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[27]_net_1\, Y
         => N_1348);
    
    \data_out_8_bm[25]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_3_rep2\, B => 
        \data_out_8_bm_1_1[25]_net_1\, C => \line4[57]_net_1\, D
         => \line4[25]_net_1\, Y => \data_out_8_bm[25]_net_1\);
    
    \data_out_8_bm[2]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_3_rep2\, B => 
        \data_out_8_bm_1_1[2]_net_1\, C => \line4[34]_net_1\, D
         => \line4[2]_net_1\, Y => \data_out_8_bm[2]_net_1\);
    
    \line3_5[38]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(6), C => \line3[38]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[38]_net_1\);
    
    \line1[11]\ : SLE
      port map(D => \line1_5[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[11]_net_1\);
    
    \data_out_6_am[18]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[18]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[18]_net_1\, Y => \data_out_6_am[18]_net_1\);
    
    \data_out_8_bm_1_1[19]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[51]_net_1\, B => \line0[19]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[19]_net_1\);
    
    \line0_RNO[29]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(29), C => \line0[29]_net_1\, 
        D => waddr_in_net_0(0), Y => N_38_i_0);
    
    \line2[50]\ : SLE
      port map(D => \line2_5[50]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[50]_net_1\);
    
    \data_out_8_am[7]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[39]_net_1\, D => \line1[7]_net_1\, Y => 
        \data_out_8_am[7]_net_1\);
    
    \line3_5[47]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(15), C => \line3[47]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[47]_net_1\);
    
    \line0[32]\ : SLE
      port map(D => \line0_6[32]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[32]_net_1\);
    
    \line2_5[10]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(10), C => \line2[10]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[10]_net_1\);
    
    \line1_5[60]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(28), C => \line1[60]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[60]_net_1\);
    
    \data_out_9_0_RNO_0[0]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[32]_net_1\, B => \line0[0]_net_1\, C
         => \raddr_pos_3_rep2\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_5_i_m2_1_1[0]\);
    
    \line3_5[8]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(8), C => \line3[8]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[8]_net_1\);
    
    \line1[56]\ : SLE
      port map(D => \line1_5[56]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[56]_net_1\);
    
    \data_out_6_ns[17]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[17]_net_1\, C => \data_out_6_am[17]_net_1\, 
        Y => N_1271);
    
    \line3[36]\ : SLE
      port map(D => \line3_5[36]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[36]_net_1\);
    
    raddr_pos_3_rep2 : SLE
      port map(D => raddr_in_net_0(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_1424_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_3_rep2\);
    
    \line3[4]\ : SLE
      port map(D => \line3_5[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[4]_net_1\);
    
    \line1_5[58]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(26), C => \line1[58]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[58]_net_1\);
    
    \line0[20]\ : SLE
      port map(D => \line0_6[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[20]_net_1\);
    
    \line2_5[12]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(12), C => \line2[12]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[12]_net_1\);
    
    \raddr_pos_fast[3]\ : SLE
      port map(D => raddr_in_net_0(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_1424_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_fast[3]_net_1\);
    
    \line1_5[62]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(30), C => \line1[62]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[62]_net_1\);
    
    \line0[56]\ : SLE
      port map(D => \line0_6[56]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[56]_net_1\);
    
    \line4_5[1]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(1), 
        C => \line4[1]_net_1\, D => N_47_i, Y => 
        \line4_5[1]_net_1\);
    
    \line2[49]\ : SLE
      port map(D => \line2_5[49]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[49]_net_1\);
    
    \data_out_8_ns[11]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[11]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[11]_net_1\, Y
         => N_1332);
    
    \data_out_8_bm[11]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_3_rep2\, B => 
        \data_out_8_bm_1_1[11]_net_1\, C => \line4[43]_net_1\, D
         => \line4[11]_net_1\, Y => \data_out_8_bm[11]_net_1\);
    
    \line2[20]\ : SLE
      port map(D => \line2_5[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[20]_net_1\);
    
    \data_out_8_bm[18]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[18]_net_1\, C => \line4[50]_net_1\, D
         => \line4[18]_net_1\, Y => \data_out_8_bm[18]_net_1\);
    
    \line4_5[56]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(24), 
        C => \line4[56]_net_1\, D => N_47_i, Y => 
        \line4_5[56]_net_1\);
    
    \data_out_8_bm_1_1[18]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[50]_net_1\, B => \line0[18]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[18]_net_1\);
    
    \line3[61]\ : SLE
      port map(D => N_1439_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[61]_net_1\);
    
    \line3[29]\ : SLE
      port map(D => N_1440_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[29]_net_1\);
    
    \line1[54]\ : SLE
      port map(D => \line1_5[54]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[54]_net_1\);
    
    \line3[34]\ : SLE
      port map(D => \line3_5[34]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[34]_net_1\);
    
    \line3[7]\ : SLE
      port map(D => \line3_5[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[7]_net_1\);
    
    \line1_5[25]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(25), C => \line1[25]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[25]_net_1\);
    
    \line0_6[15]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(15), C => \line0[15]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[15]_net_1\);
    
    \line4[61]\ : SLE
      port map(D => N_1437_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[61]_net_1\);
    
    \line0[54]\ : SLE
      port map(D => \line0_6[54]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[54]_net_1\);
    
    \line2_5[38]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(6), C => \line2[38]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[38]_net_1\);
    
    \line0[8]\ : SLE
      port map(D => \line0_6[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[8]_net_1\);
    
    \data_out_8_bm[19]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[19]_net_1\, C => \line4[51]_net_1\, D
         => \line4[19]_net_1\, Y => \data_out_8_bm[19]_net_1\);
    
    \line0[49]\ : SLE
      port map(D => \line0_6[49]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[49]_net_1\);
    
    \data_out_8_am[3]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[35]_net_1\, D => \line1[3]_net_1\, Y => 
        \data_out_8_am[3]_net_1\);
    
    \line3_5[46]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(14), C => \line3[46]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[46]_net_1\);
    
    \line1[51]\ : SLE
      port map(D => \line1_5[51]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[51]_net_1\);
    
    \line4[50]\ : SLE
      port map(D => \line4_5[50]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[50]_net_1\);
    
    \line3[31]\ : SLE
      port map(D => N_20_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD
         => GND_net_1, LAT => GND_net_1, Q => \line3[31]_net_1\);
    
    \line4_5[25]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(25), 
        C => \line4[25]_net_1\, D => N_47_i, Y => 
        \line4_5[25]_net_1\);
    
    \line0[51]\ : SLE
      port map(D => \line0_6[51]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[51]_net_1\);
    
    \line0_6[20]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(20), C => \line0[20]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[20]_net_1\);
    
    \line4_5[3]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(3), 
        C => \line4[3]_net_1\, D => N_47_i, Y => 
        \line4_5[3]_net_1\);
    
    \line2[16]\ : SLE
      port map(D => \line2_5[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[16]_net_1\);
    
    \line0_6[39]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(7), C => \line0[39]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[39]_net_1\);
    
    \line2_5[49]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(17), C => \line2[49]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[49]_net_1\);
    
    ren_pos : SLE
      port map(D => N_35_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ren_pos\);
    
    \line4_5[60]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(28), 
        C => \line4[60]_net_1\, D => N_47_i, Y => 
        \line4_5[60]_net_1\);
    
    \line0_6[22]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(22), C => \line0[22]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[22]_net_1\);
    
    \line1[23]\ : SLE
      port map(D => \line1_5[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[23]_net_1\);
    
    \data_out_8_am[4]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[36]_net_1\, D => \line1[4]_net_1\, Y => 
        \data_out_8_am[4]_net_1\);
    
    \line2_5[53]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(21), C => \line2[53]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[53]_net_1\);
    
    \data_out_8_bm_1_1[24]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[56]_net_1\, B => \line0[24]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[24]_net_1\);
    
    \line4[8]\ : SLE
      port map(D => \line4_5[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[8]_net_1\);
    
    \line3_5[11]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(11), C => \line3[11]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[11]_net_1\);
    
    \line3[55]\ : SLE
      port map(D => \line3_5[55]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[55]_net_1\);
    
    \data_out_6_am[24]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[24]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[24]_net_1\, Y => \data_out_6_am[24]_net_1\);
    
    \line4_5[62]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(30), 
        C => \line4[62]_net_1\, D => N_47_i, Y => 
        \line4_5[62]_net_1\);
    
    \line1_5[0]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(0), C => \line1[0]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[0]_net_1\);
    
    \data_out_8_am[8]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[40]_net_1\, D => \line1[8]_net_1\, Y => 
        \data_out_8_am[8]_net_1\);
    
    \line4[0]\ : SLE
      port map(D => \line4_5[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[0]_net_1\);
    
    \data_out_8_bm_1_1[15]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[47]_net_1\, B => \line0[15]_net_1\, C
         => \raddr_pos_fast[3]_net_1\, D => \raddr_pos[0]_net_1\, 
        Y => \data_out_8_bm_1_1[15]_net_1\);
    
    \line4[42]\ : SLE
      port map(D => \line4_5[42]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[42]_net_1\);
    
    \line2[14]\ : SLE
      port map(D => \line2_5[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[14]_net_1\);
    
    \data_out_8_ns[30]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[30]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[30]_net_1\, Y
         => N_1351);
    
    \data_out_6_am[16]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[16]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[16]_net_1\, Y => \data_out_6_am[16]_net_1\);
    
    \line4_5[11]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(11), 
        C => \line4[11]_net_1\, D => N_47_i, Y => 
        \line4_5[11]_net_1\);
    
    \line1[49]\ : SLE
      port map(D => \line1_5[49]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[49]_net_1\);
    
    \data_out_8_ns[18]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[18]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[18]_net_1\, Y
         => N_1339);
    
    \line2[11]\ : SLE
      port map(D => \line2_5[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[11]_net_1\);
    
    \data_out_6_bm[24]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[56]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[56]_net_1\, Y => \data_out_6_bm[24]_net_1\);
    
    \line3[2]\ : SLE
      port map(D => \line3_5[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[2]_net_1\);
    
    \data_out_8_am[10]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[42]_net_1\, D => \line1[10]_net_1\, Y => 
        \data_out_8_am[10]_net_1\);
    
    \line4[32]\ : SLE
      port map(D => \line4_5[32]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[32]_net_1\);
    
    \line4[16]\ : SLE
      port map(D => \line4_5[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[16]_net_1\);
    
    \line2[32]\ : SLE
      port map(D => \line2_5[32]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[32]_net_1\);
    
    \line4[7]\ : SLE
      port map(D => \line4_5[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[7]_net_1\);
    
    \line2_5[17]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(17), C => \line2[17]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[17]_net_1\);
    
    \data_out_8_bm[20]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[20]_net_1\, C => \line4[52]_net_1\, D
         => \line4[20]_net_1\, Y => \data_out_8_bm[20]_net_1\);
    
    \line3_5[35]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(3), C => \line3[35]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[35]_net_1\);
    
    \line3[9]\ : SLE
      port map(D => \line3_5[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[9]_net_1\);
    
    \line0[33]\ : SLE
      port map(D => \line0_6[33]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[33]_net_1\);
    
    \data_out_8_ns[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[7]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[7]_net_1\, Y
         => N_1328);
    
    \data_out_9_0[1]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_1453, B => data_out_sn_N_11_mux, C => 
        \data_out_sn_N_12_mux\, D => N_1455, Y => data_out_9_0_1);
    
    \line4[1]\ : SLE
      port map(D => \line4_5[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[1]_net_1\);
    
    \line1[35]\ : SLE
      port map(D => \line1_5[35]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[35]_net_1\);
    
    \line3[49]\ : SLE
      port map(D => \line3_5[49]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[49]_net_1\);
    
    \line1_5[20]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(20), C => \line1[20]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[20]_net_1\);
    
    \line0_6[10]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(10), C => \line0[10]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[10]_net_1\);
    
    \line0[12]\ : SLE
      port map(D => \line0_6[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[12]_net_1\);
    
    \data_out_6_am[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[5]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[5]_net_1\, Y => \data_out_6_am[5]_net_1\);
    
    \line4[14]\ : SLE
      port map(D => \line4_5[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[14]_net_1\);
    
    \line1_5[22]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(22), C => \line1[22]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[22]_net_1\);
    
    \line0_6[12]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(12), C => \line0[12]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[12]_net_1\);
    
    \line1_5[55]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(23), C => \line1[55]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[55]_net_1\);
    
    \line1[28]\ : SLE
      port map(D => \line1_5[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[28]_net_1\);
    
    \line4_5[20]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(20), 
        C => \line4[20]_net_1\, D => N_47_i, Y => 
        \line4_5[20]_net_1\);
    
    \line2[4]\ : SLE
      port map(D => \line2_5[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[4]_net_1\);
    
    \data_out_8_bm_1_1[7]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[39]_net_1\, B => \line0[7]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[7]_net_1\);
    
    \line4[11]\ : SLE
      port map(D => \line4_5[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[11]_net_1\);
    
    \line4_5[39]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(7), 
        C => \line4[39]_net_1\, D => N_47_i, Y => 
        \line4_5[39]_net_1\);
    
    \line4_5[22]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(22), 
        C => \line4[22]_net_1\, D => N_47_i, Y => 
        \line4_5[22]_net_1\);
    
    \line2_5[16]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(16), C => \line2[16]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[16]_net_1\);
    
    \data_out_6_am[25]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[25]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[25]_net_1\, Y => \data_out_6_am[25]_net_1\);
    
    \data_out_6_am[22]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[22]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[22]_net_1\, Y => \data_out_6_am[22]_net_1\);
    
    \line4_RNO[29]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(29), 
        C => \line4[29]_net_1\, D => N_47_i, Y => N_1438_i_0);
    
    \data_out_6_ns[23]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[23]_net_1\, C => \data_out_6_am[23]_net_1\, 
        Y => N_1277);
    
    \data_out_8_ns[20]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[20]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[20]_net_1\, Y
         => N_1341);
    
    \data_out_8_ns[19]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[19]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[19]_net_1\, Y
         => N_1340);
    
    \line1[19]\ : SLE
      port map(D => \line1_5[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[19]_net_1\);
    
    \line2_5[35]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(3), C => \line2[35]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[35]_net_1\);
    
    \line0_6[27]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(27), C => \line0[27]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[27]_net_1\);
    
    \line1[0]\ : SLE
      port map(D => \line1_5[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[0]_net_1\);
    
    \data_out_6_ns[12]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[12]_net_1\, C => \data_out_6_am[12]_net_1\, 
        Y => N_1266);
    
    \line4[20]\ : SLE
      port map(D => \line4_5[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[20]_net_1\);
    
    \line2[55]\ : SLE
      port map(D => \line2_5[55]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[55]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line3[1]\ : SLE
      port map(D => \line3_5[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[1]_net_1\);
    
    \line0[38]\ : SLE
      port map(D => \line0_6[38]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[38]_net_1\);
    
    \line2[47]\ : SLE
      port map(D => \line2_5[47]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[47]_net_1\);
    
    \line0[25]\ : SLE
      port map(D => \line0_6[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[25]_net_1\);
    
    \data_out_6_bm[9]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[41]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[41]_net_1\, Y => \data_out_6_bm[9]_net_1\);
    
    \line2_5[58]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(26), C => \line2[58]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[58]_net_1\);
    
    \data_out_6_ns[21]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[21]_net_1\, C => \data_out_6_am[21]_net_1\, 
        Y => N_1275);
    
    \line3[27]\ : SLE
      port map(D => \line3_5[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[27]_net_1\);
    
    \data_out_6_am[10]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[10]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[10]_net_1\, Y => \data_out_6_am[10]_net_1\);
    
    \line3_5[30]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(30), C => \line3[30]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[30]_net_1\);
    
    \line2[25]\ : SLE
      port map(D => \line2_5[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[25]_net_1\);
    
    N_1424_i : CFG2
      generic map(INIT => x"B")

      port map(A => AHB_slave_dummy_0_read_en, B => 
        sha256_system_sb_0_POWER_ON_RESET_N, Y => N_1424_i_0);
    
    \line4[43]\ : SLE
      port map(D => \line4_5[43]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[43]_net_1\);
    
    \data_out_8_bm[7]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[7]_net_1\, C => \line4[39]_net_1\, D
         => \line4[7]_net_1\, Y => \data_out_8_bm[7]_net_1\);
    
    \line3[12]\ : SLE
      port map(D => \line3_5[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[12]_net_1\);
    
    \line3_5[32]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(0), C => \line3[32]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[32]_net_1\);
    
    \line0[47]\ : SLE
      port map(D => \line0_6[47]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[47]_net_1\);
    
    \line3_5[13]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(13), C => \line3[13]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[13]_net_1\);
    
    \data_out_6_ns[9]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[9]_net_1\, C => \data_out_6_am[9]_net_1\, 
        Y => N_1263);
    
    \line4_5[54]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(22), 
        C => \line4[54]_net_1\, D => N_47_i, Y => 
        \line4_5[54]_net_1\);
    
    \line0_6[26]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(26), C => \line0[26]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[26]_net_1\);
    
    \line3_5[5]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(5), C => \line3[5]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[5]_net_1\);
    
    \line4[33]\ : SLE
      port map(D => \line4_5[33]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[33]_net_1\);
    
    \line2[33]\ : SLE
      port map(D => \line2_5[33]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[33]_net_1\);
    
    \line1_5[50]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(18), C => \line1[50]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[50]_net_1\);
    
    \data_out_6_am[28]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[28]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[28]_net_1\, Y => \data_out_6_am[28]_net_1\);
    
    \line4[55]\ : SLE
      port map(D => \line4_5[55]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[55]_net_1\);
    
    \line1[59]\ : SLE
      port map(D => \line1_5[59]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[59]_net_1\);
    
    \line4_5[13]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(13), 
        C => \line4[13]_net_1\, D => N_47_i, Y => 
        \line4_5[13]_net_1\);
    
    \line3[39]\ : SLE
      port map(D => \line3_5[39]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[39]_net_1\);
    
    \data_out_8_bm_1_1[11]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[43]_net_1\, B => \line0[11]_net_1\, C
         => \raddr_pos_fast[3]_net_1\, D => \raddr_pos[0]_net_1\, 
        Y => \data_out_8_bm_1_1[11]_net_1\);
    
    \line1_5[52]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(20), C => \line1[52]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[52]_net_1\);
    
    \line1_5[27]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(27), C => \line1[27]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[27]_net_1\);
    
    \line3_5[44]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(12), C => \line3[44]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[44]_net_1\);
    
    \line0_6[17]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(17), C => \line0[17]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[17]_net_1\);
    
    \line0[59]\ : SLE
      port map(D => \line0_6[59]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[59]_net_1\);
    
    \line0[13]\ : SLE
      port map(D => \line0_6[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[13]_net_1\);
    
    \data_out_8_bm[30]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[30]_net_1\, C => \line4[62]_net_1\, D
         => \line4[30]_net_1\, Y => \data_out_8_bm[30]_net_1\);
    
    \data_out_8_bm_1_1[26]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[58]_net_1\, B => \line0[26]_net_1\, C
         => \raddr_pos_3_rep2\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[26]_net_1\);
    
    \data_out_8_ns[14]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[14]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[14]_net_1\, Y
         => N_1335);
    
    \line3_5[2]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(2), C => \line3[2]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[2]_net_1\);
    
    \data_out_8_bm[3]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[3]_net_1\, C => \line4[35]_net_1\, D
         => \line4[3]_net_1\, Y => \data_out_8_bm[3]_net_1\);
    
    \line1[9]\ : SLE
      port map(D => \line1_5[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[9]_net_1\);
    
    \line4_5[27]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(27), 
        C => \line4[27]_net_1\, D => N_47_i, Y => 
        \line4_5[27]_net_1\);
    
    \data_out_6_am[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[2]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[2]_net_1\, Y => \data_out_6_am[2]_net_1\);
    
    \data_out_8_bm_1_1[9]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[41]_net_1\, B => \line0[9]_net_1\, C
         => \raddr_pos_fast[3]_net_1\, D => \raddr_pos[0]_net_1\, 
        Y => \data_out_8_bm_1_1[9]_net_1\);
    
    \data_out_6_bm[18]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[50]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[50]_net_1\, Y => \data_out_6_bm[18]_net_1\);
    
    \line2_5[30]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(30), C => \line2[30]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[30]_net_1\);
    
    \data_out_8_bm[21]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[21]_net_1\, C => \line4[53]_net_1\, D
         => \line4[21]_net_1\, Y => \data_out_8_bm[21]_net_1\);
    
    \line3[5]\ : SLE
      port map(D => \line3_5[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[5]_net_1\);
    
    \line3[8]\ : SLE
      port map(D => \line3_5[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[8]_net_1\);
    
    \data_out_8_bm[28]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[28]_net_1\, C => \line4[60]_net_1\, D
         => \line4[28]_net_1\, Y => \data_out_8_bm[28]_net_1\);
    
    \line2_5[32]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(0), C => \line2[32]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[32]_net_1\);
    
    \line1[47]\ : SLE
      port map(D => \line1_5[47]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[47]_net_1\);
    
    \line1[7]\ : SLE
      port map(D => \line1_5[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[7]_net_1\);
    
    \line1[60]\ : SLE
      port map(D => \line1_5[60]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[60]_net_1\);
    
    \line4[48]\ : SLE
      port map(D => \line4_5[48]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[48]_net_1\);
    
    \line0[62]\ : SLE
      port map(D => \line0_6[62]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[62]_net_1\);
    
    \line1_5[7]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(7), C => \line1[7]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[7]_net_1\);
    
    \line1_5[19]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(19), C => \line1[19]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[19]_net_1\);
    
    \line1_5[39]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(7), C => \line1[39]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[39]_net_1\);
    
    \data_out_8_bm[4]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[4]_net_1\, C => \line4[36]_net_1\, D
         => \line4[4]_net_1\, Y => \data_out_8_bm[4]_net_1\);
    
    \data_out_9_m2_1_am[31]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[31]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[31]_net_1\, Y => 
        \data_out_9_m2_1_am[31]_net_1\);
    
    \line1_5[26]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(26), C => \line1[26]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[26]_net_1\);
    
    \line2[6]\ : SLE
      port map(D => \line2_5[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[6]_net_1\);
    
    \line0_6[16]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(16), C => \line0[16]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[16]_net_1\);
    
    \data_out_9_a4_1_1[31]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \raddr_pos_fast[3]_net_1\, B => \ren_pos\, Y
         => N_1423_1);
    
    \line2[19]\ : SLE
      port map(D => \line2_5[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[19]_net_1\);
    
    \line2_5[2]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(2), C => \line2[2]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[2]_net_1\);
    
    \data_out_8_bm[8]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[8]_net_1\, C => \line4[40]_net_1\, D
         => \line4[8]_net_1\, Y => \data_out_8_bm[8]_net_1\);
    
    \line3_5[59]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(27), C => \line3[59]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[59]_net_1\);
    
    \line2_RNO[63]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(31), C => \line2[63]_net_1\, 
        D => waddr_in_net_0(0), Y => N_22_i_0);
    
    un1_wen_19_or_0_m2 : CFG3
      generic map(INIT => x"D8")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(3), C
         => waddr_in_net_0(2), Y => N_61);
    
    \line4[38]\ : SLE
      port map(D => \line4_5[38]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[38]_net_1\);
    
    \line3[47]\ : SLE
      port map(D => \line3_5[47]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[47]_net_1\);
    
    \line2[38]\ : SLE
      port map(D => \line2_5[38]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[38]_net_1\);
    
    \line0_6[49]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(17), C => \line0[49]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[49]_net_1\);
    
    \line4_5[26]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(26), 
        C => \line4[26]_net_1\, D => N_47_i, Y => 
        \line4_5[26]_net_1\);
    
    \line2_5[41]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(9), C => \line2[41]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[41]_net_1\);
    
    \data_out_9_a4_1_3[31]\ : CFG4
      generic map(INIT => x"2400")

      port map(A => \raddr_pos[2]_net_1\, B => 
        \raddr_pos[1]_net_1\, C => \raddr_pos[0]_net_1\, D => 
        N_1423_1, Y => N_1423_3);
    
    \line4_5[0]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(0), 
        C => \line4[0]_net_1\, D => N_47_i, Y => 
        \line4_5[0]_net_1\);
    
    \data_out_8_bm[17]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[17]_net_1\, C => \line4[49]_net_1\, D
         => \line4[17]_net_1\, Y => \data_out_8_bm[17]_net_1\);
    
    \line3_5[37]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(5), C => \line3[37]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[37]_net_1\);
    
    \line0[18]\ : SLE
      port map(D => \line0_6[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[18]_net_1\);
    
    \line1_5[49]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(17), C => \line1[49]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[49]_net_1\);
    
    \line2[3]\ : SLE
      port map(D => \line2_5[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[3]_net_1\);
    
    \data_out_6_ns[14]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[14]_net_1\, C => \data_out_6_am[14]_net_1\, 
        Y => N_1268);
    
    \data_out_6_bm[15]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[47]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[47]_net_1\, Y => \data_out_6_bm[15]_net_1\);
    
    \line3[13]\ : SLE
      port map(D => \line3_5[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[13]_net_1\);
    
    \data_out_9_m2_0_ns[29]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_9_m2_0_bm[29]_net_1\, C => 
        \data_out_9_m2_0_am[29]_net_1\, Y => N_1467);
    
    \line2_5[55]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(23), C => \line2[55]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[55]_net_1\);
    
    \line1[26]\ : SLE
      port map(D => \line1_5[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[26]_net_1\);
    
    \data_out_6_am[17]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[17]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[17]_net_1\, Y => \data_out_6_am[17]_net_1\);
    
    \data_out_6_am[13]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[13]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[13]_net_1\, Y => \data_out_6_am[13]_net_1\);
    
    \line4_5[49]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(17), 
        C => \line4[49]_net_1\, D => N_47_i, Y => 
        \line4_5[49]_net_1\);
    
    \line4[19]\ : SLE
      port map(D => \line4_5[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[19]_net_1\);
    
    \line3_5[18]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(18), C => \line3[18]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[18]_net_1\);
    
    \line1_5[57]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(25), C => \line1[57]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[57]_net_1\);
    
    \data_out_6_am[26]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[26]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[26]_net_1\, Y => \data_out_6_am[26]_net_1\);
    
    \line1[17]\ : SLE
      port map(D => \line1_5[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[17]_net_1\);
    
    \data_out_8_ns[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[3]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[3]_net_1\, Y
         => N_1324);
    
    \data_out_8_am[20]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[52]_net_1\, D => \line1[20]_net_1\, Y => 
        \data_out_8_am[20]_net_1\);
    
    \line2_5[14]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(14), C => \line2[14]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[14]_net_1\);
    
    \line3_5[3]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(3), C => \line3[3]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[3]_net_1\);
    
    \line4_5[18]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(18), 
        C => \line4[18]_net_1\, D => N_47_i, Y => 
        \line4_5[18]_net_1\);
    
    \line4[25]\ : SLE
      port map(D => \line4_5[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[25]_net_1\);
    
    \line3[52]\ : SLE
      port map(D => \line3_5[52]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[52]_net_1\);
    
    \line1[24]\ : SLE
      port map(D => \line1_5[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[24]_net_1\);
    
    \line3_5[36]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(4), C => \line3[36]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[36]_net_1\);
    
    \data_out_8_am[14]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[46]_net_1\, D => \line1[14]_net_1\, Y => 
        \data_out_8_am[14]_net_1\);
    
    \line2_5[37]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(5), C => \line2[37]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[37]_net_1\);
    
    \line1[21]\ : SLE
      port map(D => \line1_5[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[21]_net_1\);
    
    \data_out_8_ns[8]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[8]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[8]_net_1\, Y
         => N_1329);
    
    \line0[36]\ : SLE
      port map(D => \line0_6[36]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[36]_net_1\);
    
    \line3_5[60]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(28), C => \line3[60]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[60]_net_1\);
    
    \line1_5[56]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(24), C => \line1[56]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[56]_net_1\);
    
    \data_out_8_am[9]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[41]_net_1\, D => \line1[9]_net_1\, Y => 
        \data_out_8_am[9]_net_1\);
    
    \line1[2]\ : SLE
      port map(D => \line1_5[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[2]_net_1\);
    
    \line3_5[62]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(30), C => \line3[62]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[62]_net_1\);
    
    \line0[63]\ : SLE
      port map(D => N_30_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => un1_wen_7_or, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[63]_net_1\);
    
    \line3[18]\ : SLE
      port map(D => \line3_5[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[18]_net_1\);
    
    \line1[32]\ : SLE
      port map(D => \line1_5[32]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[32]_net_1\);
    
    \data_out_9_m2_1_ns[31]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_9_m2_1_bm[31]_net_1\, C => 
        \data_out_9_m2_1_am[31]_net_1\, Y => N_60);
    
    \line1[57]\ : SLE
      port map(D => \line1_5[57]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[57]_net_1\);
    
    \line0[34]\ : SLE
      port map(D => \line0_6[34]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[34]_net_1\);
    
    \line3[37]\ : SLE
      port map(D => \line3_5[37]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[37]_net_1\);
    
    \data_out_8_ns[17]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[17]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[17]_net_1\, Y
         => N_1338);
    
    \line0[57]\ : SLE
      port map(D => \line0_6[57]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[57]_net_1\);
    
    \line0_6[24]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(24), C => \line0[24]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[24]_net_1\);
    
    \data_out_8_am[11]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[43]_net_1\, D => \line1[11]_net_1\, Y => 
        \data_out_8_am[11]_net_1\);
    
    \data_out_8_am[15]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[47]_net_1\, D => \line1[15]_net_1\, Y => 
        \data_out_8_am[15]_net_1\);
    
    \line2_5[50]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(18), C => \line2[50]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[50]_net_1\);
    
    \line2_5[36]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(4), C => \line2[36]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[36]_net_1\);
    
    \line1_RNO[61]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(29), C => \line1[61]_net_1\, 
        D => waddr_in_net_0(0), Y => N_1443_i_0);
    
    \line0[31]\ : SLE
      port map(D => N_32_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => un1_wen_7_or, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[31]_net_1\);
    
    \line2_5[52]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(20), C => \line2[52]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[52]_net_1\);
    
    \line0_6[59]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(27), C => \line0[59]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[59]_net_1\);
    
    \data_out_6_ns[19]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[19]_net_1\, C => \data_out_6_am[19]_net_1\, 
        Y => N_1273);
    
    \line0_6[33]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(1), C => \line0[33]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[33]_net_1\);
    
    \data_out_6_bm[17]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[49]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[49]_net_1\, Y => \data_out_6_bm[17]_net_1\);
    
    \line2_5[43]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(11), C => \line2[43]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[43]_net_1\);
    
    \line2[7]\ : SLE
      port map(D => \line2_5[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[7]_net_1\);
    
    \line0_6[3]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(3), C => \line0[3]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[3]_net_1\);
    
    \data_out_8_am[16]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[48]_net_1\, D => \line1[16]_net_1\, Y => 
        \data_out_8_am[16]_net_1\);
    
    \data_out_6_am[20]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[20]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[20]_net_1\, Y => \data_out_6_am[20]_net_1\);
    
    \data_out_8_ns[26]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[26]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[26]_net_1\, Y
         => N_1347);
    
    \line4[6]\ : SLE
      port map(D => \line4_5[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[6]_net_1\);
    
    \data_out_8_bm[16]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[16]_net_1\, C => \line4[48]_net_1\, D
         => \line4[16]_net_1\, Y => \data_out_8_bm[16]_net_1\);
    
    \line2[52]\ : SLE
      port map(D => \line2_5[52]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[52]_net_1\);
    
    \line2[17]\ : SLE
      port map(D => \line2_5[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[17]_net_1\);
    
    \line4_5_1_o2[63]\ : CFG3
      generic map(INIT => x"64")

      port map(A => waddr_in_net_0(3), B => N_44, C => 
        waddr_in_net_0(0), Y => N_46);
    
    \line4[46]\ : SLE
      port map(D => \line4_5[46]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[46]_net_1\);
    
    \line0[22]\ : SLE
      port map(D => \line0_6[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[22]_net_1\);
    
    \line3_5[15]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(15), C => \line3[15]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[15]_net_1\);
    
    \line3[53]\ : SLE
      port map(D => \line3_5[53]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[53]_net_1\);
    
    \line1_5[24]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(24), C => \line1[24]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[24]_net_1\);
    
    \line0_6[14]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(14), C => \line0[14]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[14]_net_1\);
    
    \data_out_6_am[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[7]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[7]_net_1\, Y => \data_out_6_am[7]_net_1\);
    
    \data_out_8_am[30]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[62]_net_1\, D => \line1[30]_net_1\, Y => 
        \data_out_8_am[30]_net_1\);
    
    \line2[22]\ : SLE
      port map(D => \line2_5[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[22]_net_1\);
    
    \line4[36]\ : SLE
      port map(D => \line4_5[36]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[36]_net_1\);
    
    \line2[36]\ : SLE
      port map(D => \line2_5[36]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[36]_net_1\);
    
    \line4_5[15]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(15), 
        C => \line4[15]_net_1\, D => N_47_i, Y => 
        \line4_5[15]_net_1\);
    
    \line2[2]\ : SLE
      port map(D => \line2_5[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[2]_net_1\);
    
    \line1_5[1]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(1), C => \line1[1]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[1]_net_1\);
    
    \line4[9]\ : SLE
      port map(D => \line4_5[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[9]_net_1\);
    
    \line4_5[24]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(24), 
        C => \line4[24]_net_1\, D => N_47_i, Y => 
        \line4_5[24]_net_1\);
    
    \line4[44]\ : SLE
      port map(D => \line4_5[44]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[44]_net_1\);
    
    \line2_5[6]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(6), C => \line2[6]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[6]_net_1\);
    
    \data_out_6_bm[28]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[60]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[60]_net_1\, Y => \data_out_6_bm[28]_net_1\);
    
    un1_wen_4_or_0 : CFG3
      generic map(INIT => x"8F")

      port map(A => N_1434, B => waddr_in_net_0(3), C => 
        sha256_system_sb_0_POWER_ON_RESET_N, Y => un1_wen_4_or);
    
    \data_out_6_ns[7]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[7]_net_1\, C => \data_out_6_am[7]_net_1\, 
        Y => N_1261);
    
    \line0[16]\ : SLE
      port map(D => \line0_6[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[16]_net_1\);
    
    \line2_RNO[29]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(29), C => \line2[29]_net_1\, 
        D => waddr_in_net_0(0), Y => N_1442_i_0);
    
    \line4[17]\ : SLE
      port map(D => \line4_5[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[17]_net_1\);
    
    \line4[41]\ : SLE
      port map(D => \line4_5[41]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[41]_net_1\);
    
    \line2[40]\ : SLE
      port map(D => \line2_5[40]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[40]_net_1\);
    
    \line4[52]\ : SLE
      port map(D => \line4_5[52]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[52]_net_1\);
    
    \data_out_6_bm[19]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[51]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[51]_net_1\, Y => \data_out_6_bm[19]_net_1\);
    
    \line3_RNO[29]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(29), C => \line3[29]_net_1\, 
        D => waddr_in_net_0(0), Y => N_1440_i_0);
    
    \line4[34]\ : SLE
      port map(D => \line4_5[34]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[34]_net_1\);
    
    \line0[0]\ : SLE
      port map(D => \line0_6[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[0]_net_1\);
    
    \line2[34]\ : SLE
      port map(D => \line2_5[34]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[34]_net_1\);
    
    \line1_5[11]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(11), C => \line1[11]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[11]_net_1\);
    
    \line1[33]\ : SLE
      port map(D => \line1_5[33]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[33]_net_1\);
    
    \line3[20]\ : SLE
      port map(D => \line3_5[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[20]_net_1\);
    
    \data_out_6_am[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[3]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[3]_net_1\, Y => \data_out_6_am[3]_net_1\);
    
    \line4_5[33]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(1), 
        C => \line4[33]_net_1\, D => N_47_i, Y => 
        \line4_5[33]_net_1\);
    
    \line4[31]\ : SLE
      port map(D => \line4_5[31]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[31]_net_1\);
    
    \line2_5[57]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(25), C => \line2[57]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[57]_net_1\);
    
    \line2[31]\ : SLE
      port map(D => N_24_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => un1_wen_19_or, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[31]_net_1\);
    
    \line3_5[51]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(19), C => \line3[51]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[51]_net_1\);
    
    \line0[14]\ : SLE
      port map(D => \line0_6[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[14]_net_1\);
    
    \data_out_9_0_RNO_0[31]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[63]_net_1\, B => \line0[31]_net_1\, C
         => \raddr_pos_fast[3]_net_1\, D => \raddr_pos[0]_net_1\, 
        Y => \data_out_9_m2_0_1_1[31]\);
    
    \data_out_6_bm[12]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[44]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[44]_net_1\, Y => \data_out_6_bm[12]_net_1\);
    
    \line0[40]\ : SLE
      port map(D => \line0_6[40]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[40]_net_1\);
    
    \line0_6[41]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(9), C => \line0[41]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[41]_net_1\);
    
    \data_out_8_bm_1_1[28]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[60]_net_1\, B => \line0[28]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[28]_net_1\);
    
    \line4_5[2]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(2), 
        C => \line4[2]_net_1\, D => N_47_i, Y => 
        \line4_5[2]_net_1\);
    
    un1_wen_20_or_0 : CFG3
      generic map(INIT => x"D5")

      port map(A => sha256_system_sb_0_POWER_ON_RESET_N, B => 
        N_1434, C => N_62, Y => un1_wen_20_or);
    
    \line3[58]\ : SLE
      port map(D => \line3_5[58]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[58]_net_1\);
    
    \line0[11]\ : SLE
      port map(D => \line0_6[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[11]_net_1\);
    
    \data_out_9_0[31]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_56, B => \data_out_sn_N_12_mux\, C => 
        data_out_sn_N_11_mux, D => N_60, Y => data_out_9_0_31);
    
    \data_out_8_bm[27]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[27]_net_1\, C => \line4[59]_net_1\, D
         => \line4[27]_net_1\, Y => \data_out_8_bm[27]_net_1\);
    
    \line3_5[34]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(2), C => \line3[34]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[34]_net_1\);
    
    \line1_5[41]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(9), C => \line1[41]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[41]_net_1\);
    
    \data_out_6_am[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[4]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[4]_net_1\, Y => \data_out_6_am[4]_net_1\);
    
    \line3_5[10]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(10), C => \line3[10]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[10]_net_1\);
    
    \line0_6[38]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(6), C => \line0[38]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[38]_net_1\);
    
    \line1[29]\ : SLE
      port map(D => N_34_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => un1_wen_20_or, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[29]_net_1\);
    
    \line2_5[48]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(16), C => \line2[48]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[48]_net_1\);
    
    \line2[60]\ : SLE
      port map(D => \line2_5[60]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[60]_net_1\);
    
    \line2_5[9]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(9), C => \line2[9]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[9]_net_1\);
    
    \data_out_6_am[8]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[8]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[8]_net_1\, Y => \data_out_6_am[8]_net_1\);
    
    \line3_5[0]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(0), C => \line3[0]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[0]_net_1\);
    
    \data_out_6_bm[25]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[57]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[57]_net_1\, Y => \data_out_6_bm[25]_net_1\);
    
    \line3_5[12]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(12), C => \line3[12]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[12]_net_1\);
    
    \line2[53]\ : SLE
      port map(D => \line2_5[53]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[53]_net_1\);
    
    \line1_5[6]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(6), C => \line1[6]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[6]_net_1\);
    
    \line1[8]\ : SLE
      port map(D => \line1_5[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[8]_net_1\);
    
    \data_out_6_am[30]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[30]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[30]_net_1\, Y => \data_out_6_am[30]_net_1\);
    
    \line4_5[41]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(9), 
        C => \line4[41]_net_1\, D => N_47_i, Y => 
        \line4_5[41]_net_1\);
    
    \line2_5[56]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(24), C => \line2[56]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[56]_net_1\);
    
    \data_out_6_am[27]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[27]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[27]_net_1\, Y => \data_out_6_am[27]_net_1\);
    
    \data_out_6_am[23]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[23]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[23]_net_1\, Y => \data_out_6_am[23]_net_1\);
    
    \line1_5[4]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(4), C => \line1[4]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[4]_net_1\);
    
    \line4_5[10]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(10), 
        C => \line4[10]_net_1\, D => N_47_i, Y => 
        \line4_5[10]_net_1\);
    
    \line1_5[54]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(22), C => \line1[54]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[54]_net_1\);
    
    \data_out_8_ns[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[2]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[2]_net_1\, Y
         => N_1323);
    
    \data_out_9_0_RNO[29]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_9_m2_1_1_1[29]\, C => \line0[61]_net_1\, D => 
        \line0[29]_net_1\, Y => N_1468);
    
    \line0[23]\ : SLE
      port map(D => \line0_6[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[23]_net_1\);
    
    \line3[16]\ : SLE
      port map(D => \line3_5[16]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[16]_net_1\);
    
    \line4_5[12]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(12), 
        C => \line4[12]_net_1\, D => N_47_i, Y => 
        \line4_5[12]_net_1\);
    
    \line1[38]\ : SLE
      port map(D => \line1_5[38]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[38]_net_1\);
    
    \line1[40]\ : SLE
      port map(D => \line1_5[40]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[40]_net_1\);
    
    \data_out_8_bm[9]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_3_rep2\, B => 
        \data_out_8_bm_1_1[9]_net_1\, C => \line4[41]_net_1\, D
         => \line4[9]_net_1\, Y => \data_out_8_bm[9]_net_1\);
    
    \data_out_6_ns[13]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[13]_net_1\, C => \data_out_6_am[13]_net_1\, 
        Y => N_1267);
    
    \data_out_8_ns[10]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[10]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[10]_net_1\, Y
         => N_1331);
    
    \line2_5[1]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(1), C => \line2[1]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[1]_net_1\);
    
    \line2[23]\ : SLE
      port map(D => \line2_5[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[23]_net_1\);
    
    \data_out_8_bm_1_1[25]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[57]_net_1\, B => \line0[25]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[25]_net_1\);
    
    \line2_5[5]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(5), C => \line2[5]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[5]_net_1\);
    
    \line0[39]\ : SLE
      port map(D => \line0_6[39]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[39]_net_1\);
    
    \line2_5[34]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(2), C => \line2[34]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[34]_net_1\);
    
    \data_out_8_am[24]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[56]_net_1\, D => \line1[24]_net_1\, Y => 
        \data_out_8_am[24]_net_1\);
    
    \line3[14]\ : SLE
      port map(D => \line3_5[14]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[14]_net_1\);
    
    un1_wen_7_or_0_a2 : CFG2
      generic map(INIT => x"4")

      port map(A => AHB_slave_dummy_0_read_en, B => 
        AHB_slave_dummy_0_write_en, Y => N_1434);
    
    \line3[40]\ : SLE
      port map(D => \line3_5[40]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[40]_net_1\);
    
    \data_out_9_0[0]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_1454, B => data_out_sn_N_11_mux, C => 
        \data_out_sn_N_12_mux\, D => N_1456, Y => data_out_9_0_0);
    
    \line3_RNO[61]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(29), C => \line3[61]_net_1\, 
        D => waddr_in_net_0(0), Y => N_1439_i_0);
    
    \data_out_9_m2[31]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[31]_net_1\, B => \raddr_pos[0]_net_1\, 
        C => \line2[63]_net_1\, Y => N_53);
    
    \data_out_8_bm_1_1[12]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[44]_net_1\, B => \line0[12]_net_1\, C
         => \raddr_pos_3_rep2\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[12]_net_1\);
    
    \data_out_6_bm[10]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[42]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[42]_net_1\, Y => \data_out_6_bm[10]_net_1\);
    
    \data_out_6_ns[11]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[11]_net_1\, C => \data_out_6_am[11]_net_1\, 
        Y => N_1265);
    
    \data_out_6_am[19]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[19]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[19]_net_1\, Y => \data_out_6_am[19]_net_1\);
    
    \line4[53]\ : SLE
      port map(D => \line4_5[53]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[53]_net_1\);
    
    \line3[11]\ : SLE
      port map(D => \line3_5[11]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[11]_net_1\);
    
    \data_out_4_i_m2[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[1]_net_1\, B => \raddr_pos[0]_net_1\, 
        C => \line2[33]_net_1\, Y => N_1457);
    
    \line4_RNO[61]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(29), 
        C => \line4[61]_net_1\, D => N_47_i, Y => N_1437_i_0);
    
    \line4[22]\ : SLE
      port map(D => \line4_5[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[22]_net_1\);
    
    \line2_5[21]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(21), C => \line2[21]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[21]_net_1\);
    
    \line2[58]\ : SLE
      port map(D => \line2_5[58]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[58]_net_1\);
    
    \data_out_8_bm_1_1[2]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[34]_net_1\, B => \line0[2]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[2]_net_1\);
    
    \line4_5[38]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(6), 
        C => \line4[38]_net_1\, D => N_47_i, Y => 
        \line4_5[38]_net_1\);
    
    \line1_5[13]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(13), C => \line1[13]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[13]_net_1\);
    
    \line2[8]\ : SLE
      port map(D => \line2_5[8]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[8]_net_1\);
    
    \line1_RNO[31]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(31), C => \line1[31]_net_1\, 
        D => waddr_in_net_0(0), Y => N_28_i_0);
    
    \line1_5[33]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(1), C => \line1[33]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[33]_net_1\);
    
    \data_out_8_ns[23]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[23]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[23]_net_1\, Y
         => N_1344);
    
    \line0[28]\ : SLE
      port map(D => \line0_6[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[28]_net_1\);
    
    \data_out_8_bm_1_1[3]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[35]_net_1\, B => \line0[3]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[3]_net_1\);
    
    \data_out_8_am[21]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[53]_net_1\, D => \line1[21]_net_1\, Y => 
        \data_out_8_am[21]_net_1\);
    
    \data_out_8_am[25]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[57]_net_1\, D => \line1[25]_net_1\, Y => 
        \data_out_8_am[25]_net_1\);
    
    \data_out_8_bm_1_1[30]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[62]_net_1\, B => \line0[30]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[30]_net_1\);
    
    \line1[10]\ : SLE
      port map(D => \line1_5[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[10]_net_1\);
    
    \data_out_8_ns[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[4]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[4]_net_1\, Y
         => N_1325);
    
    \line3_5[53]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(21), C => \line3[53]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[53]_net_1\);
    
    \line4_5_1[63]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(31), 
        C => \line4[63]_net_1\, D => N_46, Y => \line4_5[63]\);
    
    \line3_5[17]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(17), C => \line3[17]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[17]_net_1\);
    
    \line2[28]\ : SLE
      port map(D => \line2_5[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[28]_net_1\);
    
    \line0_6[51]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(19), C => \line0[51]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[51]_net_1\);
    
    \line0_6[43]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(11), C => \line0[43]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[43]_net_1\);
    
    \line0_RNO[61]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(29), C => \line0[61]_net_1\, 
        D => waddr_in_net_0(0), Y => N_36_i_0);
    
    \line0[6]\ : SLE
      port map(D => \line0_6[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[6]_net_1\);
    
    \data_out_6_bm[27]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[59]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[59]_net_1\, Y => \data_out_6_bm[27]_net_1\);
    
    \line0_6[2]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(2), C => \line0[2]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[2]_net_1\);
    
    \data_out_8_am[26]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[58]_net_1\, D => \line1[26]_net_1\, Y => 
        \data_out_8_am[26]_net_1\);
    
    un1_wen_18_or_0_0 : CFG4
      generic map(INIT => x"B333")

      port map(A => waddr_in_net_0(2), B => 
        sha256_system_sb_0_POWER_ON_RESET_N, C => N_1434, D => 
        waddr_in_net_0(1), Y => \un1_wen_18_or_0_0\);
    
    \data_out_8_am[12]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[44]_net_1\, D => \line1[12]_net_1\, Y => 
        \data_out_8_am[12]_net_1\);
    
    \line1_5[43]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(11), C => \line1[43]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[43]_net_1\);
    
    \line4_5[17]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(17), 
        C => \line4[17]_net_1\, D => N_47_i, Y => 
        \line4_5[17]_net_1\);
    
    \data_out_8_bm[26]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[26]_net_1\, C => \line4[58]_net_1\, D
         => \line4[26]_net_1\, Y => \data_out_8_bm[26]_net_1\);
    
    \line0_6[35]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(3), C => \line0[35]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[35]_net_1\);
    
    \line2[1]\ : SLE
      port map(D => \line2_5[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[1]_net_1\);
    
    \line2_5[45]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(13), C => \line2[45]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[45]_net_1\);
    
    \line2[45]\ : SLE
      port map(D => \line2_5[45]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[45]_net_1\);
    
    \line4[49]\ : SLE
      port map(D => \line4_5[49]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[49]_net_1\);
    
    \line0[61]\ : SLE
      port map(D => N_36_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => un1_wen_7_or, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[61]_net_1\);
    
    \data_out_6_i_m2_bm[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[33]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[33]_net_1\, Y => 
        \data_out_6_i_m2_bm[1]_net_1\);
    
    \line4[58]\ : SLE
      port map(D => \line4_5[58]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[58]_net_1\);
    
    \line3_RNO[31]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(31), C => \line3[31]_net_1\, 
        D => waddr_in_net_0(0), Y => N_20_i_0);
    
    \line3[25]\ : SLE
      port map(D => \line3_5[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[25]_net_1\);
    
    \line3[60]\ : SLE
      port map(D => \line3_5[60]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[60]_net_1\);
    
    \line4_5[59]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(27), 
        C => \line4[59]_net_1\, D => N_47_i, Y => 
        \line4_5[59]_net_1\);
    
    \line4_5[43]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(11), 
        C => \line4[43]_net_1\, D => N_47_i, Y => 
        \line4_5[43]_net_1\);
    
    \line3_5[21]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(21), C => \line3[21]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[21]_net_1\);
    
    \data_out_9_m2[29]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[29]_net_1\, B => \raddr_pos[0]_net_1\, 
        C => \line2[61]_net_1\, Y => N_1446);
    
    \line4[39]\ : SLE
      port map(D => \line4_5[39]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[39]_net_1\);
    
    \line2[39]\ : SLE
      port map(D => \line2_5[39]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[39]_net_1\);
    
    \data_out_8_am[13]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[45]_net_1\, D => \line1[13]_net_1\, Y => 
        \data_out_8_am[13]_net_1\);
    
    \line3_5[16]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(16), C => \line3[16]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[16]_net_1\);
    
    \line4[60]\ : SLE
      port map(D => \line4_5[60]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[60]_net_1\);
    
    \line0[45]\ : SLE
      port map(D => \line0_6[45]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[45]_net_1\);
    
    \data_out_9_0_RNO[0]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_5_i_m2_1_1[0]\, C => \line4[32]_net_1\, D => 
        \line4[0]_net_1\, Y => N_1456);
    
    \data_out_8_bm[12]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[12]_net_1\, C => \line4[44]_net_1\, D
         => \line4[12]_net_1\, Y => \data_out_8_bm[12]_net_1\);
    
    \line2_5[60]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(28), C => \line2[60]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[60]_net_1\);
    
    \data_out_9_0_RNO[31]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_3_rep2\, B => 
        \data_out_9_m2_0_1_1[31]\, C => \line4[63]_net_1\, D => 
        \line4[31]_net_1\, Y => N_56);
    
    \line1[50]\ : SLE
      port map(D => \line1_5[50]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[50]_net_1\);
    
    \line3[30]\ : SLE
      port map(D => \line3_5[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[30]_net_1\);
    
    \line3_5[49]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(17), C => \line3[49]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[49]_net_1\);
    
    \line1[27]\ : SLE
      port map(D => \line1_5[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[27]_net_1\);
    
    \data_out_6_ns[3]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[3]_net_1\, C => \data_out_6_am[3]_net_1\, 
        Y => N_1257);
    
    \line0[50]\ : SLE
      port map(D => \line0_6[50]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[50]_net_1\);
    
    \line0[19]\ : SLE
      port map(D => \line0_6[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[19]_net_1\);
    
    \line2_5[62]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(30), C => \line2[62]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[62]_net_1\);
    
    \line3[56]\ : SLE
      port map(D => \line3_5[56]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[56]_net_1\);
    
    \line1[62]\ : SLE
      port map(D => \line1_5[62]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[62]_net_1\);
    
    \line4_5[16]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(16), 
        C => \line4[16]_net_1\, D => N_47_i, Y => 
        \line4_5[16]_net_1\);
    
    \line4[4]\ : SLE
      port map(D => \line4_5[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[4]_net_1\);
    
    \raddr_pos[3]\ : SLE
      port map(D => raddr_in_net_0(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_1424_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos[3]_net_1\);
    
    \data_out_6_ns[30]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[30]_net_1\, C => \data_out_6_am[30]_net_1\, 
        Y => N_1284);
    
    \data_out_6_bm[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[38]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[38]_net_1\, Y => \data_out_6_bm[6]_net_1\);
    
    \data_out_8_bm_1_1[21]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[53]_net_1\, B => \line0[21]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[21]_net_1\);
    
    \line4[23]\ : SLE
      port map(D => \line4_5[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[23]_net_1\);
    
    \data_out_9_m2_1_bm[31]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[63]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[63]_net_1\, Y => 
        \data_out_9_m2_1_bm[31]_net_1\);
    
    \data_out_6_ns[8]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[8]_net_1\, C => \data_out_6_am[8]_net_1\, 
        Y => N_1262);
    
    \line3[54]\ : SLE
      port map(D => \line3_5[54]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[54]_net_1\);
    
    \data_out_6_ns[28]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[28]_net_1\, C => \data_out_6_am[28]_net_1\, 
        Y => N_1282);
    
    \data_out_6_ns[26]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[26]_net_1\, C => \data_out_6_am[26]_net_1\, 
        Y => N_1280);
    
    \line2_5[54]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(22), C => \line2[54]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[54]_net_1\);
    
    \data_out_8_bm_1_1[10]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[42]_net_1\, B => \line0[10]_net_1\, C
         => \raddr_pos_fast[3]_net_1\, D => \raddr_pos[0]_net_1\, 
        Y => \data_out_8_bm_1_1[10]_net_1\);
    
    \line2_5[23]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(23), C => \line2[23]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[23]_net_1\);
    
    \line0[37]\ : SLE
      port map(D => \line0_6[37]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[37]_net_1\);
    
    \line2_5[0]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(0), C => \line2[0]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[0]_net_1\);
    
    \line1_5[18]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(18), C => \line1[18]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[18]_net_1\);
    
    \data_out_6_bm[22]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[54]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[54]_net_1\, Y => \data_out_6_bm[22]_net_1\);
    
    \line1_5[38]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(6), C => \line1[38]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[38]_net_1\);
    
    \line1[45]\ : SLE
      port map(D => \line1_5[45]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[45]_net_1\);
    
    \line3[51]\ : SLE
      port map(D => \line3_5[51]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[51]_net_1\);
    
    \line1[36]\ : SLE
      port map(D => \line1_5[36]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[36]_net_1\);
    
    \line0_6[30]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(30), C => \line0[30]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[30]_net_1\);
    
    \line2_5[40]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(8), C => \line2[40]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[40]_net_1\);
    
    \line4_5[35]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(3), 
        C => \line4[35]_net_1\, D => N_47_i, Y => 
        \line4_5[35]_net_1\);
    
    \line2[10]\ : SLE
      port map(D => \line2_5[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[10]_net_1\);
    
    \data_out_8_ns[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[5]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[5]_net_1\, Y
         => N_1326);
    
    \line3_5[58]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(26), C => \line3[58]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[58]_net_1\);
    
    \line0_6[32]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(0), C => \line0[32]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[32]_net_1\);
    
    \line2_5[42]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(10), C => \line2[42]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[42]_net_1\);
    
    \line0_6[48]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(16), C => \line0[48]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[48]_net_1\);
    
    un1_wen_18_or_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(2), Y
         => N_44);
    
    \line3[45]\ : SLE
      port map(D => \line3_5[45]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[45]_net_1\);
    
    \line0_6[53]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(21), C => \line0[53]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[53]_net_1\);
    
    \data_out_8_ns[25]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[25]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[25]_net_1\, Y
         => N_1346);
    
    \line1[34]\ : SLE
      port map(D => \line1_5[34]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[34]_net_1\);
    
    \data_out_8_bm_1_1[6]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[38]_net_1\, B => \line0[6]_net_1\, C
         => \raddr_pos_3_rep2\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[6]_net_1\);
    
    \line1_5[8]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(8), C => \line1[8]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[8]_net_1\);
    
    \line1_5[48]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(16), C => \line1[48]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[48]_net_1\);
    
    \line0_6[60]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(28), C => \line0[60]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[60]_net_1\);
    
    \line3[19]\ : SLE
      port map(D => \line3_5[19]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[19]_net_1\);
    
    \data_out_9_0_RNO_0[1]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[33]_net_1\, B => \line0[1]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_5_i_m2_1_1[1]\);
    
    \data_out_6_ns[20]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[20]_net_1\, C => \data_out_6_am[20]_net_1\, 
        Y => N_1274);
    
    \data_out_4_i_m2[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[0]_net_1\, B => \raddr_pos[0]_net_1\, 
        C => \line2[32]_net_1\, Y => N_1458);
    
    \line4[28]\ : SLE
      port map(D => \line4_5[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[28]_net_1\);
    
    \line1[31]\ : SLE
      port map(D => N_28_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => un1_wen_20_or, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[31]_net_1\);
    
    \line0_6[62]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(30), C => \line0[62]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[62]_net_1\);
    
    \data_out_8_bm_1_1[17]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[49]_net_1\, B => \line0[17]_net_1\, C
         => \raddr_pos_3_rep2\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[17]_net_1\);
    
    \line4[10]\ : SLE
      port map(D => \line4_5[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[10]_net_1\);
    
    \line2[56]\ : SLE
      port map(D => \line2_5[56]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[56]_net_1\);
    
    \line4_5[48]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(16), 
        C => \line4[48]_net_1\, D => N_47_i, Y => 
        \line4_5[48]_net_1\);
    
    \line4[3]\ : SLE
      port map(D => \line4_5[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[3]_net_1\);
    
    \line2_5[19]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(19), C => \line2[19]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[19]_net_1\);
    
    \data_out_8_am[18]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[50]_net_1\, D => \line1[18]_net_1\, Y => 
        \data_out_8_am[18]_net_1\);
    
    \line3_5[23]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(23), C => \line3[23]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[23]_net_1\);
    
    \line0[26]\ : SLE
      port map(D => \line0_6[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[26]_net_1\);
    
    \line1[15]\ : SLE
      port map(D => \line1_5[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[15]_net_1\);
    
    \data_out_6_bm[11]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[43]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[43]_net_1\, Y => \data_out_6_bm[11]_net_1\);
    
    \line1[63]\ : SLE
      port map(D => N_26_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => un1_wen_20_or, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[63]_net_1\);
    
    \line0_6[5]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(5), C => \line0[5]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[5]_net_1\);
    
    \line2[54]\ : SLE
      port map(D => \line2_5[54]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[54]_net_1\);
    
    \line2[26]\ : SLE
      port map(D => \line2_5[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[26]_net_1\);
    
    \data_out_6_ns[25]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[25]_net_1\, C => \data_out_6_am[25]_net_1\, 
        Y => N_1279);
    
    \line4[47]\ : SLE
      port map(D => \line4_5[47]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[47]_net_1\);
    
    \data_out_6_bm[20]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[52]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[52]_net_1\, Y => \data_out_6_bm[20]_net_1\);
    
    \data_out_6_am[9]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[9]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[9]_net_1\, Y => \data_out_6_am[9]_net_1\);
    
    \line4_5[30]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(30), 
        C => \line4[30]_net_1\, D => N_47_i, Y => 
        \line4_5[30]_net_1\);
    
    \line0[24]\ : SLE
      port map(D => \line0_6[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[24]_net_1\);
    
    \line2[51]\ : SLE
      port map(D => \line2_5[51]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[51]_net_1\);
    
    \data_out_8_ns[16]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[16]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[16]_net_1\, Y
         => N_1337);
    
    \line0_RNO[31]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(31), C => \line0[31]_net_1\, 
        D => waddr_in_net_0(0), Y => N_32_i_0);
    
    \line4[37]\ : SLE
      port map(D => \line4_5[37]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[37]_net_1\);
    
    \line2[37]\ : SLE
      port map(D => \line2_5[37]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[37]_net_1\);
    
    \data_out_8_bm_1_1[13]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[45]_net_1\, B => \line0[13]_net_1\, C
         => \raddr_pos_fast[3]_net_1\, D => \raddr_pos[0]_net_1\, 
        Y => \data_out_8_bm_1_1[13]_net_1\);
    
    \line4[56]\ : SLE
      port map(D => \line4_5[56]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[56]_net_1\);
    
    \line2[24]\ : SLE
      port map(D => \line2_5[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[24]_net_1\);
    
    \line0[21]\ : SLE
      port map(D => \line0_6[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[21]_net_1\);
    
    \line0_6[37]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(5), C => \line0[37]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[37]_net_1\);
    
    \line2_5[47]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(15), C => \line2[47]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[47]_net_1\);
    
    \line2_5[28]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(28), C => \line2[28]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[28]_net_1\);
    
    \data_out_8_ns[22]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[22]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[22]_net_1\, Y
         => N_1343);
    
    \line2[21]\ : SLE
      port map(D => \line2_5[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[21]_net_1\);
    
    \line0[17]\ : SLE
      port map(D => \line0_6[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[17]_net_1\);
    
    \line1_5[15]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(15), C => \line1[15]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[15]_net_1\);
    
    \line1_5[35]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(3), C => \line1[35]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[35]_net_1\);
    
    \line1[55]\ : SLE
      port map(D => \line1_5[55]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[55]_net_1\);
    
    \line3_5[14]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(14), C => \line3[14]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[14]_net_1\);
    
    \line3[35]\ : SLE
      port map(D => \line3_5[35]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[35]_net_1\);
    
    \line4[54]\ : SLE
      port map(D => \line4_5[54]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[54]_net_1\);
    
    \line0[55]\ : SLE
      port map(D => \line0_6[55]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[55]_net_1\);
    
    \line3_5[55]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(23), C => \line3[55]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[55]_net_1\);
    
    \line4_5[4]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(4), 
        C => \line4[4]_net_1\, D => N_47_i, Y => 
        \line4_5[4]_net_1\);
    
    \line0_6[45]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(13), C => \line0[45]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[45]_net_1\);
    
    \data_out_9_0_RNO_0[29]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => \line4[61]_net_1\, B => \line4[29]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_9_m2_1_1_1[29]\);
    
    \data_out_8_am[22]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[54]_net_1\, D => \line1[22]_net_1\, Y => 
        \data_out_8_am[22]_net_1\);
    
    \line4_5[14]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(14), 
        C => \line4[14]_net_1\, D => N_47_i, Y => 
        \line4_5[14]_net_1\);
    
    \line0_6[58]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(26), C => \line0[58]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[58]_net_1\);
    
    \line4[51]\ : SLE
      port map(D => \line4_5[51]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[51]_net_1\);
    
    \line0_6[36]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(4), C => \line0[36]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[36]_net_1\);
    
    \line2_5[46]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(14), C => \line2[46]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[46]_net_1\);
    
    \data_out_8_am[6]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[38]_net_1\, D => \line1[6]_net_1\, Y => 
        \data_out_8_am[6]_net_1\);
    
    \line1_5[45]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(13), C => \line1[45]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[45]_net_1\);
    
    \data_out_6_i_m2_bm[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[32]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[32]_net_1\, Y => 
        \data_out_6_i_m2_bm[0]_net_1\);
    
    \line0_6[6]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(6), C => \line0[6]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[6]_net_1\);
    
    \line4_5[51]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(19), 
        C => \line4[51]_net_1\, D => N_47_i, Y => 
        \line4_5[51]_net_1\);
    
    \data_out_8_bm_1_1[4]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[36]_net_1\, B => \line0[4]_net_1\, C
         => \raddr_pos_3_rep2\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[4]_net_1\);
    
    \data_out_8_am[23]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[55]_net_1\, D => \line1[23]_net_1\, Y => 
        \data_out_8_am[23]_net_1\);
    
    \raddr_pos[0]\ : SLE
      port map(D => raddr_in_net_0(0), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_1424_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos[0]_net_1\);
    
    \data_out_8_bm[22]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[22]_net_1\, C => \line4[54]_net_1\, D
         => \line4[22]_net_1\, Y => \data_out_8_bm[22]_net_1\);
    
    \line3[59]\ : SLE
      port map(D => \line3_5[59]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[59]_net_1\);
    
    \line4_5[45]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(13), 
        C => \line4[45]_net_1\, D => N_47_i, Y => 
        \line4_5[45]_net_1\);
    
    \line2[15]\ : SLE
      port map(D => \line2_5[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[15]_net_1\);
    
    \data_out_6_ns[2]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[2]_net_1\, C => \data_out_6_am[2]_net_1\, 
        Y => N_1256);
    
    \line3_5[41]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(9), C => \line3[41]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[41]_net_1\);
    
    \line3_5[28]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(28), C => \line3[28]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[28]_net_1\);
    
    \line0_6[19]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(19), C => \line0[19]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[19]_net_1\);
    
    \line2[42]\ : SLE
      port map(D => \line2_5[42]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[42]_net_1\);
    
    \data_out_8_bm[13]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_3_rep2\, B => 
        \data_out_8_bm_1_1[13]_net_1\, C => \line4[45]_net_1\, D
         => \line4[13]_net_1\, Y => \data_out_8_bm[13]_net_1\);
    
    \data_out_8_bm_1_1[5]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[37]_net_1\, B => \line0[5]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[5]_net_1\);
    
    \line4_5[37]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(5), 
        C => \line4[37]_net_1\, D => N_47_i, Y => 
        \line4_5[37]_net_1\);
    
    \line3_5[1]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(1), C => \line3[1]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[1]_net_1\);
    
    \line3[22]\ : SLE
      port map(D => \line3_5[22]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[22]_net_1\);
    
    \line3[17]\ : SLE
      port map(D => \line3_5[17]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[17]_net_1\);
    
    \line1_5[10]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(10), C => \line1[10]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[10]_net_1\);
    
    \line0[42]\ : SLE
      port map(D => \line0_6[42]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[42]_net_1\);
    
    \line1_5[30]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(30), C => \line1[30]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[30]_net_1\);
    
    \line0_6[0]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(0), C => \line0[0]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[0]_net_1\);
    
    \data_out_9_a4_1_1_RNIIPHT[31]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => \raddr_pos[2]_net_1\, B => 
        \raddr_pos[1]_net_1\, C => \raddr_pos[0]_net_1\, D => 
        N_1423_1, Y => \data_out_sn_N_12_mux\);
    
    \data_out_6_bm[30]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[62]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[62]_net_1\, Y => \data_out_6_bm[30]_net_1\);
    
    \line4_5[7]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(7), 
        C => \line4[7]_net_1\, D => N_47_i, Y => 
        \line4_5[7]_net_1\);
    
    \line3_5[4]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(4), C => \line3[4]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[4]_net_1\);
    
    \line2[5]\ : SLE
      port map(D => \line2_5[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[5]_net_1\);
    
    \line1_5[12]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(12), C => \line1[12]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[12]_net_1\);
    
    \line1_5[32]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(0), C => \line1[32]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[32]_net_1\);
    
    \line1[39]\ : SLE
      port map(D => \line1_5[39]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[39]_net_1\);
    
    \data_out_6_i_m2_am[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[1]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[1]_net_1\, Y => \data_out_6_i_m2_am[1]_net_1\);
    
    \line3_5[50]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(18), C => \line3[50]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[50]_net_1\);
    
    \line4[26]\ : SLE
      port map(D => \line4_5[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[26]_net_1\);
    
    \line4[15]\ : SLE
      port map(D => \line4_5[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[15]_net_1\);
    
    \line1_5[5]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(5), C => \line1[5]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[5]_net_1\);
    
    \data_out_6_bm[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[37]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[37]_net_1\, Y => \data_out_6_bm[5]_net_1\);
    
    \line0_6[40]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(8), C => \line0[40]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[40]_net_1\);
    
    un30_wen_0_x2 : CFG3
      generic map(INIT => x"1E")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(2), C
         => waddr_in_net_0(3), Y => N_47_i);
    
    \line3_5[52]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(20), C => \line3[52]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[52]_net_1\);
    
    \data_out_8_bm[14]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[14]_net_1\, C => \line4[46]_net_1\, D
         => \line4[14]_net_1\, Y => \data_out_8_bm[14]_net_1\);
    
    \line2[62]\ : SLE
      port map(D => \line2_5[62]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[62]_net_1\);
    
    \data_out_9_0_RNO[1]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_5_i_m2_1_1[1]\, C => \line4[33]_net_1\, D => 
        \line4[1]_net_1\, Y => N_1455);
    
    \line0_6[42]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(10), C => \line0[42]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[42]_net_1\);
    
    \line2_5[25]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(25), C => \line2[25]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[25]_net_1\);
    
    \line4_5[36]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(4), 
        C => \line4[36]_net_1\, D => N_47_i, Y => 
        \line4_5[36]_net_1\);
    
    ren_pos_RNI0NOS : CFG3
      generic map(INIT => x"02")

      port map(A => \ren_pos\, B => \raddr_pos[2]_net_1\, C => 
        \raddr_pos[1]_net_1\, Y => data_out_sn_N_11_mux);
    
    \line1_5[40]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(8), C => \line1[40]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[40]_net_1\);
    
    \line1[1]\ : SLE
      port map(D => \line1_5[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[1]_net_1\);
    
    \line4[24]\ : SLE
      port map(D => \line4_5[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[24]_net_1\);
    
    \line0_6[9]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(9), C => \line0[9]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[9]_net_1\);
    
    \data_out_9_m2_0_bm[29]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[61]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[61]_net_1\, Y => 
        \data_out_9_m2_0_bm[29]_net_1\);
    
    \data_out_9_0[29]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_1467, B => data_out_sn_N_11_mux, C => 
        \data_out_sn_N_12_mux\, D => N_1468, Y => data_out_9_0_29);
    
    \line1_5[42]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(10), C => \line1[42]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[42]_net_1\);
    
    \line3_5[39]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(7), C => \line3[39]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[39]_net_1\);
    
    \data_out_6_ns[4]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[4]_net_1\, C => \data_out_6_am[4]_net_1\, 
        Y => N_1258);
    
    \line1[20]\ : SLE
      port map(D => \line1_5[20]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[20]_net_1\);
    
    \line4_5[40]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(8), 
        C => \line4[40]_net_1\, D => N_47_i, Y => 
        \line4_5[40]_net_1\);
    
    \line1[42]\ : SLE
      port map(D => \line1_5[42]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[42]_net_1\);
    
    \line4[21]\ : SLE
      port map(D => \line4_5[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[21]_net_1\);
    
    \line1_5[9]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(9), C => \line1[9]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[9]_net_1\);
    
    \line2[59]\ : SLE
      port map(D => \line2_5[59]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[59]_net_1\);
    
    \line0_6[55]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(23), C => \line0[55]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[55]_net_1\);
    
    \line4_5[42]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(10), 
        C => \line4[42]_net_1\, D => N_47_i, Y => 
        \line4_5[42]_net_1\);
    
    \line0_6[1]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(1), C => \line0[1]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[1]_net_1\);
    
    \line0[3]\ : SLE
      port map(D => \line0_6[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[3]_net_1\);
    
    \line1_5[59]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(27), C => \line1[59]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[59]_net_1\);
    
    \line0[29]\ : SLE
      port map(D => N_38_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => un1_wen_7_or, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[29]_net_1\);
    
    un1_wen_18_or_0 : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_1434, B => waddr_in_net_0(3), C => N_44, D
         => \un1_wen_18_or_0_0\, Y => un1_wen_18_or);
    
    \data_out_8_ns[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[6]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[6]_net_1\, Y
         => N_1327);
    
    \line3[42]\ : SLE
      port map(D => \line3_5[42]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[42]_net_1\);
    
    \line2_5[11]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(11), C => \line2[11]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[11]_net_1\);
    
    \line4_5[53]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(21), 
        C => \line4[53]_net_1\, D => N_47_i, Y => 
        \line4_5[53]_net_1\);
    
    \data_out_8_ns[13]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[13]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[13]_net_1\, Y
         => N_1334);
    
    \line3_5[6]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(6), C => \line3[6]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[6]_net_1\);
    
    \data_out_8_am[28]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[60]_net_1\, D => \line1[28]_net_1\, Y => 
        \data_out_8_am[28]_net_1\);
    
    \line2[43]\ : SLE
      port map(D => \line2_5[43]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[43]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line2[29]\ : SLE
      port map(D => N_1442_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[29]_net_1\);
    
    \data_out_6_bm[21]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[53]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[53]_net_1\, Y => \data_out_6_bm[21]_net_1\);
    
    \line4_5_1[32]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(0), 
        C => \line4[32]_net_1\, D => N_46, Y => \line4_5[32]\);
    
    \line0[30]\ : SLE
      port map(D => \line0_6[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[30]_net_1\);
    
    \line3_5[25]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(25), C => \line3[25]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[25]_net_1\);
    
    \line3[23]\ : SLE
      port map(D => \line3_5[23]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[23]_net_1\);
    
    \line3_5[43]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(11), C => \line3[43]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[43]_net_1\);
    
    \line2_5[39]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(7), C => \line2[39]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[39]_net_1\);
    
    \line1[5]\ : SLE
      port map(D => \line1_5[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[5]_net_1\);
    
    \line1_5[17]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(17), C => \line1[17]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[17]_net_1\);
    
    \line1_RNO[29]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(29), C => \line1[29]_net_1\, 
        D => waddr_in_net_0(0), Y => N_34_i_0);
    
    \line1_5[37]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(5), C => \line1[37]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[37]_net_1\);
    
    \line4_5[8]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(8), 
        C => \line4[8]_net_1\, D => N_47_i, Y => 
        \line4_5[8]_net_1\);
    
    \line0[9]\ : SLE
      port map(D => \line0_6[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[9]_net_1\);
    
    \line0[4]\ : SLE
      port map(D => \line0_6[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[4]_net_1\);
    
    \line2_5[4]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(4), C => \line2[4]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[4]_net_1\);
    
    \line0[43]\ : SLE
      port map(D => \line0_6[43]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[43]_net_1\);
    
    \data_out_6_am[11]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[11]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[11]_net_1\, Y => \data_out_6_am[11]_net_1\);
    
    \line4[59]\ : SLE
      port map(D => \line4_5[59]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[59]_net_1\);
    
    \line2_5[20]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(20), C => \line2[20]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[20]_net_1\);
    
    \line3_or[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => un1_wen_18_or, B => 
        sha256_system_sb_0_POWER_ON_RESET_N, Y => 
        \line3_or[0]_net_1\);
    
    \line2_RNO[61]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(29), C => \line2[61]_net_1\, 
        D => waddr_in_net_0(0), Y => N_1441_i_0);
    
    \line3_5[57]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(25), C => \line3[57]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[57]_net_1\);
    
    \data_out_8_bm_1_1[14]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[46]_net_1\, B => \line0[14]_net_1\, C
         => \raddr_pos_3_rep2\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[14]_net_1\);
    
    \line3_5[9]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(9), C => \line3[9]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[9]_net_1\);
    
    \line0_6[7]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(7), C => \line0[7]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[7]_net_1\);
    
    \line1[12]\ : SLE
      port map(D => \line1_5[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[12]_net_1\);
    
    \line2_5[22]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(22), C => \line2[22]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[22]_net_1\);
    
    \line0_6[47]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(15), C => \line0[47]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[47]_net_1\);
    
    \raddr_pos[1]\ : SLE
      port map(D => raddr_in_net_0(1), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_1424_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos[1]_net_1\);
    
    \line0_6[34]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(2), C => \line0[34]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[34]_net_1\);
    
    \line2_5[44]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(12), C => \line2[44]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[44]_net_1\);
    
    \line3[57]\ : SLE
      port map(D => \line3_5[57]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[57]_net_1\);
    
    \data_out_6_ns[27]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[27]_net_1\, C => \data_out_6_am[27]_net_1\, 
        Y => N_1281);
    
    \line0[5]\ : SLE
      port map(D => \line0_6[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[5]_net_1\);
    
    \data_out_6_bm[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[34]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[34]_net_1\, Y => \data_out_6_bm[2]_net_1\);
    
    \line2[63]\ : SLE
      port map(D => N_22_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => un1_wen_19_or, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[63]_net_1\);
    
    \data_out_8_bm_1_1[22]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[54]_net_1\, B => \line0[22]_net_1\, C
         => \raddr_pos_3_rep2\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[22]_net_1\);
    
    \line0_6[21]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(21), C => \line0[21]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[21]_net_1\);
    
    \line0[2]\ : SLE
      port map(D => \line0_6[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[2]_net_1\);
    
    \data_out_8_am[17]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[49]_net_1\, D => \line1[17]_net_1\, Y => 
        \data_out_8_am[17]_net_1\);
    
    \line4_5[5]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(5), 
        C => \line4[5]_net_1\, D => N_47_i, Y => 
        \line4_5[5]_net_1\);
    
    \line1_5[47]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(15), C => \line1[47]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[47]_net_1\);
    
    \data_out_8_ns[21]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[21]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[21]_net_1\, Y
         => N_1342);
    
    \line0_6[50]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(18), C => \line0[50]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[50]_net_1\);
    
    \data_out_6_bm[16]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[48]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[48]_net_1\, Y => \data_out_6_bm[16]_net_1\);
    
    \line0_6[8]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(8), C => \line0[8]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[8]_net_1\);
    
    \data_out_8_bm[6]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[6]_net_1\, C => \line4[38]_net_1\, D
         => \line4[6]_net_1\, Y => \data_out_8_bm[6]_net_1\);
    
    \line1_RNO[63]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(31), C => \line1[63]_net_1\, 
        D => waddr_in_net_0(0), Y => N_26_i_0);
    
    \line1_5[16]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(16), C => \line1[16]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[16]_net_1\);
    
    \line1_5[36]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(4), C => \line1[36]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[36]_net_1\);
    
    \line1[61]\ : SLE
      port map(D => N_1443_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[61]_net_1\);
    
    \line2[48]\ : SLE
      port map(D => \line2_5[48]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[48]_net_1\);
    
    \line0_6[52]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(20), C => \line0[52]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[52]_net_1\);
    
    \line4_5[47]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(15), 
        C => \line4[47]_net_1\, D => N_47_i, Y => 
        \line4_5[47]_net_1\);
    
    \line3_5[56]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(24), C => \line3[56]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[56]_net_1\);
    
    \line3[62]\ : SLE
      port map(D => \line3_5[62]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[62]_net_1\);
    
    \line3[28]\ : SLE
      port map(D => \line3_5[28]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[28]_net_1\);
    
    \line1[43]\ : SLE
      port map(D => \line1_5[43]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[43]_net_1\);
    
    \line0_6[46]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(14), C => \line0[46]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[46]_net_1\);
    
    \data_out_6_ns[5]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[5]_net_1\, C => \data_out_6_am[5]_net_1\, 
        Y => N_1259);
    
    un1_wen_19_or_0 : CFG3
      generic map(INIT => x"D5")

      port map(A => sha256_system_sb_0_POWER_ON_RESET_N, B => 
        N_1434, C => N_61, Y => un1_wen_19_or);
    
    \line2_5[3]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(3), C => \line2[3]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[3]_net_1\);
    
    \data_out_6_bm[13]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[45]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[45]_net_1\, Y => \data_out_6_bm[13]_net_1\);
    
    \data_out_8_bm_1_1[8]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[40]_net_1\, B => \line0[8]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[8]_net_1\);
    
    \line4[62]\ : SLE
      port map(D => \line4_5[62]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[62]_net_1\);
    
    \line1[37]\ : SLE
      port map(D => \line1_5[37]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[37]_net_1\);
    
    \line0[48]\ : SLE
      port map(D => \line0_6[48]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[48]_net_1\);
    
    \line1[52]\ : SLE
      port map(D => \line1_5[52]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[52]_net_1\);
    
    \line4[40]\ : SLE
      port map(D => \line4_5[40]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[40]_net_1\);
    
    \line3_5[20]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(20), C => \line3[20]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[20]_net_1\);
    
    \line3[32]\ : SLE
      port map(D => \line3_5[32]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[32]_net_1\);
    
    \line1_5[46]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(14), C => \line1[46]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[46]_net_1\);
    
    \line0[52]\ : SLE
      port map(D => \line0_6[52]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[52]_net_1\);
    
    \data_out_6_ns[18]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[18]_net_1\, C => \data_out_6_am[18]_net_1\, 
        Y => N_1272);
    
    \data_out_6_ns[16]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[16]_net_1\, C => \data_out_6_am[16]_net_1\, 
        Y => N_1270);
    
    \line3[43]\ : SLE
      port map(D => \line3_5[43]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[43]_net_1\);
    
    \line3_5[22]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(22), C => \line3[22]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[22]_net_1\);
    
    \data_out_6_i_m2_ns[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_i_m2_bm[0]_net_1\, C => 
        \data_out_6_i_m2_am[0]_net_1\, Y => N_1454);
    
    \line4_5[58]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(26), 
        C => \line4[58]_net_1\, D => N_47_i, Y => 
        \line4_5[58]_net_1\);
    
    \line4[30]\ : SLE
      port map(D => \line4_5[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[30]_net_1\);
    
    \line1_5[21]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(21), C => \line1[21]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[21]_net_1\);
    
    \line2[30]\ : SLE
      port map(D => \line2_5[30]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[30]_net_1\);
    
    \line0_6[11]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(11), C => \line0[11]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[11]_net_1\);
    
    \data_out_8_am[5]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[37]_net_1\, D => \line1[5]_net_1\, Y => 
        \data_out_8_am[5]_net_1\);
    
    \line1[6]\ : SLE
      port map(D => \line1_5[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[6]_net_1\);
    
    \line4_5[46]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(14), 
        C => \line4[46]_net_1\, D => N_47_i, Y => 
        \line4_5[46]_net_1\);
    
    \line1_5[3]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(3), C => \line1[3]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[3]_net_1\);
    
    \line2_5[13]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(13), C => \line2[13]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[13]_net_1\);
    
    \data_out_8_bm[23]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_3_rep2\, B => 
        \data_out_8_bm_1_1[23]_net_1\, C => \line4[55]_net_1\, D
         => \line4[23]_net_1\, Y => \data_out_8_bm[23]_net_1\);
    
    \line4_5[34]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(2), 
        C => \line4[34]_net_1\, D => N_47_i, Y => 
        \line4_5[34]_net_1\);
    
    \line4_5[21]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(21), 
        C => \line4[21]_net_1\, D => N_47_i, Y => 
        \line4_5[21]_net_1\);
    
    \line0[10]\ : SLE
      port map(D => \line0_6[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[10]_net_1\);
    
    \line3_5[48]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(16), C => \line3[48]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[48]_net_1\);
    
    \line4[5]\ : SLE
      port map(D => \line4_5[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[5]_net_1\);
    
    \line2_5[27]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(27), C => \line2[27]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[27]_net_1\);
    
    \line1_5[2]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(2), C => \line1[2]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[2]_net_1\);
    
    \line2[57]\ : SLE
      port map(D => \line2_5[57]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[57]_net_1\);
    
    \line2[0]\ : SLE
      port map(D => \line2_5[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[0]_net_1\);
    
    \data_out_8_ns[28]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[28]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[28]_net_1\, Y
         => N_1349);
    
    \data_out_8_ns[15]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[15]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[15]_net_1\, Y
         => N_1336);
    
    un5_wen_0_a2 : CFG3
      generic map(INIT => x"02")

      port map(A => waddr_in_net_0(3), B => N_44, C => 
        waddr_in_net_0(0), Y => un5_wen);
    
    \line1[25]\ : SLE
      port map(D => \line1_5[25]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[25]_net_1\);
    
    \line4[2]\ : SLE
      port map(D => \line4_5[2]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[2]_net_1\);
    
    \line4[29]\ : SLE
      port map(D => N_1438_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[29]_net_1\);
    
    \line1[48]\ : SLE
      port map(D => \line1_5[48]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[48]_net_1\);
    
    \line1[13]\ : SLE
      port map(D => \line1_5[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[13]_net_1\);
    
    \line2[12]\ : SLE
      port map(D => \line2_5[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[12]_net_1\);
    
    \line0[27]\ : SLE
      port map(D => \line0_6[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[27]_net_1\);
    
    \data_out_6_ns[10]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[10]_net_1\, C => \data_out_6_am[10]_net_1\, 
        Y => N_1264);
    
    \line4_5[6]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(6), 
        C => \line4[6]_net_1\, D => N_47_i, Y => 
        \line4_5[6]_net_1\);
    
    \data_out_6_i_m2_am[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[0]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[0]_net_1\, Y => \data_out_6_i_m2_am[0]_net_1\);
    
    \line2[27]\ : SLE
      port map(D => \line2_5[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[27]_net_1\);
    
    \line2_5[59]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(27), C => \line2[59]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[59]_net_1\);
    
    \line0_6[57]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(25), C => \line0[57]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[57]_net_1\);
    
    \data_out_8_bm[24]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[24]_net_1\, C => \line4[56]_net_1\, D
         => \line4[24]_net_1\, Y => \data_out_8_bm[24]_net_1\);
    
    \line3[48]\ : SLE
      port map(D => \line3_5[48]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[48]_net_1\);
    
    \line2_5[7]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(7), C => \line2[7]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[7]_net_1\);
    
    \line2_5[26]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(26), C => \line2[26]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[26]_net_1\);
    
    \line0_6[23]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(23), C => \line0[23]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[23]_net_1\);
    
    un1_wen_20_or_0_m2 : CFG3
      generic map(INIT => x"CA")

      port map(A => waddr_in_net_0(1), B => waddr_in_net_0(3), C
         => waddr_in_net_0(2), Y => N_62);
    
    \line0[35]\ : SLE
      port map(D => \line0_6[35]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[35]_net_1\);
    
    \line3[63]\ : SLE
      port map(D => N_18_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => sha256_system_sb_0_POWER_ON_RESET_N, SD
         => GND_net_1, LAT => GND_net_1, Q => \line3[63]_net_1\);
    
    \data_out_8_bm_1_1[20]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[52]_net_1\, B => \line0[20]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[20]_net_1\);
    
    \line4[57]\ : SLE
      port map(D => \line4_5[57]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[57]_net_1\);
    
    raddr_pos_3_rep1 : SLE
      port map(D => raddr_in_net_0(3), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_1424_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_3_rep1\);
    
    \data_out_8_bm_1_1[16]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[48]_net_1\, B => \line0[16]_net_1\, C
         => \raddr_pos_3_rep2\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[16]_net_1\);
    
    \line4[12]\ : SLE
      port map(D => \line4_5[12]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[12]_net_1\);
    
    \data_out_6_ns[15]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[15]_net_1\, C => \data_out_6_am[15]_net_1\, 
        Y => N_1269);
    
    \line4[63]\ : SLE
      port map(D => \line4_5[63]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[63]_net_1\);
    
    \data_out_8_bm[15]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_3_rep2\, B => 
        \data_out_8_bm_1_1[15]_net_1\, C => \line4[47]_net_1\, D
         => \line4[15]_net_1\, Y => \data_out_8_bm[15]_net_1\);
    
    ren_pos_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => AHB_slave_dummy_0_read_en, B => 
        sha256_system_sb_0_POWER_ON_RESET_N, Y => N_35_i_0);
    
    \line3_5[27]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(27), C => \line3[27]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[27]_net_1\);
    
    \line1[53]\ : SLE
      port map(D => \line1_5[53]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[53]_net_1\);
    
    \data_out_6_ns[22]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[22]_net_1\, C => \data_out_6_am[22]_net_1\, 
        Y => N_1276);
    
    \line3[33]\ : SLE
      port map(D => \line3_5[33]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[33]_net_1\);
    
    \line0_6[56]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(24), C => \line0[56]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[56]_net_1\);
    
    \line1_5[51]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(19), C => \line1[51]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[51]_net_1\);
    
    \line3[10]\ : SLE
      port map(D => \line3_5[10]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[10]_net_1\);
    
    \line4_5_1[31]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(31), 
        C => \line4[31]_net_1\, D => N_46, Y => \line4_5[31]\);
    
    \line0[53]\ : SLE
      port map(D => \line0_6[53]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[53]_net_1\);
    
    \line1[18]\ : SLE
      port map(D => \line1_5[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[18]_net_1\);
    
    \data_out_8_ns[12]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[12]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[12]_net_1\, Y
         => N_1333);
    
    \data_out_6_i_m2_ns[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_i_m2_bm[1]_net_1\, C => 
        \data_out_6_i_m2_am[1]_net_1\, Y => N_1453);
    
    \data_out_8_am[2]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[34]_net_1\, D => \line1[2]_net_1\, Y => 
        \data_out_8_am[2]_net_1\);
    
    \line1[3]\ : SLE
      port map(D => \line1_5[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[3]_net_1\);
    
    \line4_5[55]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(23), 
        C => \line4[55]_net_1\, D => N_47_i, Y => 
        \line4_5[55]_net_1\);
    
    \line2_5[18]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(18), C => \line2[18]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[18]_net_1\);
    
    \data_out_8_bm_1_1[27]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[59]_net_1\, B => \line0[27]_net_1\, C
         => \raddr_pos_3_rep1\, D => \raddr_pos[0]_net_1\, Y => 
        \data_out_8_bm_1_1[27]_net_1\);
    
    \line1_5[23]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(23), C => \line1[23]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[23]_net_1\);
    
    \line0_6[13]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(13), C => \line0[13]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[13]_net_1\);
    
    \line3_5[26]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(26), C => \line3[26]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[26]_net_1\);
    
    \line2[46]\ : SLE
      port map(D => \line2_5[46]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[46]_net_1\);
    
    \line1_5[14]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(14), C => \line1[14]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[14]_net_1\);
    
    \line1_5[34]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(2), C => \line1[34]_net_1\, D
         => waddr_in_net_0(0), Y => \line1_5[34]_net_1\);
    
    \raddr_pos[2]\ : SLE
      port map(D => raddr_in_net_0(2), CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_1424_i_0, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos[2]_net_1\);
    
    \line3_RNO[63]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(31), C => \line3[63]_net_1\, 
        D => waddr_in_net_0(0), Y => N_18_i_0);
    
    \data_out_6_am[21]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[21]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[21]_net_1\, Y => \data_out_6_am[21]_net_1\);
    
    \line4_5[23]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(23), 
        C => \line4[23]_net_1\, D => N_47_i, Y => 
        \line4_5[23]_net_1\);
    
    \line3_5[45]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(13), C => \line3[45]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[45]_net_1\);
    
    \line3[3]\ : SLE
      port map(D => \line3_5[3]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[3]_net_1\);
    
    \line3[26]\ : SLE
      port map(D => \line3_5[26]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[26]_net_1\);
    
    \line3_5[54]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(22), C => \line3[54]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[54]_net_1\);
    
    \line2[13]\ : SLE
      port map(D => \line2_5[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[13]_net_1\);
    
    \data_out_6_bm[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[39]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[39]_net_1\, Y => \data_out_6_bm[7]_net_1\);
    
    \line0_6[44]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(12), C => \line0[44]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[44]_net_1\);
    
    \line4[45]\ : SLE
      port map(D => \line4_5[45]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[45]_net_1\);
    
    \line1[58]\ : SLE
      port map(D => \line1_5[58]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[58]_net_1\);
    
    \line0[46]\ : SLE
      port map(D => \line0_6[46]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[46]_net_1\);
    
    \line0[60]\ : SLE
      port map(D => \line0_6[60]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[60]_net_1\);
    
    \line3[38]\ : SLE
      port map(D => \line3_5[38]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[38]_net_1\);
    
    \line2[44]\ : SLE
      port map(D => \line2_5[44]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[44]_net_1\);
    
    \data_out_8_ns[24]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[24]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[24]_net_1\, Y
         => N_1345);
    
    \line0[58]\ : SLE
      port map(D => \line0_6[58]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[58]_net_1\);
    
    \data_out_8_am[27]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \raddr_pos[0]_net_1\, B => N_1423_1, C => 
        \line2[59]_net_1\, D => \line1[27]_net_1\, Y => 
        \data_out_8_am[27]_net_1\);
    
    \line1_5[44]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(12), C => \line1[44]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[44]_net_1\);
    
    \line0[7]\ : SLE
      port map(D => \line0_6[7]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[7]_net_1\);
    
    \line3[24]\ : SLE
      port map(D => \line3_5[24]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[24]_net_1\);
    
    \line4[35]\ : SLE
      port map(D => \line4_5[35]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[35]_net_1\);
    
    \data_out_8_ns[9]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \data_out_8_bm[9]_net_1\, B => 
        data_out_sn_N_11_mux, C => \data_out_8_am[9]_net_1\, Y
         => N_1330);
    
    \line2[41]\ : SLE
      port map(D => \line2_5[41]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[41]_net_1\);
    
    \line2[35]\ : SLE
      port map(D => \line2_5[35]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[35]_net_1\);
    
    \data_out_6_bm[26]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[58]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[58]_net_1\, Y => \data_out_6_bm[26]_net_1\);
    
    \data_out_6_am[14]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[14]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[14]_net_1\, Y => \data_out_6_am[14]_net_1\);
    
    \line0_6[28]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(28), C => \line0[28]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[28]_net_1\);
    
    \line3_5[19]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(19), C => \line3[19]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[19]_net_1\);
    
    \line0[44]\ : SLE
      port map(D => \line0_6[44]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[44]_net_1\);
    
    \data_out_8_bm_1_1[23]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line0[55]_net_1\, B => \line0[23]_net_1\, C
         => \raddr_pos_fast[3]_net_1\, D => \raddr_pos[0]_net_1\, 
        Y => \data_out_8_bm_1_1[23]_net_1\);
    
    \line3[21]\ : SLE
      port map(D => \line3_5[21]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[21]_net_1\);
    
    \line4_5[44]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(12), 
        C => \line4[44]_net_1\, D => N_47_i, Y => 
        \line4_5[44]_net_1\);
    
    \line4[13]\ : SLE
      port map(D => \line4_5[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[13]_net_1\);
    
    \line0_RNO[63]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(31), C => \line0[63]_net_1\, 
        D => waddr_in_net_0(0), Y => N_30_i_0);
    
    \line0[15]\ : SLE
      port map(D => \line0_6[15]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[15]_net_1\);
    
    \data_out_6_bm[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[35]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[35]_net_1\, Y => \data_out_6_bm[3]_net_1\);
    
    \line4[27]\ : SLE
      port map(D => \line4_5[27]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[27]_net_1\);
    
    \line0[41]\ : SLE
      port map(D => \line0_6[41]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[41]_net_1\);
    
    \data_out_8_bm[5]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \data_out_8_bm_1_1[5]_net_1\, C => \line4[37]_net_1\, D
         => \line4[5]_net_1\, Y => \data_out_8_bm[5]_net_1\);
    
    \data_out_6_bm[23]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[55]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[55]_net_1\, Y => \data_out_6_bm[23]_net_1\);
    
    \line3_5[33]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(1), C => \line3[33]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[33]_net_1\);
    
    \line3[6]\ : SLE
      port map(D => \line3_5[6]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[6]_net_1\);
    
    \line4_5[19]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(19), 
        C => \line4[19]_net_1\, D => N_47_i, Y => 
        \line4_5[19]_net_1\);
    
    \data_out_6_bm[14]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[46]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[46]_net_1\, Y => \data_out_6_bm[14]_net_1\);
    
    \data_out_6_am[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[6]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[6]_net_1\, Y => \data_out_6_am[6]_net_1\);
    
    \line4_5[50]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(18), 
        C => \line4[50]_net_1\, D => N_47_i, Y => 
        \line4_5[50]_net_1\);
    
    \line4_5[9]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(9), 
        C => \line4[9]_net_1\, D => N_47_i, Y => 
        \line4_5[9]_net_1\);
    
    un30_wen_0_x2_RNIL99T : CFG3
      generic map(INIT => x"5D")

      port map(A => sha256_system_sb_0_POWER_ON_RESET_N, B => 
        N_1434, C => N_47_i, Y => un1_wen_7_or);
    
    \data_out_8_bm[10]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_3_rep2\, B => 
        \data_out_8_bm_1_1[10]_net_1\, C => \line4[42]_net_1\, D
         => \line4[10]_net_1\, Y => \data_out_8_bm[10]_net_1\);
    
    \line2[18]\ : SLE
      port map(D => \line2_5[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[18]_net_1\);
    
    \line1[46]\ : SLE
      port map(D => \line1_5[46]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[46]_net_1\);
    
    \line0_6[4]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(4), C => \line0[4]_net_1\, D
         => waddr_in_net_0(0), Y => \line0_6[4]_net_1\);
    
    \line4_5[52]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(20), 
        C => \line4[52]_net_1\, D => N_47_i, Y => 
        \line4_5[52]_net_1\);
    
    \data_out_6_bm[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[36]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[36]_net_1\, Y => \data_out_6_bm[4]_net_1\);
    
    \line2_5[8]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(8), C => \line2[8]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[8]_net_1\);
    
    \line1_5[53]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(21), C => \line1[53]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[53]_net_1\);
    
    \line2[61]\ : SLE
      port map(D => N_1441_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[61]_net_1\);
    
    \line3_5[40]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(8), C => \line3[40]_net_1\, D
         => waddr_in_net_0(0), Y => \line3_5[40]_net_1\);
    
    \line2[9]\ : SLE
      port map(D => \line2_5[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_19_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line2[9]_net_1\);
    
    \line0[1]\ : SLE
      port map(D => \line0_6[1]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_7_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line0[1]_net_1\);
    
    \data_out_6_bm[8]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line1[40]_net_1\, B => \raddr_pos[2]_net_1\, 
        C => \line3[40]_net_1\, Y => \data_out_6_bm[8]_net_1\);
    
    \data_out_6_ns[24]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[24]_net_1\, C => \data_out_6_am[24]_net_1\, 
        Y => N_1278);
    
    \line3[50]\ : SLE
      port map(D => \line3_5[50]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[50]_net_1\);
    
    \line3[46]\ : SLE
      port map(D => \line3_5[46]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[46]_net_1\);
    
    \line3_5[42]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(10), C => \line3[42]_net_1\, 
        D => waddr_in_net_0(0), Y => \line3_5[42]_net_1\);
    
    \line1[44]\ : SLE
      port map(D => \line1_5[44]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[44]_net_1\);
    
    \data_out_9_m2_0_am[29]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[29]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[29]_net_1\, Y => 
        \data_out_9_m2_0_am[29]_net_1\);
    
    \line1_5[28]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(28), C => \line1[28]_net_1\, 
        D => waddr_in_net_0(0), Y => \line1_5[28]_net_1\);
    
    \data_out_6_ns[6]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_6_bm[6]_net_1\, C => \data_out_6_am[6]_net_1\, 
        Y => N_1260);
    
    \line0_6[18]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(18), C => \line0[18]_net_1\, 
        D => waddr_in_net_0(0), Y => \line0_6[18]_net_1\);
    
    \line2_5[24]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(24), C => \line2[24]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[24]_net_1\);
    
    \line2_5[15]\ : CFG4
      generic map(INIT => x"5044")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(15), C => \line2[15]_net_1\, 
        D => waddr_in_net_0(0), Y => \line2_5[15]_net_1\);
    
    \line2_5[33]\ : CFG4
      generic map(INIT => x"4450")

      port map(A => waddr_in_net_0(3), B => 
        AHB_slave_dummy_0_mem_wdata(1), C => \line2[33]_net_1\, D
         => waddr_in_net_0(0), Y => \line2_5[33]_net_1\);
    
    \line1[41]\ : SLE
      port map(D => \line1_5[41]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[41]_net_1\);
    
    \line4[18]\ : SLE
      port map(D => \line4_5[18]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_4_or, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line4[18]_net_1\);
    
    \data_out_6_am[15]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[15]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[15]_net_1\, Y => \data_out_6_am[15]_net_1\);
    
    \data_out_6_am[12]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \line2[12]_net_1\, B => \raddr_pos[1]_net_1\, 
        C => \line3[12]_net_1\, Y => \data_out_6_am[12]_net_1\);
    
    \line4_5[28]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un5_wen, B => AHB_slave_dummy_0_mem_wdata(28), 
        C => \line4[28]_net_1\, D => N_47_i, Y => 
        \line4_5[28]_net_1\);
    
    \line3[44]\ : SLE
      port map(D => \line3_5[44]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => \line3_or[0]_net_1\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line3[44]_net_1\);
    
    \line1[4]\ : SLE
      port map(D => \line1_5[4]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => un1_wen_20_or, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        sha256_system_sb_0_POWER_ON_RESET_N, SD => GND_net_1, LAT
         => GND_net_1, Q => \line1[4]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity AHB_slave_dummy is

    port( waddr_in_net_0                                     : out   std_logic_vector(3 downto 0);
          raddr_in_net_0                                     : out   std_logic_vector(3 downto 0);
          arbRegSMCurrentState                               : in    std_logic_vector(15 to 15);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR  : in    std_logic_vector(27 downto 24);
          masterAddrInProg                                   : in    std_logic_vector(3 downto 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS : in    std_logic_vector(1 to 1);
          sha256_system_sb_0_POWER_ON_RESET_N                : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                       : in    std_logic;
          N_42_i_0                                           : in    std_logic;
          N_44_i_0                                           : in    std_logic;
          N_46_i_0                                           : in    std_logic;
          N_48_i_0                                           : in    std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY             : out   std_logic;
          AHB_slave_dummy_0_write_en                         : out   std_logic;
          AHB_slave_dummy_0_read_en                          : out   std_logic;
          N_16_i_0                                           : in    std_logic;
          masterRegAddrSel                                   : in    std_logic;
          regHTRANS                                          : in    std_logic;
          N_359                                              : in    std_logic;
          N_344                                              : in    std_logic;
          N_253                                              : in    std_logic;
          N_321_2                                            : in    std_logic;
          N_354                                              : in    std_logic;
          N_355                                              : in    std_logic;
          N_358                                              : in    std_logic;
          N_211                                              : in    std_logic;
          N_395                                              : in    std_logic;
          N_403                                              : in    std_logic;
          N_401                                              : in    std_logic;
          N_208                                              : in    std_logic;
          regHWRITE                                          : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE : in    std_logic;
          N_36_2                                             : out   std_logic
        );

end AHB_slave_dummy;

architecture DEF_ARCH of AHB_slave_dummy is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \FSM[0]_net_1\, \FSM_i_0[0]\, VCC_net_1, N_292, 
        GND_net_1, N_290, 
        \sha256_system_sb_0_AMBA_SLAVE_0_HREADY\, N_65, N_77_i_0, 
        \hwrite_r\, N_372, \FSM[1]_net_1\, \FSM_ns[1]\, 
        \un1_lsram_waddr_0_sqmuxa_i_0_a1_0\, 
        \lsram_raddr_1_sqmuxa_i_o2_i_a2_2_1_0\, \g0_1\, 
        lsram_raddr_1_sqmuxa_i_o2_i_o2_7, \g0_2_1\, 
        \lsram_waddr_0_sqmuxa_i_i_a2_0_0\, \g0_1_3\, g0_1_2, 
        N_325_0_0_0, g0_1_5, lsram_raddr_1_sqmuxa_i_o2_i_a2_1_0, 
        N_77_i_1, \un1_lsram_waddr_0_sqmuxa_i_0\, 
        \un1_lsram_raddr_1_sqmuxa_i_i_0_1\, 
        \un1_lsram_raddr_1_sqmuxa_i_i_a2\, 
        \un1_lsram_raddr_1_sqmuxa_i_i_a2_RNO\ : std_logic;

begin 

    sha256_system_sb_0_AMBA_SLAVE_0_HREADY <= 
        \sha256_system_sb_0_AMBA_SLAVE_0_HREADY\;

    ready : SLE
      port map(D => \FSM[0]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_65, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sha256_system_sb_0_AMBA_SLAVE_0_HREADY\);
    
    lsram_raddr_1_sqmuxa_i_o2_i_a2_2 : CFG4
      generic map(INIT => x"00C8")

      port map(A => N_359, B => 
        \lsram_raddr_1_sqmuxa_i_o2_i_a2_2_1_0\, C => N_344, D => 
        \g0_1\, Y => N_372);
    
    write_en : SLE
      port map(D => \FSM_i_0[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_77_i_0, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => AHB_slave_dummy_0_write_en);
    
    \lsram_raddr[3]\ : SLE
      port map(D => N_48_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_290, ALn => sha256_system_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => raddr_in_net_0(3));
    
    \lsram_raddr[2]\ : SLE
      port map(D => N_46_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_290, ALn => sha256_system_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => raddr_in_net_0(2));
    
    g0_1 : CFG2
      generic map(INIT => x"1")

      port map(A => masterRegAddrSel, B => 
        arbRegSMCurrentState(15), Y => 
        lsram_raddr_1_sqmuxa_i_o2_i_a2_1_0);
    
    un1_lsram_waddr_0_sqmuxa_i_0 : CFG4
      generic map(INIT => x"FBAA")

      port map(A => \FSM_ns[1]\, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), C
         => masterRegAddrSel, D => 
        \un1_lsram_waddr_0_sqmuxa_i_0_a1_0\, Y => 
        \un1_lsram_waddr_0_sqmuxa_i_0\);
    
    un1_lsram_waddr_0_sqmuxa_i_0_a1_0 : CFG3
      generic map(INIT => x"15")

      port map(A => \FSM[0]_net_1\, B => masterRegAddrSel, C => 
        regHTRANS, Y => \un1_lsram_waddr_0_sqmuxa_i_0_a1_0\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \lsram_raddr[0]\ : SLE
      port map(D => N_42_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_290, ALn => sha256_system_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => raddr_in_net_0(0));
    
    un1_lsram_raddr_1_sqmuxa_i_i_0 : CFG4
      generic map(INIT => x"00DC")

      port map(A => lsram_raddr_1_sqmuxa_i_o2_i_o2_7, B => 
        \FSM_ns[1]\, C => \un1_lsram_raddr_1_sqmuxa_i_i_0_1\, D
         => \un1_lsram_raddr_1_sqmuxa_i_i_a2\, Y => N_65);
    
    \lsram_waddr[0]\ : SLE
      port map(D => N_42_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_292, ALn => sha256_system_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => waddr_in_net_0(0));
    
    \lsram_waddr[3]\ : SLE
      port map(D => N_48_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_292, ALn => sha256_system_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => waddr_in_net_0(3));
    
    \FSM_RNIR3G7[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \FSM[0]_net_1\, Y => \FSM_i_0[0]\);
    
    hwrite_r : SLE
      port map(D => N_16_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_372, ALn => sha256_system_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \hwrite_r\);
    
    \lsram_waddr[2]\ : SLE
      port map(D => N_46_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_292, ALn => sha256_system_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => waddr_in_net_0(2));
    
    \lsram_waddr[1]\ : SLE
      port map(D => N_44_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_292, ALn => sha256_system_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => waddr_in_net_0(1));
    
    \FSM[0]\ : SLE
      port map(D => N_372, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \FSM[0]_net_1\);
    
    un1_lsram_raddr_1_sqmuxa_i_i_0_1 : CFG4
      generic map(INIT => x"3F2A")

      port map(A => N_344, B => N_208, C => 
        lsram_raddr_1_sqmuxa_i_o2_i_a2_1_0, D => N_359, Y => 
        \un1_lsram_raddr_1_sqmuxa_i_i_0_1\);
    
    lsram_raddr_1_sqmuxa_i_o2_i_a2_2_1_0 : CFG2
      generic map(INIT => x"1")

      port map(A => lsram_raddr_1_sqmuxa_i_o2_i_o2_7, B => 
        \FSM[0]_net_1\, Y => 
        \lsram_raddr_1_sqmuxa_i_o2_i_a2_2_1_0\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    g0_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_354, B => N_355, C => N_358, D => N_211, Y
         => N_325_0_0_0);
    
    lsram_waddr_0_sqmuxa_i_i_a2_0_0 : CFG4
      generic map(INIT => x"4450")

      port map(A => \FSM[0]_net_1\, B => regHTRANS, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), D
         => masterRegAddrSel, Y => 
        \lsram_waddr_0_sqmuxa_i_i_a2_0_0\);
    
    un1_lsram_raddr_1_sqmuxa_i_i_a2 : CFG4
      generic map(INIT => x"1F0E")

      port map(A => \FSM[0]_net_1\, B => masterRegAddrSel, C => 
        \un1_lsram_raddr_1_sqmuxa_i_i_a2_RNO\, D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, Y => 
        \un1_lsram_raddr_1_sqmuxa_i_i_a2\);
    
    \lsram_raddr[1]\ : SLE
      port map(D => N_44_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_290, ALn => sha256_system_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => raddr_in_net_0(1));
    
    g0_2_1 : CFG3
      generic map(INIT => x"01")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(24), B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(27), 
        C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(26), Y
         => \g0_2_1\);
    
    lsram_waddr_0_sqmuxa_i_i_a2_0_0_RNILJGV7_0 : CFG4
      generic map(INIT => x"0100")

      port map(A => N_253, B => \g0_1\, C => 
        lsram_raddr_1_sqmuxa_i_o2_i_o2_7, D => 
        \lsram_waddr_0_sqmuxa_i_i_a2_0_0\, Y => N_290);
    
    read_en : SLE
      port map(D => \FSM_i_0[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_65, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => AHB_slave_dummy_0_read_en);
    
    g0_1_3 : CFG3
      generic map(INIT => x"FE")

      port map(A => masterAddrInProg(3), B => masterAddrInProg(2), 
        C => N_321_2, Y => \g0_1_3\);
    
    lsram_raddr_1_sqmuxa_i_o2_i_o2_2 : CFG2
      generic map(INIT => x"E")

      port map(A => N_401, B => N_403, Y => N_36_2);
    
    \FSM_RNI4AE85[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => N_403, B => N_325_0_0_0, C => g0_1_5, D => 
        N_401, Y => lsram_raddr_1_sqmuxa_i_o2_i_o2_7);
    
    write_en_RNO : CFG4
      generic map(INIT => x"D0F0")

      port map(A => lsram_raddr_1_sqmuxa_i_o2_i_a2_1_0, B => 
        \FSM[0]_net_1\, C => N_77_i_1, D => N_208, Y => N_77_i_0);
    
    lsram_waddr_0_sqmuxa_i_i_a2_0_0_RNILJGV7 : CFG4
      generic map(INIT => x"0200")

      port map(A => N_253, B => \g0_1\, C => 
        lsram_raddr_1_sqmuxa_i_o2_i_o2_7, D => 
        \lsram_waddr_0_sqmuxa_i_i_a2_0_0\, Y => N_292);
    
    write_en_RNO_0 : CFG4
      generic map(INIT => x"0B0A")

      port map(A => \FSM[0]_net_1\, B => 
        lsram_raddr_1_sqmuxa_i_o2_i_o2_7, C => 
        \un1_lsram_waddr_0_sqmuxa_i_0\, D => N_253, Y => N_77_i_1);
    
    \FSM[1]\ : SLE
      port map(D => \FSM_ns[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \FSM[1]_net_1\);
    
    \FSM_RNIN40P2[1]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => N_358, B => g0_1_2, C => N_395, D => \g0_1_3\, 
        Y => g0_1_5);
    
    \FSM_RNI5UTQ[1]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \FSM[1]_net_1\, B => masterAddrInProg(1), C
         => \sha256_system_sb_0_AMBA_SLAVE_0_HREADY\, Y => g0_1_2);
    
    g0_2 : CFG4
      generic map(INIT => x"000B")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(25), B
         => \g0_2_1\, C => arbRegSMCurrentState(15), D => 
        masterRegAddrSel, Y => \g0_1\);
    
    un1_lsram_raddr_1_sqmuxa_i_i_a2_RNO : CFG3
      generic map(INIT => x"35")

      port map(A => regHWRITE, B => \hwrite_r\, C => 
        \FSM[0]_net_1\, Y => 
        \un1_lsram_raddr_1_sqmuxa_i_i_a2_RNO\);
    
    un1_lsram_waddr_0_sqmuxa_i_0_a4 : CFG2
      generic map(INIT => x"2")

      port map(A => \FSM[0]_net_1\, B => \hwrite_r\, Y => 
        \FSM_ns[1]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_system_sb_MSS is

    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : inout std_logic_vector(1 to 1) := (others => 'Z');
          arbRegSMCurrentState_ns_i_0_0_0_a0_0                 : out   std_logic_vector(1 to 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : out   std_logic_vector(31 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : in    std_logic_vector(0 to 0);
          data_out_9_0_29                                      : in    std_logic;
          data_out_9_0_31                                      : in    std_logic;
          data_out_9_0_1                                       : in    std_logic;
          data_out_9_0_0                                       : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_26 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_27 : out   std_logic;
          masterRegAddrSel                                     : in    std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic;
          N_1256                                               : in    std_logic;
          data_out_sn_N_12_mux                                 : in    std_logic;
          N_1323                                               : in    std_logic;
          hready_m_xhdl339                                     : in    std_logic;
          N_1257                                               : in    std_logic;
          N_1324                                               : in    std_logic;
          N_1258                                               : in    std_logic;
          N_1325                                               : in    std_logic;
          N_1259                                               : in    std_logic;
          N_1326                                               : in    std_logic;
          N_1260                                               : in    std_logic;
          N_1327                                               : in    std_logic;
          N_1261                                               : in    std_logic;
          N_1328                                               : in    std_logic;
          N_1262                                               : in    std_logic;
          N_1329                                               : in    std_logic;
          N_1263                                               : in    std_logic;
          N_1330                                               : in    std_logic;
          N_1264                                               : in    std_logic;
          N_1331                                               : in    std_logic;
          N_1265                                               : in    std_logic;
          N_1332                                               : in    std_logic;
          N_1266                                               : in    std_logic;
          N_1333                                               : in    std_logic;
          N_1267                                               : in    std_logic;
          N_1334                                               : in    std_logic;
          N_1268                                               : in    std_logic;
          N_1335                                               : in    std_logic;
          N_1269                                               : in    std_logic;
          N_1336                                               : in    std_logic;
          N_1270                                               : in    std_logic;
          N_1337                                               : in    std_logic;
          N_1271                                               : in    std_logic;
          N_1338                                               : in    std_logic;
          N_1272                                               : in    std_logic;
          N_1339                                               : in    std_logic;
          N_1273                                               : in    std_logic;
          N_1340                                               : in    std_logic;
          N_1274                                               : in    std_logic;
          N_1341                                               : in    std_logic;
          N_1275                                               : in    std_logic;
          N_1342                                               : in    std_logic;
          N_1276                                               : in    std_logic;
          N_1343                                               : in    std_logic;
          N_1277                                               : in    std_logic;
          N_1344                                               : in    std_logic;
          N_1278                                               : in    std_logic;
          N_1345                                               : in    std_logic;
          N_1279                                               : in    std_logic;
          N_1346                                               : in    std_logic;
          N_1280                                               : in    std_logic;
          N_1347                                               : in    std_logic;
          N_1281                                               : in    std_logic;
          N_1348                                               : in    std_logic;
          N_1282                                               : in    std_logic;
          N_1349                                               : in    std_logic;
          N_1284                                               : in    std_logic;
          N_1351                                               : in    std_logic;
          N_1446                                               : in    std_logic;
          N_1423_3                                             : in    std_logic;
          N_53                                                 : in    std_logic;
          N_1457                                               : in    std_logic;
          N_1458                                               : in    std_logic;
          GPIO_2_M2F_c                                         : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N      : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : out   std_logic;
          sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F           : out   std_logic;
          GPIO_1_M2F_c                                         : out   std_logic;
          GPIO_0_M2F_c                                         : out   std_logic;
          N_23_i_0                                             : in    std_logic;
          FIC_0_LOCK                                           : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic
        );

end sha256_system_sb_MSS;

architecture DEF_ARCH of sha256_system_sb_MSS is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MSS_060

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MGPIO0B_IN                              : in    std_logic := 'U';
          MGPIO10B_IN                             : in    std_logic := 'U';
          MGPIO1B_IN                              : in    std_logic := 'U';
          MGPIO25A_IN                             : in    std_logic := 'U';
          MGPIO26A_IN                             : in    std_logic := 'U';
          MGPIO27A_IN                             : in    std_logic := 'U';
          MGPIO28A_IN                             : in    std_logic := 'U';
          MGPIO29A_IN                             : in    std_logic := 'U';
          MGPIO2B_IN                              : in    std_logic := 'U';
          MGPIO30A_IN                             : in    std_logic := 'U';
          MGPIO31A_IN                             : in    std_logic := 'U';
          MGPIO3B_IN                              : in    std_logic := 'U';
          MGPIO4B_IN                              : in    std_logic := 'U';
          MGPIO5B_IN                              : in    std_logic := 'U';
          MGPIO6B_IN                              : in    std_logic := 'U';
          MGPIO7B_IN                              : in    std_logic := 'U';
          MGPIO8B_IN                              : in    std_logic := 'U';
          MGPIO9B_IN                              : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_CTS_MGPIO13B_IN                 : in    std_logic := 'U';
          MMUART1_DCD_MGPIO16B_IN                 : in    std_logic := 'U';
          MMUART1_DSR_MGPIO14B_IN                 : in    std_logic := 'U';
          MMUART1_DTR_MGPIO12B_IN                 : in    std_logic := 'U';
          MMUART1_RI_MGPIO15B_IN                  : in    std_logic := 'U';
          MMUART1_RTS_MGPIO11B_IN                 : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI0_SS4_MGPIO19A_IN                    : in    std_logic := 'U';
          SPI0_SS5_MGPIO20A_IN                    : in    std_logic := 'U';
          SPI0_SS6_MGPIO21A_IN                    : in    std_logic := 'U';
          SPI0_SS7_MGPIO22A_IN                    : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          USBD_DATA0_IN                           : in    std_logic := 'U';
          USBD_DATA1_IN                           : in    std_logic := 'U';
          USBD_DATA2_IN                           : in    std_logic := 'U';
          USBD_DATA3_IN                           : in    std_logic := 'U';
          USBD_DATA4_IN                           : in    std_logic := 'U';
          USBD_DATA5_IN                           : in    std_logic := 'U';
          USBD_DATA6_IN                           : in    std_logic := 'U';
          USBD_DATA7_MGPIO23B_IN                  : in    std_logic := 'U';
          USBD_DIR_IN                             : in    std_logic := 'U';
          USBD_NXT_IN                             : in    std_logic := 'U';
          USBD_STP_IN                             : in    std_logic := 'U';
          USBD_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MGPIO0B_OUT                             : out   std_logic;
          MGPIO10B_OUT                            : out   std_logic;
          MGPIO1B_OUT                             : out   std_logic;
          MGPIO25A_OUT                            : out   std_logic;
          MGPIO26A_OUT                            : out   std_logic;
          MGPIO27A_OUT                            : out   std_logic;
          MGPIO28A_OUT                            : out   std_logic;
          MGPIO29A_OUT                            : out   std_logic;
          MGPIO2B_OUT                             : out   std_logic;
          MGPIO30A_OUT                            : out   std_logic;
          MGPIO31A_OUT                            : out   std_logic;
          MGPIO3B_OUT                             : out   std_logic;
          MGPIO4B_OUT                             : out   std_logic;
          MGPIO5B_OUT                             : out   std_logic;
          MGPIO6B_OUT                             : out   std_logic;
          MGPIO7B_OUT                             : out   std_logic;
          MGPIO8B_OUT                             : out   std_logic;
          MGPIO9B_OUT                             : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_CTS_MGPIO13B_OUT                : out   std_logic;
          MMUART1_DCD_MGPIO16B_OUT                : out   std_logic;
          MMUART1_DSR_MGPIO14B_OUT                : out   std_logic;
          MMUART1_DTR_MGPIO12B_OUT                : out   std_logic;
          MMUART1_RI_MGPIO15B_OUT                 : out   std_logic;
          MMUART1_RTS_MGPIO11B_OUT                : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI0_SS4_MGPIO19A_OUT                   : out   std_logic;
          SPI0_SS5_MGPIO20A_OUT                   : out   std_logic;
          SPI0_SS6_MGPIO21A_OUT                   : out   std_logic;
          SPI0_SS7_MGPIO22A_OUT                   : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          USBD_DATA0_OUT                          : out   std_logic;
          USBD_DATA1_OUT                          : out   std_logic;
          USBD_DATA2_OUT                          : out   std_logic;
          USBD_DATA3_OUT                          : out   std_logic;
          USBD_DATA4_OUT                          : out   std_logic;
          USBD_DATA5_OUT                          : out   std_logic;
          USBD_DATA6_OUT                          : out   std_logic;
          USBD_DATA7_MGPIO23B_OUT                 : out   std_logic;
          USBD_DIR_OUT                            : out   std_logic;
          USBD_NXT_OUT                            : out   std_logic;
          USBD_STP_OUT                            : out   std_logic;
          USBD_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MGPIO0B_OE                              : out   std_logic;
          MGPIO10B_OE                             : out   std_logic;
          MGPIO1B_OE                              : out   std_logic;
          MGPIO25A_OE                             : out   std_logic;
          MGPIO26A_OE                             : out   std_logic;
          MGPIO27A_OE                             : out   std_logic;
          MGPIO28A_OE                             : out   std_logic;
          MGPIO29A_OE                             : out   std_logic;
          MGPIO2B_OE                              : out   std_logic;
          MGPIO30A_OE                             : out   std_logic;
          MGPIO31A_OE                             : out   std_logic;
          MGPIO3B_OE                              : out   std_logic;
          MGPIO4B_OE                              : out   std_logic;
          MGPIO5B_OE                              : out   std_logic;
          MGPIO6B_OE                              : out   std_logic;
          MGPIO7B_OE                              : out   std_logic;
          MGPIO8B_OE                              : out   std_logic;
          MGPIO9B_OE                              : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_CTS_MGPIO13B_OE                 : out   std_logic;
          MMUART1_DCD_MGPIO16B_OE                 : out   std_logic;
          MMUART1_DSR_MGPIO14B_OE                 : out   std_logic;
          MMUART1_DTR_MGPIO12B_OE                 : out   std_logic;
          MMUART1_RI_MGPIO15B_OE                  : out   std_logic;
          MMUART1_RTS_MGPIO11B_OE                 : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI0_SS4_MGPIO19A_OE                    : out   std_logic;
          SPI0_SS5_MGPIO20A_OE                    : out   std_logic;
          SPI0_SS6_MGPIO21A_OE                    : out   std_logic;
          SPI0_SS7_MGPIO22A_OE                    : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic;
          USBD_DATA0_OE                           : out   std_logic;
          USBD_DATA1_OE                           : out   std_logic;
          USBD_DATA2_OE                           : out   std_logic;
          USBD_DATA3_OE                           : out   std_logic;
          USBD_DATA4_OE                           : out   std_logic;
          USBD_DATA5_OE                           : out   std_logic;
          USBD_DATA6_OE                           : out   std_logic;
          USBD_DATA7_MGPIO23B_OE                  : out   std_logic;
          USBD_DIR_OE                             : out   std_logic;
          USBD_NXT_OE                             : out   std_logic;
          USBD_STP_OE                             : out   std_logic;
          USBD_XCLK_OE                            : out   std_logic
        );
  end component;

    signal \AMBA_SLAVE_0_HRDATA_S0_m[2]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[3]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[4]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[5]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[6]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[7]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[8]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[9]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[10]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[11]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[12]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[13]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[14]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[15]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[16]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[17]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[18]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[19]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[20]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[21]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[22]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[23]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[24]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[25]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[26]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[27]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[28]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[30]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[29]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[31]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[1]\, 
        \AMBA_SLAVE_0_HRDATA_S0_m[0]\, VCC_net_1, GND_net_1
         : std_logic;
    signal nc228, nc203, nc265, nc216, nc194, nc151, nc23, nc175, 
        nc250, nc58, nc116, nc74, nc133, nc238, nc167, nc84, nc39, 
        nc72, nc256, nc212, nc205, nc82, nc145, nc181, nc160, 
        nc57, nc156, nc280, nc125, nc211, nc73, nc107, nc329, 
        nc66, nc83, nc9, nc252, nc171, nc54, nc286, nc307, nc135, 
        nc41, nc100, nc270, nc52, nc251, nc186, nc29, nc269, 
        nc118, nc60, nc141, nc311, nc276, nc193, nc214, nc298, 
        nc282, nc240, nc45, nc53, nc121, nc176, nc220, nc158, 
        nc281, nc209, nc246, nc162, nc11, nc272, nc131, nc254, 
        nc267, nc96, nc79, nc226, nc146, nc230, nc89, nc119, nc48, 
        nc271, nc213, nc300, nc126, nc195, nc188, nc242, nc15, 
        nc308, nc236, nc102, nc304, nc3, nc207, nc47, nc90, nc284, 
        nc222, nc159, nc136, nc241, nc253, nc178, nc306, nc215, 
        nc59, nc221, nc232, nc274, nc18, nc44, nc117, nc189, 
        nc164, nc148, nc42, nc231, nc191, nc255, nc283, nc317, 
        nc290, nc17, nc2, nc302, nc110, nc128, nc244, nc321, nc43, 
        nc179, nc157, nc36, nc224, nc296, nc273, nc61, nc104, 
        nc138, nc14, nc285, nc303, nc150, nc331, nc196, nc234, 
        nc149, nc12, nc219, nc30, nc243, nc187, nc65, nc7, nc292, 
        nc129, nc275, nc8, nc223, nc13, nc305, nc180, nc26, nc291, 
        nc177, nc139, nc310, nc259, nc245, nc233, nc163, nc318, 
        nc268, nc112, nc68, nc49, nc314, nc217, nc170, nc91, 
        nc225, nc5, nc20, nc198, nc147, nc316, nc67, nc289, nc294, 
        nc152, nc127, nc103, nc235, nc76, nc208, nc140, nc257, 
        nc86, nc95, nc327, nc120, nc165, nc279, nc137, nc64, nc19, 
        nc312, nc70, nc182, nc62, nc199, nc80, nc130, nc287, nc98, 
        nc293, nc249, nc114, nc56, nc105, nc63, nc313, nc309, 
        nc172, nc229, nc277, nc97, nc161, nc31, nc295, nc154, 
        nc50, nc260, nc239, nc142, nc320, nc315, nc247, nc94, 
        nc197, nc328, nc122, nc266, nc35, nc324, nc4, nc227, nc92, 
        nc101, nc330, nc184, nc200, nc190, nc166, nc326, nc132, 
        nc334, nc21, nc237, nc93, nc262, nc69, nc206, nc174, nc38, 
        nc113, nc218, nc106, nc261, nc25, nc1, nc322, nc299, nc37, 
        nc202, nc144, nc153, nc46, nc258, nc71, nc124, nc332, 
        nc81, nc201, nc168, nc323, nc34, nc28, nc115, nc264, 
        nc192, nc319, nc134, nc32, nc40, nc297, nc99, nc75, nc183, 
        nc333, nc288, nc85, nc27, nc108, nc325, nc16, nc155, nc51, 
        nc301, nc33, nc204, nc173, nc278, nc169, nc78, nc263, 
        nc335, nc24, nc88, nc111, nc55, nc10, nc22, nc210, nc185, 
        nc143, nc248, nc77, nc6, nc109, nc87, nc123 : std_logic;

begin 


    MSS_ADLIB_INST_RNO_20 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1275, B => data_out_sn_N_12_mux, C => 
        N_1342, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[21]\);
    
    MSS_ADLIB_INST_RNO_23 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1278, B => data_out_sn_N_12_mux, C => 
        N_1345, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[24]\);
    
    MSS_ADLIB_INST_RNO_29 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1284, B => data_out_sn_N_12_mux, C => 
        N_1351, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[30]\);
    
    MSS_ADLIB_INST_RNO_21 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1276, B => data_out_sn_N_12_mux, C => 
        N_1343, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[22]\);
    
    MSS_ADLIB_INST_RNO : CFG4
      generic map(INIT => x"F080")

      port map(A => N_1458, B => N_1423_3, C => hready_m_xhdl339, 
        D => data_out_9_0_0, Y => \AMBA_SLAVE_0_HRDATA_S0_m[0]\);
    
    MSS_ADLIB_INST_RNO_22 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1277, B => data_out_sn_N_12_mux, C => 
        N_1344, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[23]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    MSS_ADLIB_INST_RNO_27 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1282, B => data_out_sn_N_12_mux, C => 
        N_1349, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[28]\);
    
    MSS_ADLIB_INST_RNO_10 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1265, B => data_out_sn_N_12_mux, C => 
        N_1332, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[11]\);
    
    MSS_ADLIB_INST_RNO_13 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1268, B => data_out_sn_N_12_mux, C => 
        N_1335, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[14]\);
    
    MSS_ADLIB_INST_RNO_19 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1274, B => data_out_sn_N_12_mux, C => 
        N_1341, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[20]\);
    
    MSS_ADLIB_INST_RNO_11 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1266, B => data_out_sn_N_12_mux, C => 
        N_1333, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[12]\);
    
    MSS_ADLIB_INST_RNO_12 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1267, B => data_out_sn_N_12_mux, C => 
        N_1334, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[13]\);
    
    MSS_ADLIB_INST_RNO_2 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1257, B => data_out_sn_N_12_mux, C => 
        N_1324, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[3]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    MSS_ADLIB_INST_RNO_4 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1259, B => data_out_sn_N_12_mux, C => 
        N_1326, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[5]\);
    
    MSS_ADLIB_INST_RNO_17 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1272, B => data_out_sn_N_12_mux, C => 
        N_1339, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[18]\);
    
    MSS_ADLIB_INST_RNO_7 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1262, B => data_out_sn_N_12_mux, C => 
        N_1329, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[8]\);
    
    MSS_ADLIB_INST_RNI4I5R : CFG3
      generic map(INIT => x"02")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), B
         => masterRegAddrSel, C => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, Y => 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1));
    
    MSS_ADLIB_INST : MSS_060

              generic map(INIT => "00" & x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C000000006092C0104003FFFFE4000000000000100000000F0F15C00000182DFFC010842108421000001FE34001FF8000000400000000020891007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem", RTC_MAIN_XTL_FREQ => 0.0,
         DDR_CLK_FREQ => 100.0)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => OPEN, CAN_TX_EBL_MGPIO4A_H2F_A
         => OPEN, CAN_TX_EBL_MGPIO4A_H2F_B => OPEN, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => GPIO_2_M2F_c, CLK_CONFIG_APB => OPEN, COMMS_INT => 
        OPEN, CONFIG_PRESET_N => 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        EDAC_ERROR(7) => nc228, EDAC_ERROR(6) => nc203, 
        EDAC_ERROR(5) => nc265, EDAC_ERROR(4) => nc216, 
        EDAC_ERROR(3) => nc194, EDAC_ERROR(2) => nc151, 
        EDAC_ERROR(1) => nc23, EDAC_ERROR(0) => nc175, 
        F_FM0_RDATA(31) => nc250, F_FM0_RDATA(30) => nc58, 
        F_FM0_RDATA(29) => nc116, F_FM0_RDATA(28) => nc74, 
        F_FM0_RDATA(27) => nc133, F_FM0_RDATA(26) => nc238, 
        F_FM0_RDATA(25) => nc167, F_FM0_RDATA(24) => nc84, 
        F_FM0_RDATA(23) => nc39, F_FM0_RDATA(22) => nc72, 
        F_FM0_RDATA(21) => nc256, F_FM0_RDATA(20) => nc212, 
        F_FM0_RDATA(19) => nc205, F_FM0_RDATA(18) => nc82, 
        F_FM0_RDATA(17) => nc145, F_FM0_RDATA(16) => nc181, 
        F_FM0_RDATA(15) => nc160, F_FM0_RDATA(14) => nc57, 
        F_FM0_RDATA(13) => nc156, F_FM0_RDATA(12) => nc280, 
        F_FM0_RDATA(11) => nc125, F_FM0_RDATA(10) => nc211, 
        F_FM0_RDATA(9) => nc73, F_FM0_RDATA(8) => nc107, 
        F_FM0_RDATA(7) => nc329, F_FM0_RDATA(6) => nc66, 
        F_FM0_RDATA(5) => nc83, F_FM0_RDATA(4) => nc9, 
        F_FM0_RDATA(3) => nc252, F_FM0_RDATA(2) => nc171, 
        F_FM0_RDATA(1) => nc54, F_FM0_RDATA(0) => nc286, 
        F_FM0_READYOUT => OPEN, F_FM0_RESP => OPEN, 
        F_HM0_ADDR(31) => nc307, F_HM0_ADDR(30) => nc135, 
        F_HM0_ADDR(29) => nc41, F_HM0_ADDR(28) => nc100, 
        F_HM0_ADDR(27) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_27, 
        F_HM0_ADDR(26) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_26, 
        F_HM0_ADDR(25) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, 
        F_HM0_ADDR(24) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        F_HM0_ADDR(23) => nc270, F_HM0_ADDR(22) => nc52, 
        F_HM0_ADDR(21) => nc251, F_HM0_ADDR(20) => nc186, 
        F_HM0_ADDR(19) => nc29, F_HM0_ADDR(18) => nc269, 
        F_HM0_ADDR(17) => nc118, F_HM0_ADDR(16) => nc60, 
        F_HM0_ADDR(15) => nc141, F_HM0_ADDR(14) => nc311, 
        F_HM0_ADDR(13) => nc276, F_HM0_ADDR(12) => nc193, 
        F_HM0_ADDR(11) => nc214, F_HM0_ADDR(10) => nc298, 
        F_HM0_ADDR(9) => nc282, F_HM0_ADDR(8) => nc240, 
        F_HM0_ADDR(7) => nc45, F_HM0_ADDR(6) => nc53, 
        F_HM0_ADDR(5) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        F_HM0_ADDR(4) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        F_HM0_ADDR(3) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        F_HM0_ADDR(2) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        F_HM0_ADDR(1) => nc121, F_HM0_ADDR(0) => nc176, 
        F_HM0_ENABLE => OPEN, F_HM0_SEL => OPEN, F_HM0_SIZE(1)
         => nc220, F_HM0_SIZE(0) => nc158, F_HM0_TRANS1 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        F_HM0_WDATA(31) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        F_HM0_WDATA(30) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        F_HM0_WDATA(29) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        F_HM0_WDATA(28) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        F_HM0_WDATA(27) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        F_HM0_WDATA(26) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        F_HM0_WDATA(25) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        F_HM0_WDATA(24) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        F_HM0_WDATA(23) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        F_HM0_WDATA(22) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        F_HM0_WDATA(21) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        F_HM0_WDATA(20) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        F_HM0_WDATA(19) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        F_HM0_WDATA(18) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        F_HM0_WDATA(17) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        F_HM0_WDATA(16) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        F_HM0_WDATA(15) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        F_HM0_WDATA(14) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        F_HM0_WDATA(13) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        F_HM0_WDATA(12) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        F_HM0_WDATA(11) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        F_HM0_WDATA(10) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        F_HM0_WDATA(9) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        F_HM0_WDATA(8) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        F_HM0_WDATA(7) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        F_HM0_WDATA(6) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        F_HM0_WDATA(5) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        F_HM0_WDATA(4) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        F_HM0_WDATA(3) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        F_HM0_WDATA(2) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        F_HM0_WDATA(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        F_HM0_WDATA(0) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        F_HM0_WRITE => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        FAB_CHRGVBUS => OPEN, FAB_DISCHRGVBUS => OPEN, 
        FAB_DMPULLDOWN => OPEN, FAB_DPPULLDOWN => OPEN, 
        FAB_DRVVBUS => OPEN, FAB_IDPULLUP => OPEN, FAB_OPMODE(1)
         => nc281, FAB_OPMODE(0) => nc209, FAB_SUSPENDM => OPEN, 
        FAB_TERMSEL => OPEN, FAB_TXVALID => OPEN, FAB_VCONTROL(3)
         => nc246, FAB_VCONTROL(2) => nc162, FAB_VCONTROL(1) => 
        nc11, FAB_VCONTROL(0) => nc272, FAB_VCONTROLLOADM => OPEN, 
        FAB_XCVRSEL(1) => nc131, FAB_XCVRSEL(0) => nc254, 
        FAB_XDATAOUT(7) => nc267, FAB_XDATAOUT(6) => nc96, 
        FAB_XDATAOUT(5) => nc79, FAB_XDATAOUT(4) => nc226, 
        FAB_XDATAOUT(3) => nc146, FAB_XDATAOUT(2) => nc230, 
        FAB_XDATAOUT(1) => nc89, FAB_XDATAOUT(0) => nc119, 
        FACC_GLMUX_SEL => OPEN, FIC32_0_MASTER(1) => nc48, 
        FIC32_0_MASTER(0) => nc271, FIC32_1_MASTER(1) => nc213, 
        FIC32_1_MASTER(0) => nc300, FPGA_RESET_N => 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, GTX_CLK => 
        OPEN, H2F_INTERRUPT(15) => nc126, H2F_INTERRUPT(14) => 
        nc195, H2F_INTERRUPT(13) => nc188, H2F_INTERRUPT(12) => 
        nc242, H2F_INTERRUPT(11) => nc15, H2F_INTERRUPT(10) => 
        nc308, H2F_INTERRUPT(9) => nc236, H2F_INTERRUPT(8) => 
        nc102, H2F_INTERRUPT(7) => nc304, H2F_INTERRUPT(6) => nc3, 
        H2F_INTERRUPT(5) => nc207, H2F_INTERRUPT(4) => nc47, 
        H2F_INTERRUPT(3) => nc90, H2F_INTERRUPT(2) => nc284, 
        H2F_INTERRUPT(1) => nc222, H2F_INTERRUPT(0) => nc159, 
        H2F_NMI => OPEN, H2FCALIB => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_A => OPEN, I2C0_SCL_MGPIO31B_H2F_B
         => OPEN, I2C0_SDA_MGPIO30B_H2F_A => OPEN, 
        I2C0_SDA_MGPIO30B_H2F_B => OPEN, I2C1_SCL_MGPIO1A_H2F_A
         => OPEN, I2C1_SCL_MGPIO1A_H2F_B => GPIO_1_M2F_c, 
        I2C1_SDA_MGPIO0A_H2F_A => OPEN, I2C1_SDA_MGPIO0A_H2F_B
         => GPIO_0_M2F_c, MDCF => OPEN, MDOENF => OPEN, MDOF => 
        OPEN, MMUART0_CTS_MGPIO19B_H2F_A => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => OPEN, MPLL_LOCK => OPEN, 
        PER2_FABRIC_PADDR(15) => nc136, PER2_FABRIC_PADDR(14) => 
        nc241, PER2_FABRIC_PADDR(13) => nc253, 
        PER2_FABRIC_PADDR(12) => nc178, PER2_FABRIC_PADDR(11) => 
        nc306, PER2_FABRIC_PADDR(10) => nc215, 
        PER2_FABRIC_PADDR(9) => nc59, PER2_FABRIC_PADDR(8) => 
        nc221, PER2_FABRIC_PADDR(7) => nc232, 
        PER2_FABRIC_PADDR(6) => nc274, PER2_FABRIC_PADDR(5) => 
        nc18, PER2_FABRIC_PADDR(4) => nc44, PER2_FABRIC_PADDR(3)
         => nc117, PER2_FABRIC_PADDR(2) => nc189, 
        PER2_FABRIC_PENABLE => OPEN, PER2_FABRIC_PSEL => OPEN, 
        PER2_FABRIC_PWDATA(31) => nc164, PER2_FABRIC_PWDATA(30)
         => nc148, PER2_FABRIC_PWDATA(29) => nc42, 
        PER2_FABRIC_PWDATA(28) => nc231, PER2_FABRIC_PWDATA(27)
         => nc191, PER2_FABRIC_PWDATA(26) => nc255, 
        PER2_FABRIC_PWDATA(25) => nc283, PER2_FABRIC_PWDATA(24)
         => nc317, PER2_FABRIC_PWDATA(23) => nc290, 
        PER2_FABRIC_PWDATA(22) => nc17, PER2_FABRIC_PWDATA(21)
         => nc2, PER2_FABRIC_PWDATA(20) => nc302, 
        PER2_FABRIC_PWDATA(19) => nc110, PER2_FABRIC_PWDATA(18)
         => nc128, PER2_FABRIC_PWDATA(17) => nc244, 
        PER2_FABRIC_PWDATA(16) => nc321, PER2_FABRIC_PWDATA(15)
         => nc43, PER2_FABRIC_PWDATA(14) => nc179, 
        PER2_FABRIC_PWDATA(13) => nc157, PER2_FABRIC_PWDATA(12)
         => nc36, PER2_FABRIC_PWDATA(11) => nc224, 
        PER2_FABRIC_PWDATA(10) => nc296, PER2_FABRIC_PWDATA(9)
         => nc273, PER2_FABRIC_PWDATA(8) => nc61, 
        PER2_FABRIC_PWDATA(7) => nc104, PER2_FABRIC_PWDATA(6) => 
        nc138, PER2_FABRIC_PWDATA(5) => nc14, 
        PER2_FABRIC_PWDATA(4) => nc285, PER2_FABRIC_PWDATA(3) => 
        nc303, PER2_FABRIC_PWDATA(2) => nc150, 
        PER2_FABRIC_PWDATA(1) => nc331, PER2_FABRIC_PWDATA(0) => 
        nc196, PER2_FABRIC_PWRITE => OPEN, RTC_MATCH => OPEN, 
        SLEEPDEEP => OPEN, SLEEPHOLDACK => OPEN, SLEEPING => OPEN, 
        SMBALERT_NO0 => OPEN, SMBALERT_NO1 => OPEN, SMBSUS_NO0
         => OPEN, SMBSUS_NO1 => OPEN, SPI0_CLK_OUT => OPEN, 
        SPI0_SDI_MGPIO5A_H2F_A => OPEN, SPI0_SDI_MGPIO5A_H2F_B
         => OPEN, SPI0_SDO_MGPIO6A_H2F_A => OPEN, 
        SPI0_SDO_MGPIO6A_H2F_B => OPEN, SPI0_SS0_MGPIO7A_H2F_A
         => OPEN, SPI0_SS0_MGPIO7A_H2F_B => OPEN, 
        SPI0_SS1_MGPIO8A_H2F_A => OPEN, SPI0_SS1_MGPIO8A_H2F_B
         => OPEN, SPI0_SS2_MGPIO9A_H2F_A => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_B => OPEN, SPI0_SS3_MGPIO10A_H2F_A
         => OPEN, SPI0_SS3_MGPIO10A_H2F_B => OPEN, 
        SPI0_SS4_MGPIO19A_H2F_A => OPEN, SPI0_SS5_MGPIO20A_H2F_A
         => OPEN, SPI0_SS6_MGPIO21A_H2F_A => OPEN, 
        SPI0_SS7_MGPIO22A_H2F_A => OPEN, SPI1_CLK_OUT => OPEN, 
        SPI1_SDI_MGPIO11A_H2F_A => OPEN, SPI1_SDI_MGPIO11A_H2F_B
         => OPEN, SPI1_SDO_MGPIO12A_H2F_A => OPEN, 
        SPI1_SDO_MGPIO12A_H2F_B => OPEN, SPI1_SS0_MGPIO13A_H2F_A
         => OPEN, SPI1_SS0_MGPIO13A_H2F_B => OPEN, 
        SPI1_SS1_MGPIO14A_H2F_A => OPEN, SPI1_SS1_MGPIO14A_H2F_B
         => OPEN, SPI1_SS2_MGPIO15A_H2F_A => OPEN, 
        SPI1_SS2_MGPIO15A_H2F_B => OPEN, SPI1_SS3_MGPIO16A_H2F_A
         => OPEN, SPI1_SS3_MGPIO16A_H2F_B => OPEN, 
        SPI1_SS4_MGPIO17A_H2F_A => OPEN, SPI1_SS5_MGPIO18A_H2F_A
         => OPEN, SPI1_SS6_MGPIO23A_H2F_A => OPEN, 
        SPI1_SS7_MGPIO24A_H2F_A => OPEN, TCGF(9) => nc234, 
        TCGF(8) => nc149, TCGF(7) => nc12, TCGF(6) => nc219, 
        TCGF(5) => nc30, TCGF(4) => nc243, TCGF(3) => nc187, 
        TCGF(2) => nc65, TCGF(1) => nc7, TCGF(0) => nc292, 
        TRACECLK => OPEN, TRACEDATA(3) => nc129, TRACEDATA(2) => 
        nc275, TRACEDATA(1) => nc8, TRACEDATA(0) => nc223, TX_CLK
         => OPEN, TX_ENF => OPEN, TX_ERRF => OPEN, TXCTL_EN_RIF
         => OPEN, TXD_RIF(3) => nc13, TXD_RIF(2) => nc305, 
        TXD_RIF(1) => nc180, TXD_RIF(0) => nc26, TXDF(7) => nc291, 
        TXDF(6) => nc177, TXDF(5) => nc139, TXDF(4) => nc310, 
        TXDF(3) => nc259, TXDF(2) => nc245, TXDF(1) => nc233, 
        TXDF(0) => nc163, TXEV => OPEN, WDOGTIMEOUT => OPEN, 
        F_ARREADY_HREADYOUT1 => OPEN, F_AWREADY_HREADYOUT0 => 
        OPEN, F_BID(3) => nc318, F_BID(2) => nc268, F_BID(1) => 
        nc112, F_BID(0) => nc68, F_BRESP_HRESP0(1) => nc49, 
        F_BRESP_HRESP0(0) => nc314, F_BVALID => OPEN, 
        F_RDATA_HRDATA01(63) => nc217, F_RDATA_HRDATA01(62) => 
        nc170, F_RDATA_HRDATA01(61) => nc91, F_RDATA_HRDATA01(60)
         => nc225, F_RDATA_HRDATA01(59) => nc5, 
        F_RDATA_HRDATA01(58) => nc20, F_RDATA_HRDATA01(57) => 
        nc198, F_RDATA_HRDATA01(56) => nc147, 
        F_RDATA_HRDATA01(55) => nc316, F_RDATA_HRDATA01(54) => 
        nc67, F_RDATA_HRDATA01(53) => nc289, F_RDATA_HRDATA01(52)
         => nc294, F_RDATA_HRDATA01(51) => nc152, 
        F_RDATA_HRDATA01(50) => nc127, F_RDATA_HRDATA01(49) => 
        nc103, F_RDATA_HRDATA01(48) => nc235, 
        F_RDATA_HRDATA01(47) => nc76, F_RDATA_HRDATA01(46) => 
        nc208, F_RDATA_HRDATA01(45) => nc140, 
        F_RDATA_HRDATA01(44) => nc257, F_RDATA_HRDATA01(43) => 
        nc86, F_RDATA_HRDATA01(42) => nc95, F_RDATA_HRDATA01(41)
         => nc327, F_RDATA_HRDATA01(40) => nc120, 
        F_RDATA_HRDATA01(39) => nc165, F_RDATA_HRDATA01(38) => 
        nc279, F_RDATA_HRDATA01(37) => nc137, 
        F_RDATA_HRDATA01(36) => nc64, F_RDATA_HRDATA01(35) => 
        nc19, F_RDATA_HRDATA01(34) => nc312, F_RDATA_HRDATA01(33)
         => nc70, F_RDATA_HRDATA01(32) => nc182, 
        F_RDATA_HRDATA01(31) => nc62, F_RDATA_HRDATA01(30) => 
        nc199, F_RDATA_HRDATA01(29) => nc80, F_RDATA_HRDATA01(28)
         => nc130, F_RDATA_HRDATA01(27) => nc287, 
        F_RDATA_HRDATA01(26) => nc98, F_RDATA_HRDATA01(25) => 
        nc293, F_RDATA_HRDATA01(24) => nc249, 
        F_RDATA_HRDATA01(23) => nc114, F_RDATA_HRDATA01(22) => 
        nc56, F_RDATA_HRDATA01(21) => nc105, F_RDATA_HRDATA01(20)
         => nc63, F_RDATA_HRDATA01(19) => nc313, 
        F_RDATA_HRDATA01(18) => nc309, F_RDATA_HRDATA01(17) => 
        nc172, F_RDATA_HRDATA01(16) => nc229, 
        F_RDATA_HRDATA01(15) => nc277, F_RDATA_HRDATA01(14) => 
        nc97, F_RDATA_HRDATA01(13) => nc161, F_RDATA_HRDATA01(12)
         => nc31, F_RDATA_HRDATA01(11) => nc295, 
        F_RDATA_HRDATA01(10) => nc154, F_RDATA_HRDATA01(9) => 
        nc50, F_RDATA_HRDATA01(8) => nc260, F_RDATA_HRDATA01(7)
         => nc239, F_RDATA_HRDATA01(6) => nc142, 
        F_RDATA_HRDATA01(5) => nc320, F_RDATA_HRDATA01(4) => 
        nc315, F_RDATA_HRDATA01(3) => nc247, F_RDATA_HRDATA01(2)
         => nc94, F_RDATA_HRDATA01(1) => nc197, 
        F_RDATA_HRDATA01(0) => nc328, F_RID(3) => nc122, F_RID(2)
         => nc266, F_RID(1) => nc35, F_RID(0) => nc324, F_RLAST
         => OPEN, F_RRESP_HRESP1(1) => nc4, F_RRESP_HRESP1(0) => 
        nc227, F_RVALID => OPEN, F_WREADY => OPEN, 
        MDDR_FABRIC_PRDATA(15) => nc92, MDDR_FABRIC_PRDATA(14)
         => nc101, MDDR_FABRIC_PRDATA(13) => nc330, 
        MDDR_FABRIC_PRDATA(12) => nc184, MDDR_FABRIC_PRDATA(11)
         => nc200, MDDR_FABRIC_PRDATA(10) => nc190, 
        MDDR_FABRIC_PRDATA(9) => nc166, MDDR_FABRIC_PRDATA(8) => 
        nc326, MDDR_FABRIC_PRDATA(7) => nc132, 
        MDDR_FABRIC_PRDATA(6) => nc334, MDDR_FABRIC_PRDATA(5) => 
        nc21, MDDR_FABRIC_PRDATA(4) => nc237, 
        MDDR_FABRIC_PRDATA(3) => nc93, MDDR_FABRIC_PRDATA(2) => 
        nc262, MDDR_FABRIC_PRDATA(1) => nc69, 
        MDDR_FABRIC_PRDATA(0) => nc206, MDDR_FABRIC_PREADY => 
        OPEN, MDDR_FABRIC_PSLVERR => OPEN, CAN_RXBUS_F2H_SCP => 
        VCC_net_1, CAN_TX_EBL_F2H_SCP => VCC_net_1, 
        CAN_TXBUS_F2H_SCP => VCC_net_1, COLF => VCC_net_1, CRSF
         => VCC_net_1, F2_DMAREADY(1) => VCC_net_1, 
        F2_DMAREADY(0) => VCC_net_1, F2H_INTERRUPT(15) => 
        GND_net_1, F2H_INTERRUPT(14) => GND_net_1, 
        F2H_INTERRUPT(13) => GND_net_1, F2H_INTERRUPT(12) => 
        GND_net_1, F2H_INTERRUPT(11) => GND_net_1, 
        F2H_INTERRUPT(10) => GND_net_1, F2H_INTERRUPT(9) => 
        GND_net_1, F2H_INTERRUPT(8) => GND_net_1, 
        F2H_INTERRUPT(7) => GND_net_1, F2H_INTERRUPT(6) => 
        GND_net_1, F2H_INTERRUPT(5) => GND_net_1, 
        F2H_INTERRUPT(4) => GND_net_1, F2H_INTERRUPT(3) => 
        GND_net_1, F2H_INTERRUPT(2) => GND_net_1, 
        F2H_INTERRUPT(1) => GND_net_1, F2H_INTERRUPT(0) => 
        GND_net_1, F2HCALIB => VCC_net_1, F_DMAREADY(1) => 
        VCC_net_1, F_DMAREADY(0) => VCC_net_1, F_FM0_ADDR(31) => 
        GND_net_1, F_FM0_ADDR(30) => GND_net_1, F_FM0_ADDR(29)
         => GND_net_1, F_FM0_ADDR(28) => GND_net_1, 
        F_FM0_ADDR(27) => GND_net_1, F_FM0_ADDR(26) => GND_net_1, 
        F_FM0_ADDR(25) => GND_net_1, F_FM0_ADDR(24) => GND_net_1, 
        F_FM0_ADDR(23) => GND_net_1, F_FM0_ADDR(22) => GND_net_1, 
        F_FM0_ADDR(21) => GND_net_1, F_FM0_ADDR(20) => GND_net_1, 
        F_FM0_ADDR(19) => GND_net_1, F_FM0_ADDR(18) => GND_net_1, 
        F_FM0_ADDR(17) => GND_net_1, F_FM0_ADDR(16) => GND_net_1, 
        F_FM0_ADDR(15) => GND_net_1, F_FM0_ADDR(14) => GND_net_1, 
        F_FM0_ADDR(13) => GND_net_1, F_FM0_ADDR(12) => GND_net_1, 
        F_FM0_ADDR(11) => GND_net_1, F_FM0_ADDR(10) => GND_net_1, 
        F_FM0_ADDR(9) => GND_net_1, F_FM0_ADDR(8) => GND_net_1, 
        F_FM0_ADDR(7) => GND_net_1, F_FM0_ADDR(6) => GND_net_1, 
        F_FM0_ADDR(5) => GND_net_1, F_FM0_ADDR(4) => GND_net_1, 
        F_FM0_ADDR(3) => GND_net_1, F_FM0_ADDR(2) => GND_net_1, 
        F_FM0_ADDR(1) => GND_net_1, F_FM0_ADDR(0) => GND_net_1, 
        F_FM0_ENABLE => GND_net_1, F_FM0_MASTLOCK => GND_net_1, 
        F_FM0_READY => VCC_net_1, F_FM0_SEL => GND_net_1, 
        F_FM0_SIZE(1) => GND_net_1, F_FM0_SIZE(0) => GND_net_1, 
        F_FM0_TRANS1 => GND_net_1, F_FM0_WDATA(31) => GND_net_1, 
        F_FM0_WDATA(30) => GND_net_1, F_FM0_WDATA(29) => 
        GND_net_1, F_FM0_WDATA(28) => GND_net_1, F_FM0_WDATA(27)
         => GND_net_1, F_FM0_WDATA(26) => GND_net_1, 
        F_FM0_WDATA(25) => GND_net_1, F_FM0_WDATA(24) => 
        GND_net_1, F_FM0_WDATA(23) => GND_net_1, F_FM0_WDATA(22)
         => GND_net_1, F_FM0_WDATA(21) => GND_net_1, 
        F_FM0_WDATA(20) => GND_net_1, F_FM0_WDATA(19) => 
        GND_net_1, F_FM0_WDATA(18) => GND_net_1, F_FM0_WDATA(17)
         => GND_net_1, F_FM0_WDATA(16) => GND_net_1, 
        F_FM0_WDATA(15) => GND_net_1, F_FM0_WDATA(14) => 
        GND_net_1, F_FM0_WDATA(13) => GND_net_1, F_FM0_WDATA(12)
         => GND_net_1, F_FM0_WDATA(11) => GND_net_1, 
        F_FM0_WDATA(10) => GND_net_1, F_FM0_WDATA(9) => GND_net_1, 
        F_FM0_WDATA(8) => GND_net_1, F_FM0_WDATA(7) => GND_net_1, 
        F_FM0_WDATA(6) => GND_net_1, F_FM0_WDATA(5) => GND_net_1, 
        F_FM0_WDATA(4) => GND_net_1, F_FM0_WDATA(3) => GND_net_1, 
        F_FM0_WDATA(2) => GND_net_1, F_FM0_WDATA(1) => GND_net_1, 
        F_FM0_WDATA(0) => GND_net_1, F_FM0_WRITE => GND_net_1, 
        F_HM0_RDATA(31) => \AMBA_SLAVE_0_HRDATA_S0_m[31]\, 
        F_HM0_RDATA(30) => \AMBA_SLAVE_0_HRDATA_S0_m[30]\, 
        F_HM0_RDATA(29) => \AMBA_SLAVE_0_HRDATA_S0_m[29]\, 
        F_HM0_RDATA(28) => \AMBA_SLAVE_0_HRDATA_S0_m[28]\, 
        F_HM0_RDATA(27) => \AMBA_SLAVE_0_HRDATA_S0_m[27]\, 
        F_HM0_RDATA(26) => \AMBA_SLAVE_0_HRDATA_S0_m[26]\, 
        F_HM0_RDATA(25) => \AMBA_SLAVE_0_HRDATA_S0_m[25]\, 
        F_HM0_RDATA(24) => \AMBA_SLAVE_0_HRDATA_S0_m[24]\, 
        F_HM0_RDATA(23) => \AMBA_SLAVE_0_HRDATA_S0_m[23]\, 
        F_HM0_RDATA(22) => \AMBA_SLAVE_0_HRDATA_S0_m[22]\, 
        F_HM0_RDATA(21) => \AMBA_SLAVE_0_HRDATA_S0_m[21]\, 
        F_HM0_RDATA(20) => \AMBA_SLAVE_0_HRDATA_S0_m[20]\, 
        F_HM0_RDATA(19) => \AMBA_SLAVE_0_HRDATA_S0_m[19]\, 
        F_HM0_RDATA(18) => \AMBA_SLAVE_0_HRDATA_S0_m[18]\, 
        F_HM0_RDATA(17) => \AMBA_SLAVE_0_HRDATA_S0_m[17]\, 
        F_HM0_RDATA(16) => \AMBA_SLAVE_0_HRDATA_S0_m[16]\, 
        F_HM0_RDATA(15) => \AMBA_SLAVE_0_HRDATA_S0_m[15]\, 
        F_HM0_RDATA(14) => \AMBA_SLAVE_0_HRDATA_S0_m[14]\, 
        F_HM0_RDATA(13) => \AMBA_SLAVE_0_HRDATA_S0_m[13]\, 
        F_HM0_RDATA(12) => \AMBA_SLAVE_0_HRDATA_S0_m[12]\, 
        F_HM0_RDATA(11) => \AMBA_SLAVE_0_HRDATA_S0_m[11]\, 
        F_HM0_RDATA(10) => \AMBA_SLAVE_0_HRDATA_S0_m[10]\, 
        F_HM0_RDATA(9) => \AMBA_SLAVE_0_HRDATA_S0_m[9]\, 
        F_HM0_RDATA(8) => \AMBA_SLAVE_0_HRDATA_S0_m[8]\, 
        F_HM0_RDATA(7) => \AMBA_SLAVE_0_HRDATA_S0_m[7]\, 
        F_HM0_RDATA(6) => \AMBA_SLAVE_0_HRDATA_S0_m[6]\, 
        F_HM0_RDATA(5) => \AMBA_SLAVE_0_HRDATA_S0_m[5]\, 
        F_HM0_RDATA(4) => \AMBA_SLAVE_0_HRDATA_S0_m[4]\, 
        F_HM0_RDATA(3) => \AMBA_SLAVE_0_HRDATA_S0_m[3]\, 
        F_HM0_RDATA(2) => \AMBA_SLAVE_0_HRDATA_S0_m[2]\, 
        F_HM0_RDATA(1) => \AMBA_SLAVE_0_HRDATA_S0_m[1]\, 
        F_HM0_RDATA(0) => \AMBA_SLAVE_0_HRDATA_S0_m[0]\, 
        F_HM0_READY => N_23_i_0, F_HM0_RESP => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        FAB_AVALID => VCC_net_1, FAB_HOSTDISCON => VCC_net_1, 
        FAB_IDDIG => VCC_net_1, FAB_LINESTATE(1) => VCC_net_1, 
        FAB_LINESTATE(0) => VCC_net_1, FAB_M3_RESET_N => 
        VCC_net_1, FAB_PLL_LOCK => FIC_0_LOCK, FAB_RXACTIVE => 
        VCC_net_1, FAB_RXERROR => VCC_net_1, FAB_RXVALID => 
        VCC_net_1, FAB_RXVALIDH => GND_net_1, FAB_SESSEND => 
        VCC_net_1, FAB_TXREADY => VCC_net_1, FAB_VBUSVALID => 
        VCC_net_1, FAB_VSTATUS(7) => VCC_net_1, FAB_VSTATUS(6)
         => VCC_net_1, FAB_VSTATUS(5) => VCC_net_1, 
        FAB_VSTATUS(4) => VCC_net_1, FAB_VSTATUS(3) => VCC_net_1, 
        FAB_VSTATUS(2) => VCC_net_1, FAB_VSTATUS(1) => VCC_net_1, 
        FAB_VSTATUS(0) => VCC_net_1, FAB_XDATAIN(7) => VCC_net_1, 
        FAB_XDATAIN(6) => VCC_net_1, FAB_XDATAIN(5) => VCC_net_1, 
        FAB_XDATAIN(4) => VCC_net_1, FAB_XDATAIN(3) => VCC_net_1, 
        FAB_XDATAIN(2) => VCC_net_1, FAB_XDATAIN(1) => VCC_net_1, 
        FAB_XDATAIN(0) => VCC_net_1, GTX_CLKPF => VCC_net_1, 
        I2C0_BCLK => VCC_net_1, I2C0_SCL_F2H_SCP => VCC_net_1, 
        I2C0_SDA_F2H_SCP => VCC_net_1, I2C1_BCLK => VCC_net_1, 
        I2C1_SCL_F2H_SCP => VCC_net_1, I2C1_SDA_F2H_SCP => 
        VCC_net_1, MDIF => VCC_net_1, MGPIO0A_F2H_GPIN => 
        VCC_net_1, MGPIO10A_F2H_GPIN => VCC_net_1, 
        MGPIO11A_F2H_GPIN => VCC_net_1, MGPIO11B_F2H_GPIN => 
        VCC_net_1, MGPIO12A_F2H_GPIN => VCC_net_1, 
        MGPIO13A_F2H_GPIN => VCC_net_1, MGPIO14A_F2H_GPIN => 
        VCC_net_1, MGPIO15A_F2H_GPIN => VCC_net_1, 
        MGPIO16A_F2H_GPIN => VCC_net_1, MGPIO17B_F2H_GPIN => 
        VCC_net_1, MGPIO18B_F2H_GPIN => VCC_net_1, 
        MGPIO19B_F2H_GPIN => VCC_net_1, MGPIO1A_F2H_GPIN => 
        VCC_net_1, MGPIO20B_F2H_GPIN => VCC_net_1, 
        MGPIO21B_F2H_GPIN => VCC_net_1, MGPIO22B_F2H_GPIN => 
        VCC_net_1, MGPIO24B_F2H_GPIN => VCC_net_1, 
        MGPIO25B_F2H_GPIN => VCC_net_1, MGPIO26B_F2H_GPIN => 
        VCC_net_1, MGPIO27B_F2H_GPIN => VCC_net_1, 
        MGPIO28B_F2H_GPIN => VCC_net_1, MGPIO29B_F2H_GPIN => 
        VCC_net_1, MGPIO2A_F2H_GPIN => VCC_net_1, 
        MGPIO30B_F2H_GPIN => VCC_net_1, MGPIO31B_F2H_GPIN => 
        VCC_net_1, MGPIO3A_F2H_GPIN => VCC_net_1, 
        MGPIO4A_F2H_GPIN => VCC_net_1, MGPIO5A_F2H_GPIN => 
        VCC_net_1, MGPIO6A_F2H_GPIN => VCC_net_1, 
        MGPIO7A_F2H_GPIN => VCC_net_1, MGPIO8A_F2H_GPIN => 
        VCC_net_1, MGPIO9A_F2H_GPIN => VCC_net_1, 
        MMUART0_CTS_F2H_SCP => VCC_net_1, MMUART0_DCD_F2H_SCP => 
        VCC_net_1, MMUART0_DSR_F2H_SCP => VCC_net_1, 
        MMUART0_DTR_F2H_SCP => VCC_net_1, MMUART0_RI_F2H_SCP => 
        VCC_net_1, MMUART0_RTS_F2H_SCP => VCC_net_1, 
        MMUART0_RXD_F2H_SCP => VCC_net_1, MMUART0_SCK_F2H_SCP => 
        VCC_net_1, MMUART0_TXD_F2H_SCP => VCC_net_1, 
        MMUART1_CTS_F2H_SCP => VCC_net_1, MMUART1_DCD_F2H_SCP => 
        VCC_net_1, MMUART1_DSR_F2H_SCP => VCC_net_1, 
        MMUART1_RI_F2H_SCP => VCC_net_1, MMUART1_RTS_F2H_SCP => 
        VCC_net_1, MMUART1_RXD_F2H_SCP => VCC_net_1, 
        MMUART1_SCK_F2H_SCP => VCC_net_1, MMUART1_TXD_F2H_SCP => 
        VCC_net_1, PER2_FABRIC_PRDATA(31) => GND_net_1, 
        PER2_FABRIC_PRDATA(30) => GND_net_1, 
        PER2_FABRIC_PRDATA(29) => GND_net_1, 
        PER2_FABRIC_PRDATA(28) => GND_net_1, 
        PER2_FABRIC_PRDATA(27) => GND_net_1, 
        PER2_FABRIC_PRDATA(26) => GND_net_1, 
        PER2_FABRIC_PRDATA(25) => GND_net_1, 
        PER2_FABRIC_PRDATA(24) => GND_net_1, 
        PER2_FABRIC_PRDATA(23) => GND_net_1, 
        PER2_FABRIC_PRDATA(22) => GND_net_1, 
        PER2_FABRIC_PRDATA(21) => GND_net_1, 
        PER2_FABRIC_PRDATA(20) => GND_net_1, 
        PER2_FABRIC_PRDATA(19) => GND_net_1, 
        PER2_FABRIC_PRDATA(18) => GND_net_1, 
        PER2_FABRIC_PRDATA(17) => GND_net_1, 
        PER2_FABRIC_PRDATA(16) => GND_net_1, 
        PER2_FABRIC_PRDATA(15) => GND_net_1, 
        PER2_FABRIC_PRDATA(14) => GND_net_1, 
        PER2_FABRIC_PRDATA(13) => GND_net_1, 
        PER2_FABRIC_PRDATA(12) => GND_net_1, 
        PER2_FABRIC_PRDATA(11) => GND_net_1, 
        PER2_FABRIC_PRDATA(10) => GND_net_1, 
        PER2_FABRIC_PRDATA(9) => GND_net_1, PER2_FABRIC_PRDATA(8)
         => GND_net_1, PER2_FABRIC_PRDATA(7) => GND_net_1, 
        PER2_FABRIC_PRDATA(6) => GND_net_1, PER2_FABRIC_PRDATA(5)
         => GND_net_1, PER2_FABRIC_PRDATA(4) => GND_net_1, 
        PER2_FABRIC_PRDATA(3) => GND_net_1, PER2_FABRIC_PRDATA(2)
         => GND_net_1, PER2_FABRIC_PRDATA(1) => GND_net_1, 
        PER2_FABRIC_PRDATA(0) => GND_net_1, PER2_FABRIC_PREADY
         => VCC_net_1, PER2_FABRIC_PSLVERR => GND_net_1, RCGF(9)
         => VCC_net_1, RCGF(8) => VCC_net_1, RCGF(7) => VCC_net_1, 
        RCGF(6) => VCC_net_1, RCGF(5) => VCC_net_1, RCGF(4) => 
        VCC_net_1, RCGF(3) => VCC_net_1, RCGF(2) => VCC_net_1, 
        RCGF(1) => VCC_net_1, RCGF(0) => VCC_net_1, RX_CLKPF => 
        VCC_net_1, RX_DVF => VCC_net_1, RX_ERRF => VCC_net_1, 
        RX_EV => VCC_net_1, RXDF(7) => VCC_net_1, RXDF(6) => 
        VCC_net_1, RXDF(5) => VCC_net_1, RXDF(4) => VCC_net_1, 
        RXDF(3) => VCC_net_1, RXDF(2) => VCC_net_1, RXDF(1) => 
        VCC_net_1, RXDF(0) => VCC_net_1, SLEEPHOLDREQ => 
        GND_net_1, SMBALERT_NI0 => VCC_net_1, SMBALERT_NI1 => 
        VCC_net_1, SMBSUS_NI0 => VCC_net_1, SMBSUS_NI1 => 
        VCC_net_1, SPI0_CLK_IN => VCC_net_1, SPI0_SDI_F2H_SCP => 
        VCC_net_1, SPI0_SDO_F2H_SCP => VCC_net_1, 
        SPI0_SS0_F2H_SCP => VCC_net_1, SPI0_SS1_F2H_SCP => 
        VCC_net_1, SPI0_SS2_F2H_SCP => VCC_net_1, 
        SPI0_SS3_F2H_SCP => VCC_net_1, SPI1_CLK_IN => VCC_net_1, 
        SPI1_SDI_F2H_SCP => VCC_net_1, SPI1_SDO_F2H_SCP => 
        VCC_net_1, SPI1_SS0_F2H_SCP => VCC_net_1, 
        SPI1_SS1_F2H_SCP => VCC_net_1, SPI1_SS2_F2H_SCP => 
        VCC_net_1, SPI1_SS3_F2H_SCP => VCC_net_1, TX_CLKPF => 
        VCC_net_1, USER_MSS_GPIO_RESET_N => VCC_net_1, 
        USER_MSS_RESET_N => VCC_net_1, XCLK_FAB => VCC_net_1, 
        CLK_BASE => sha256_system_sb_0_FIC_0_CLK, CLK_MDDR_APB
         => VCC_net_1, F_ARADDR_HADDR1(31) => VCC_net_1, 
        F_ARADDR_HADDR1(30) => VCC_net_1, F_ARADDR_HADDR1(29) => 
        VCC_net_1, F_ARADDR_HADDR1(28) => VCC_net_1, 
        F_ARADDR_HADDR1(27) => VCC_net_1, F_ARADDR_HADDR1(26) => 
        VCC_net_1, F_ARADDR_HADDR1(25) => VCC_net_1, 
        F_ARADDR_HADDR1(24) => VCC_net_1, F_ARADDR_HADDR1(23) => 
        VCC_net_1, F_ARADDR_HADDR1(22) => VCC_net_1, 
        F_ARADDR_HADDR1(21) => VCC_net_1, F_ARADDR_HADDR1(20) => 
        VCC_net_1, F_ARADDR_HADDR1(19) => VCC_net_1, 
        F_ARADDR_HADDR1(18) => VCC_net_1, F_ARADDR_HADDR1(17) => 
        VCC_net_1, F_ARADDR_HADDR1(16) => VCC_net_1, 
        F_ARADDR_HADDR1(15) => VCC_net_1, F_ARADDR_HADDR1(14) => 
        VCC_net_1, F_ARADDR_HADDR1(13) => VCC_net_1, 
        F_ARADDR_HADDR1(12) => VCC_net_1, F_ARADDR_HADDR1(11) => 
        VCC_net_1, F_ARADDR_HADDR1(10) => VCC_net_1, 
        F_ARADDR_HADDR1(9) => VCC_net_1, F_ARADDR_HADDR1(8) => 
        VCC_net_1, F_ARADDR_HADDR1(7) => VCC_net_1, 
        F_ARADDR_HADDR1(6) => VCC_net_1, F_ARADDR_HADDR1(5) => 
        VCC_net_1, F_ARADDR_HADDR1(4) => VCC_net_1, 
        F_ARADDR_HADDR1(3) => VCC_net_1, F_ARADDR_HADDR1(2) => 
        VCC_net_1, F_ARADDR_HADDR1(1) => VCC_net_1, 
        F_ARADDR_HADDR1(0) => VCC_net_1, F_ARBURST_HTRANS1(1) => 
        GND_net_1, F_ARBURST_HTRANS1(0) => GND_net_1, 
        F_ARID_HSEL1(3) => GND_net_1, F_ARID_HSEL1(2) => 
        GND_net_1, F_ARID_HSEL1(1) => GND_net_1, F_ARID_HSEL1(0)
         => GND_net_1, F_ARLEN_HBURST1(3) => GND_net_1, 
        F_ARLEN_HBURST1(2) => GND_net_1, F_ARLEN_HBURST1(1) => 
        GND_net_1, F_ARLEN_HBURST1(0) => GND_net_1, 
        F_ARLOCK_HMASTLOCK1(1) => GND_net_1, 
        F_ARLOCK_HMASTLOCK1(0) => GND_net_1, F_ARSIZE_HSIZE1(1)
         => GND_net_1, F_ARSIZE_HSIZE1(0) => GND_net_1, 
        F_ARVALID_HWRITE1 => GND_net_1, F_AWADDR_HADDR0(31) => 
        VCC_net_1, F_AWADDR_HADDR0(30) => VCC_net_1, 
        F_AWADDR_HADDR0(29) => VCC_net_1, F_AWADDR_HADDR0(28) => 
        VCC_net_1, F_AWADDR_HADDR0(27) => VCC_net_1, 
        F_AWADDR_HADDR0(26) => VCC_net_1, F_AWADDR_HADDR0(25) => 
        VCC_net_1, F_AWADDR_HADDR0(24) => VCC_net_1, 
        F_AWADDR_HADDR0(23) => VCC_net_1, F_AWADDR_HADDR0(22) => 
        VCC_net_1, F_AWADDR_HADDR0(21) => VCC_net_1, 
        F_AWADDR_HADDR0(20) => VCC_net_1, F_AWADDR_HADDR0(19) => 
        VCC_net_1, F_AWADDR_HADDR0(18) => VCC_net_1, 
        F_AWADDR_HADDR0(17) => VCC_net_1, F_AWADDR_HADDR0(16) => 
        VCC_net_1, F_AWADDR_HADDR0(15) => VCC_net_1, 
        F_AWADDR_HADDR0(14) => VCC_net_1, F_AWADDR_HADDR0(13) => 
        VCC_net_1, F_AWADDR_HADDR0(12) => VCC_net_1, 
        F_AWADDR_HADDR0(11) => VCC_net_1, F_AWADDR_HADDR0(10) => 
        VCC_net_1, F_AWADDR_HADDR0(9) => VCC_net_1, 
        F_AWADDR_HADDR0(8) => VCC_net_1, F_AWADDR_HADDR0(7) => 
        VCC_net_1, F_AWADDR_HADDR0(6) => VCC_net_1, 
        F_AWADDR_HADDR0(5) => VCC_net_1, F_AWADDR_HADDR0(4) => 
        VCC_net_1, F_AWADDR_HADDR0(3) => VCC_net_1, 
        F_AWADDR_HADDR0(2) => VCC_net_1, F_AWADDR_HADDR0(1) => 
        VCC_net_1, F_AWADDR_HADDR0(0) => VCC_net_1, 
        F_AWBURST_HTRANS0(1) => GND_net_1, F_AWBURST_HTRANS0(0)
         => GND_net_1, F_AWID_HSEL0(3) => GND_net_1, 
        F_AWID_HSEL0(2) => GND_net_1, F_AWID_HSEL0(1) => 
        GND_net_1, F_AWID_HSEL0(0) => GND_net_1, 
        F_AWLEN_HBURST0(3) => GND_net_1, F_AWLEN_HBURST0(2) => 
        GND_net_1, F_AWLEN_HBURST0(1) => GND_net_1, 
        F_AWLEN_HBURST0(0) => GND_net_1, F_AWLOCK_HMASTLOCK0(1)
         => GND_net_1, F_AWLOCK_HMASTLOCK0(0) => GND_net_1, 
        F_AWSIZE_HSIZE0(1) => GND_net_1, F_AWSIZE_HSIZE0(0) => 
        GND_net_1, F_AWVALID_HWRITE0 => GND_net_1, F_BREADY => 
        GND_net_1, F_RMW_AXI => GND_net_1, F_RREADY => GND_net_1, 
        F_WDATA_HWDATA01(63) => VCC_net_1, F_WDATA_HWDATA01(62)
         => VCC_net_1, F_WDATA_HWDATA01(61) => VCC_net_1, 
        F_WDATA_HWDATA01(60) => VCC_net_1, F_WDATA_HWDATA01(59)
         => VCC_net_1, F_WDATA_HWDATA01(58) => VCC_net_1, 
        F_WDATA_HWDATA01(57) => VCC_net_1, F_WDATA_HWDATA01(56)
         => VCC_net_1, F_WDATA_HWDATA01(55) => VCC_net_1, 
        F_WDATA_HWDATA01(54) => VCC_net_1, F_WDATA_HWDATA01(53)
         => VCC_net_1, F_WDATA_HWDATA01(52) => VCC_net_1, 
        F_WDATA_HWDATA01(51) => VCC_net_1, F_WDATA_HWDATA01(50)
         => VCC_net_1, F_WDATA_HWDATA01(49) => VCC_net_1, 
        F_WDATA_HWDATA01(48) => VCC_net_1, F_WDATA_HWDATA01(47)
         => VCC_net_1, F_WDATA_HWDATA01(46) => VCC_net_1, 
        F_WDATA_HWDATA01(45) => VCC_net_1, F_WDATA_HWDATA01(44)
         => VCC_net_1, F_WDATA_HWDATA01(43) => VCC_net_1, 
        F_WDATA_HWDATA01(42) => VCC_net_1, F_WDATA_HWDATA01(41)
         => VCC_net_1, F_WDATA_HWDATA01(40) => VCC_net_1, 
        F_WDATA_HWDATA01(39) => VCC_net_1, F_WDATA_HWDATA01(38)
         => VCC_net_1, F_WDATA_HWDATA01(37) => VCC_net_1, 
        F_WDATA_HWDATA01(36) => VCC_net_1, F_WDATA_HWDATA01(35)
         => VCC_net_1, F_WDATA_HWDATA01(34) => VCC_net_1, 
        F_WDATA_HWDATA01(33) => VCC_net_1, F_WDATA_HWDATA01(32)
         => VCC_net_1, F_WDATA_HWDATA01(31) => VCC_net_1, 
        F_WDATA_HWDATA01(30) => VCC_net_1, F_WDATA_HWDATA01(29)
         => VCC_net_1, F_WDATA_HWDATA01(28) => VCC_net_1, 
        F_WDATA_HWDATA01(27) => VCC_net_1, F_WDATA_HWDATA01(26)
         => VCC_net_1, F_WDATA_HWDATA01(25) => VCC_net_1, 
        F_WDATA_HWDATA01(24) => VCC_net_1, F_WDATA_HWDATA01(23)
         => VCC_net_1, F_WDATA_HWDATA01(22) => VCC_net_1, 
        F_WDATA_HWDATA01(21) => VCC_net_1, F_WDATA_HWDATA01(20)
         => VCC_net_1, F_WDATA_HWDATA01(19) => VCC_net_1, 
        F_WDATA_HWDATA01(18) => VCC_net_1, F_WDATA_HWDATA01(17)
         => VCC_net_1, F_WDATA_HWDATA01(16) => VCC_net_1, 
        F_WDATA_HWDATA01(15) => VCC_net_1, F_WDATA_HWDATA01(14)
         => VCC_net_1, F_WDATA_HWDATA01(13) => VCC_net_1, 
        F_WDATA_HWDATA01(12) => VCC_net_1, F_WDATA_HWDATA01(11)
         => VCC_net_1, F_WDATA_HWDATA01(10) => VCC_net_1, 
        F_WDATA_HWDATA01(9) => VCC_net_1, F_WDATA_HWDATA01(8) => 
        VCC_net_1, F_WDATA_HWDATA01(7) => VCC_net_1, 
        F_WDATA_HWDATA01(6) => VCC_net_1, F_WDATA_HWDATA01(5) => 
        VCC_net_1, F_WDATA_HWDATA01(4) => VCC_net_1, 
        F_WDATA_HWDATA01(3) => VCC_net_1, F_WDATA_HWDATA01(2) => 
        VCC_net_1, F_WDATA_HWDATA01(1) => VCC_net_1, 
        F_WDATA_HWDATA01(0) => VCC_net_1, F_WID_HREADY01(3) => 
        GND_net_1, F_WID_HREADY01(2) => GND_net_1, 
        F_WID_HREADY01(1) => GND_net_1, F_WID_HREADY01(0) => 
        GND_net_1, F_WLAST => GND_net_1, F_WSTRB(7) => GND_net_1, 
        F_WSTRB(6) => GND_net_1, F_WSTRB(5) => GND_net_1, 
        F_WSTRB(4) => GND_net_1, F_WSTRB(3) => GND_net_1, 
        F_WSTRB(2) => GND_net_1, F_WSTRB(1) => GND_net_1, 
        F_WSTRB(0) => GND_net_1, F_WVALID => GND_net_1, 
        FPGA_MDDR_ARESET_N => VCC_net_1, MDDR_FABRIC_PADDR(10)
         => VCC_net_1, MDDR_FABRIC_PADDR(9) => VCC_net_1, 
        MDDR_FABRIC_PADDR(8) => VCC_net_1, MDDR_FABRIC_PADDR(7)
         => VCC_net_1, MDDR_FABRIC_PADDR(6) => VCC_net_1, 
        MDDR_FABRIC_PADDR(5) => VCC_net_1, MDDR_FABRIC_PADDR(4)
         => VCC_net_1, MDDR_FABRIC_PADDR(3) => VCC_net_1, 
        MDDR_FABRIC_PADDR(2) => VCC_net_1, MDDR_FABRIC_PENABLE
         => VCC_net_1, MDDR_FABRIC_PSEL => VCC_net_1, 
        MDDR_FABRIC_PWDATA(15) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(14) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(13) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(12) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(11) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(10) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(9) => VCC_net_1, MDDR_FABRIC_PWDATA(8)
         => VCC_net_1, MDDR_FABRIC_PWDATA(7) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(6) => VCC_net_1, MDDR_FABRIC_PWDATA(5)
         => VCC_net_1, MDDR_FABRIC_PWDATA(4) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(3) => VCC_net_1, MDDR_FABRIC_PWDATA(2)
         => VCC_net_1, MDDR_FABRIC_PWDATA(1) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(0) => VCC_net_1, MDDR_FABRIC_PWRITE
         => VCC_net_1, PRESET_N => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => GND_net_1, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => GND_net_1, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => GND_net_1, DM_IN(2)
         => GND_net_1, DM_IN(1) => GND_net_1, DM_IN(0) => 
        GND_net_1, DRAM_DQ_IN(17) => GND_net_1, DRAM_DQ_IN(16)
         => GND_net_1, DRAM_DQ_IN(15) => GND_net_1, 
        DRAM_DQ_IN(14) => GND_net_1, DRAM_DQ_IN(13) => GND_net_1, 
        DRAM_DQ_IN(12) => GND_net_1, DRAM_DQ_IN(11) => GND_net_1, 
        DRAM_DQ_IN(10) => GND_net_1, DRAM_DQ_IN(9) => GND_net_1, 
        DRAM_DQ_IN(8) => GND_net_1, DRAM_DQ_IN(7) => GND_net_1, 
        DRAM_DQ_IN(6) => GND_net_1, DRAM_DQ_IN(5) => GND_net_1, 
        DRAM_DQ_IN(4) => GND_net_1, DRAM_DQ_IN(3) => GND_net_1, 
        DRAM_DQ_IN(2) => GND_net_1, DRAM_DQ_IN(1) => GND_net_1, 
        DRAM_DQ_IN(0) => GND_net_1, DRAM_DQS_IN(2) => GND_net_1, 
        DRAM_DQS_IN(1) => GND_net_1, DRAM_DQS_IN(0) => GND_net_1, 
        DRAM_FIFO_WE_IN(1) => GND_net_1, DRAM_FIFO_WE_IN(0) => 
        GND_net_1, I2C0_SCL_USBC_DATA1_MGPIO31B_IN => GND_net_1, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => GND_net_1, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => GND_net_1, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => GND_net_1, MGPIO0B_IN
         => GND_net_1, MGPIO10B_IN => GND_net_1, MGPIO1B_IN => 
        GND_net_1, MGPIO25A_IN => GND_net_1, MGPIO26A_IN => 
        GND_net_1, MGPIO27A_IN => GND_net_1, MGPIO28A_IN => 
        GND_net_1, MGPIO29A_IN => GND_net_1, MGPIO2B_IN => 
        GND_net_1, MGPIO30A_IN => GND_net_1, MGPIO31A_IN => 
        GND_net_1, MGPIO3B_IN => GND_net_1, MGPIO4B_IN => 
        GND_net_1, MGPIO5B_IN => GND_net_1, MGPIO6B_IN => 
        GND_net_1, MGPIO7B_IN => GND_net_1, MGPIO8B_IN => 
        GND_net_1, MGPIO9B_IN => GND_net_1, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => GND_net_1, 
        MMUART0_DCD_MGPIO22B_IN => GND_net_1, 
        MMUART0_DSR_MGPIO20B_IN => GND_net_1, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => GND_net_1, 
        MMUART0_RI_MGPIO21B_IN => GND_net_1, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => GND_net_1, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => GND_net_1, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => GND_net_1, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => GND_net_1, 
        MMUART1_CTS_MGPIO13B_IN => GND_net_1, 
        MMUART1_DCD_MGPIO16B_IN => GND_net_1, 
        MMUART1_DSR_MGPIO14B_IN => GND_net_1, 
        MMUART1_DTR_MGPIO12B_IN => GND_net_1, 
        MMUART1_RI_MGPIO15B_IN => GND_net_1, 
        MMUART1_RTS_MGPIO11B_IN => GND_net_1, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => GND_net_1, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => GND_net_1, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => GND_net_1, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => GND_net_1, 
        RGMII_MDC_RMII_MDC_IN => GND_net_1, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => GND_net_1, 
        RGMII_RX_CLK_IN => GND_net_1, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => GND_net_1, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => GND_net_1, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => GND_net_1, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => GND_net_1, 
        RGMII_RXD3_USBB_DATA4_IN => GND_net_1, RGMII_TX_CLK_IN
         => GND_net_1, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => 
        GND_net_1, RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => GND_net_1, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => GND_net_1, 
        RGMII_TXD2_USBB_DATA5_IN => GND_net_1, 
        RGMII_TXD3_USBB_DATA6_IN => GND_net_1, 
        SPI0_SCK_USBA_XCLK_IN => GND_net_1, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => GND_net_1, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => GND_net_1, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => GND_net_1, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => GND_net_1, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => GND_net_1, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => GND_net_1, 
        SPI0_SS4_MGPIO19A_IN => GND_net_1, SPI0_SS5_MGPIO20A_IN
         => GND_net_1, SPI0_SS6_MGPIO21A_IN => GND_net_1, 
        SPI0_SS7_MGPIO22A_IN => GND_net_1, SPI1_SCK_IN => 
        GND_net_1, SPI1_SDI_MGPIO11A_IN => GND_net_1, 
        SPI1_SDO_MGPIO12A_IN => GND_net_1, SPI1_SS0_MGPIO13A_IN
         => GND_net_1, SPI1_SS1_MGPIO14A_IN => GND_net_1, 
        SPI1_SS2_MGPIO15A_IN => GND_net_1, SPI1_SS3_MGPIO16A_IN
         => GND_net_1, SPI1_SS4_MGPIO17A_IN => GND_net_1, 
        SPI1_SS5_MGPIO18A_IN => GND_net_1, SPI1_SS6_MGPIO23A_IN
         => GND_net_1, SPI1_SS7_MGPIO24A_IN => GND_net_1, 
        USBC_XCLK_IN => GND_net_1, USBD_DATA0_IN => GND_net_1, 
        USBD_DATA1_IN => GND_net_1, USBD_DATA2_IN => GND_net_1, 
        USBD_DATA3_IN => GND_net_1, USBD_DATA4_IN => GND_net_1, 
        USBD_DATA5_IN => GND_net_1, USBD_DATA6_IN => GND_net_1, 
        USBD_DATA7_MGPIO23B_IN => GND_net_1, USBD_DIR_IN => 
        GND_net_1, USBD_NXT_IN => GND_net_1, USBD_STP_IN => 
        GND_net_1, USBD_XCLK_IN => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => OPEN, DRAM_ADDR(15)
         => nc174, DRAM_ADDR(14) => nc38, DRAM_ADDR(13) => nc113, 
        DRAM_ADDR(12) => nc218, DRAM_ADDR(11) => nc106, 
        DRAM_ADDR(10) => nc261, DRAM_ADDR(9) => nc25, 
        DRAM_ADDR(8) => nc1, DRAM_ADDR(7) => nc322, DRAM_ADDR(6)
         => nc299, DRAM_ADDR(5) => nc37, DRAM_ADDR(4) => nc202, 
        DRAM_ADDR(3) => nc144, DRAM_ADDR(2) => nc153, 
        DRAM_ADDR(1) => nc46, DRAM_ADDR(0) => nc258, DRAM_BA(2)
         => nc71, DRAM_BA(1) => nc124, DRAM_BA(0) => nc332, 
        DRAM_CASN => OPEN, DRAM_CKE => OPEN, DRAM_CLK => OPEN, 
        DRAM_CSN => OPEN, DRAM_DM_RDQS_OUT(2) => nc81, 
        DRAM_DM_RDQS_OUT(1) => nc201, DRAM_DM_RDQS_OUT(0) => 
        nc168, DRAM_DQ_OUT(17) => nc323, DRAM_DQ_OUT(16) => nc34, 
        DRAM_DQ_OUT(15) => nc28, DRAM_DQ_OUT(14) => nc115, 
        DRAM_DQ_OUT(13) => nc264, DRAM_DQ_OUT(12) => nc192, 
        DRAM_DQ_OUT(11) => nc319, DRAM_DQ_OUT(10) => nc134, 
        DRAM_DQ_OUT(9) => nc32, DRAM_DQ_OUT(8) => nc40, 
        DRAM_DQ_OUT(7) => nc297, DRAM_DQ_OUT(6) => nc99, 
        DRAM_DQ_OUT(5) => nc75, DRAM_DQ_OUT(4) => nc183, 
        DRAM_DQ_OUT(3) => nc333, DRAM_DQ_OUT(2) => nc288, 
        DRAM_DQ_OUT(1) => nc85, DRAM_DQ_OUT(0) => nc27, 
        DRAM_DQS_OUT(2) => nc108, DRAM_DQS_OUT(1) => nc325, 
        DRAM_DQS_OUT(0) => nc16, DRAM_FIFO_WE_OUT(1) => nc155, 
        DRAM_FIFO_WE_OUT(0) => nc51, DRAM_ODT => OPEN, DRAM_RASN
         => OPEN, DRAM_RSTN => OPEN, DRAM_WEN => OPEN, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OUT => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => OPEN, MGPIO0B_OUT => 
        OPEN, MGPIO10B_OUT => OPEN, MGPIO1B_OUT => OPEN, 
        MGPIO25A_OUT => OPEN, MGPIO26A_OUT => OPEN, MGPIO27A_OUT
         => OPEN, MGPIO28A_OUT => OPEN, MGPIO29A_OUT => OPEN, 
        MGPIO2B_OUT => OPEN, MGPIO30A_OUT => OPEN, MGPIO31A_OUT
         => OPEN, MGPIO3B_OUT => OPEN, MGPIO4B_OUT => OPEN, 
        MGPIO5B_OUT => OPEN, MGPIO6B_OUT => OPEN, MGPIO7B_OUT => 
        OPEN, MGPIO8B_OUT => OPEN, MGPIO9B_OUT => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT => OPEN, 
        MMUART0_DCD_MGPIO22B_OUT => OPEN, 
        MMUART0_DSR_MGPIO20B_OUT => OPEN, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => OPEN, 
        MMUART1_CTS_MGPIO13B_OUT => OPEN, 
        MMUART1_DCD_MGPIO16B_OUT => OPEN, 
        MMUART1_DSR_MGPIO14B_OUT => OPEN, 
        MMUART1_DTR_MGPIO12B_OUT => OPEN, MMUART1_RI_MGPIO15B_OUT
         => OPEN, MMUART1_RTS_MGPIO11B_OUT => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => OPEN, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => OPEN, 
        RGMII_RXD3_USBB_DATA4_OUT => OPEN, RGMII_TX_CLK_OUT => 
        OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => OPEN, 
        RGMII_TXD2_USBB_DATA5_OUT => OPEN, 
        RGMII_TXD3_USBB_DATA6_OUT => OPEN, SPI0_SCK_USBA_XCLK_OUT
         => OPEN, SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => OPEN, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => OPEN, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => OPEN, 
        SPI0_SS4_MGPIO19A_OUT => OPEN, SPI0_SS5_MGPIO20A_OUT => 
        OPEN, SPI0_SS6_MGPIO21A_OUT => OPEN, 
        SPI0_SS7_MGPIO22A_OUT => OPEN, SPI1_SCK_OUT => OPEN, 
        SPI1_SDI_MGPIO11A_OUT => OPEN, SPI1_SDO_MGPIO12A_OUT => 
        OPEN, SPI1_SS0_MGPIO13A_OUT => OPEN, 
        SPI1_SS1_MGPIO14A_OUT => OPEN, SPI1_SS2_MGPIO15A_OUT => 
        OPEN, SPI1_SS3_MGPIO16A_OUT => OPEN, 
        SPI1_SS4_MGPIO17A_OUT => OPEN, SPI1_SS5_MGPIO18A_OUT => 
        OPEN, SPI1_SS6_MGPIO23A_OUT => OPEN, 
        SPI1_SS7_MGPIO24A_OUT => OPEN, USBC_XCLK_OUT => OPEN, 
        USBD_DATA0_OUT => OPEN, USBD_DATA1_OUT => OPEN, 
        USBD_DATA2_OUT => OPEN, USBD_DATA3_OUT => OPEN, 
        USBD_DATA4_OUT => OPEN, USBD_DATA5_OUT => OPEN, 
        USBD_DATA6_OUT => OPEN, USBD_DATA7_MGPIO23B_OUT => OPEN, 
        USBD_DIR_OUT => OPEN, USBD_NXT_OUT => OPEN, USBD_STP_OUT
         => OPEN, USBD_XCLK_OUT => OPEN, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => OPEN, DM_OE(2) => 
        nc301, DM_OE(1) => nc33, DM_OE(0) => nc204, 
        DRAM_DQ_OE(17) => nc173, DRAM_DQ_OE(16) => nc278, 
        DRAM_DQ_OE(15) => nc169, DRAM_DQ_OE(14) => nc78, 
        DRAM_DQ_OE(13) => nc263, DRAM_DQ_OE(12) => nc335, 
        DRAM_DQ_OE(11) => nc24, DRAM_DQ_OE(10) => nc88, 
        DRAM_DQ_OE(9) => nc111, DRAM_DQ_OE(8) => nc55, 
        DRAM_DQ_OE(7) => nc10, DRAM_DQ_OE(6) => nc22, 
        DRAM_DQ_OE(5) => nc210, DRAM_DQ_OE(4) => nc185, 
        DRAM_DQ_OE(3) => nc143, DRAM_DQ_OE(2) => nc248, 
        DRAM_DQ_OE(1) => nc77, DRAM_DQ_OE(0) => nc6, 
        DRAM_DQS_OE(2) => nc109, DRAM_DQS_OE(1) => nc87, 
        DRAM_DQS_OE(0) => nc123, I2C0_SCL_USBC_DATA1_MGPIO31B_OE
         => OPEN, I2C0_SDA_USBC_DATA0_MGPIO30B_OE => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => OPEN, MGPIO0B_OE => 
        OPEN, MGPIO10B_OE => OPEN, MGPIO1B_OE => OPEN, 
        MGPIO25A_OE => OPEN, MGPIO26A_OE => OPEN, MGPIO27A_OE => 
        OPEN, MGPIO28A_OE => OPEN, MGPIO29A_OE => OPEN, 
        MGPIO2B_OE => OPEN, MGPIO30A_OE => OPEN, MGPIO31A_OE => 
        OPEN, MGPIO3B_OE => OPEN, MGPIO4B_OE => OPEN, MGPIO5B_OE
         => OPEN, MGPIO6B_OE => OPEN, MGPIO7B_OE => OPEN, 
        MGPIO8B_OE => OPEN, MGPIO9B_OE => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => OPEN, 
        MMUART0_DCD_MGPIO22B_OE => OPEN, MMUART0_DSR_MGPIO20B_OE
         => OPEN, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => OPEN, 
        MMUART1_CTS_MGPIO13B_OE => OPEN, MMUART1_DCD_MGPIO16B_OE
         => OPEN, MMUART1_DSR_MGPIO14B_OE => OPEN, 
        MMUART1_DTR_MGPIO12B_OE => OPEN, MMUART1_RI_MGPIO15B_OE
         => OPEN, MMUART1_RTS_MGPIO11B_OE => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => OPEN, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => OPEN, 
        RGMII_RXD3_USBB_DATA4_OE => OPEN, RGMII_TX_CLK_OE => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => OPEN, 
        RGMII_TXD2_USBB_DATA5_OE => OPEN, 
        RGMII_TXD3_USBB_DATA6_OE => OPEN, SPI0_SCK_USBA_XCLK_OE
         => OPEN, SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => OPEN, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => OPEN, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => OPEN, 
        SPI0_SS4_MGPIO19A_OE => OPEN, SPI0_SS5_MGPIO20A_OE => 
        OPEN, SPI0_SS6_MGPIO21A_OE => OPEN, SPI0_SS7_MGPIO22A_OE
         => OPEN, SPI1_SCK_OE => OPEN, SPI1_SDI_MGPIO11A_OE => 
        OPEN, SPI1_SDO_MGPIO12A_OE => OPEN, SPI1_SS0_MGPIO13A_OE
         => OPEN, SPI1_SS1_MGPIO14A_OE => OPEN, 
        SPI1_SS2_MGPIO15A_OE => OPEN, SPI1_SS3_MGPIO16A_OE => 
        OPEN, SPI1_SS4_MGPIO17A_OE => OPEN, SPI1_SS5_MGPIO18A_OE
         => OPEN, SPI1_SS6_MGPIO23A_OE => OPEN, 
        SPI1_SS7_MGPIO24A_OE => OPEN, USBC_XCLK_OE => OPEN, 
        USBD_DATA0_OE => OPEN, USBD_DATA1_OE => OPEN, 
        USBD_DATA2_OE => OPEN, USBD_DATA3_OE => OPEN, 
        USBD_DATA4_OE => OPEN, USBD_DATA5_OE => OPEN, 
        USBD_DATA6_OE => OPEN, USBD_DATA7_MGPIO23B_OE => OPEN, 
        USBD_DIR_OE => OPEN, USBD_NXT_OE => OPEN, USBD_STP_OE => 
        OPEN, USBD_XCLK_OE => OPEN);
    
    MSS_ADLIB_INST_RNO_5 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1260, B => data_out_sn_N_12_mux, C => 
        N_1327, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[6]\);
    
    MSS_ADLIB_INST_RNO_25 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1280, B => data_out_sn_N_12_mux, C => 
        N_1347, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[26]\);
    
    MSS_ADLIB_INST_RNO_24 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1279, B => data_out_sn_N_12_mux, C => 
        N_1346, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[25]\);
    
    MSS_ADLIB_INST_RNO_1 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1256, B => data_out_sn_N_12_mux, C => 
        N_1323, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[2]\);
    
    MSS_ADLIB_INST_RNO_30 : CFG4
      generic map(INIT => x"F800")

      port map(A => N_1423_3, B => N_53, C => data_out_9_0_31, D
         => hready_m_xhdl339, Y => \AMBA_SLAVE_0_HRDATA_S0_m[31]\);
    
    MSS_ADLIB_INST_RNO_26 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1281, B => data_out_sn_N_12_mux, C => 
        N_1348, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[27]\);
    
    MSS_ADLIB_INST_RNO_8 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1263, B => data_out_sn_N_12_mux, C => 
        N_1330, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[9]\);
    
    MSS_ADLIB_INST_RNO_6 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1261, B => data_out_sn_N_12_mux, C => 
        N_1328, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[7]\);
    
    MSS_ADLIB_INST_RNO_28 : CFG4
      generic map(INIT => x"F080")

      port map(A => N_1446, B => N_1423_3, C => hready_m_xhdl339, 
        D => data_out_9_0_29, Y => \AMBA_SLAVE_0_HRDATA_S0_m[29]\);
    
    MSS_ADLIB_INST_RNO_9 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1264, B => data_out_sn_N_12_mux, C => 
        N_1331, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[10]\);
    
    MSS_ADLIB_INST_RNO_15 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1270, B => data_out_sn_N_12_mux, C => 
        N_1337, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[16]\);
    
    MSS_ADLIB_INST_RNO_0 : CFG4
      generic map(INIT => x"F080")

      port map(A => N_1457, B => N_1423_3, C => hready_m_xhdl339, 
        D => data_out_9_0_1, Y => \AMBA_SLAVE_0_HRDATA_S0_m[1]\);
    
    MSS_ADLIB_INST_RNO_14 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1269, B => data_out_sn_N_12_mux, C => 
        N_1336, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[15]\);
    
    MSS_ADLIB_INST_RNO_16 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1271, B => data_out_sn_N_12_mux, C => 
        N_1338, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[17]\);
    
    MSS_ADLIB_INST_RNO_18 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1273, B => data_out_sn_N_12_mux, C => 
        N_1340, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[19]\);
    
    MSS_ADLIB_INST_RNO_3 : CFG4
      generic map(INIT => x"B800")

      port map(A => N_1258, B => data_out_sn_N_12_mux, C => 
        N_1325, D => hready_m_xhdl339, Y => 
        \AMBA_SLAVE_0_HRDATA_S0_m[4]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_system_sb_FABOSC_0_OSC is

    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );

end sha256_system_sb_FABOSC_0_OSC;

architecture DEF_ARCH of sha256_system_sb_FABOSC_0_OSC is 

  component RCOSC_25_50MHZ
    generic (FREQUENCY:real := 50.0);

    port( CLKOUT : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    I_RCOSC_25_50MHZ : RCOSC_25_50MHZ
      generic map(FREQUENCY => 50.0)

      port map(CLKOUT => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreResetP is

    port( MSS_READY                                       : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK                    : in    std_logic;
          sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic;
          sha256_system_sb_0_POWER_ON_RESET_N             : in    std_logic
        );

end CoreResetP;

architecture DEF_ARCH of CoreResetP is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \MSS_HPMS_READY_int\, \mss_ready_select\, VCC_net_1, 
        \POWER_ON_RESET_N_clk_base\, 
        \un6_fic_2_apb_m_preset_n_clk_base\, GND_net_1, 
        \mss_ready_state\, \RESET_N_M2F_clk_base\, 
        \RESET_N_M2F_q1\, \FIC_2_APB_M_PRESET_N_clk_base\, 
        \FIC_2_APB_M_PRESET_N_q1\, \MSS_HPMS_READY_int_3\, 
        \POWER_ON_RESET_N_q1\ : std_logic;

begin 


    RESET_N_M2F_clk_base : SLE
      port map(D => \RESET_N_M2F_q1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RESET_N_M2F_clk_base\);
    
    POWER_ON_RESET_N_clk_base : SLE
      port map(D => \POWER_ON_RESET_N_q1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \POWER_ON_RESET_N_clk_base\);
    
    mss_ready_select : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => 
        \un6_fic_2_apb_m_preset_n_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_select\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    mss_ready_state : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => 
        \RESET_N_M2F_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_state\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    un6_fic_2_apb_m_preset_n_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \FIC_2_APB_M_PRESET_N_clk_base\, B => 
        \mss_ready_state\, Y => 
        \un6_fic_2_apb_m_preset_n_clk_base\);
    
    RESET_N_M2F_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RESET_N_M2F_q1\);
    
    FIC_2_APB_M_PRESET_N_clk_base : SLE
      port map(D => \FIC_2_APB_M_PRESET_N_q1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FIC_2_APB_M_PRESET_N_clk_base\);
    
    POWER_ON_RESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \POWER_ON_RESET_N_q1\);
    
    MSS_HPMS_READY_int_RNIFQTF : CLKINT
      port map(A => \MSS_HPMS_READY_int\, Y => MSS_READY);
    
    FIC_2_APB_M_PRESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FIC_2_APB_M_PRESET_N_q1\);
    
    MSS_HPMS_READY_int_3 : CFG3
      generic map(INIT => x"E0")

      port map(A => \RESET_N_M2F_clk_base\, B => 
        \mss_ready_select\, C => \FIC_2_APB_M_PRESET_N_clk_base\, 
        Y => \MSS_HPMS_READY_int_3\);
    
    MSS_HPMS_READY_int : SLE
      port map(D => \MSS_HPMS_READY_int_3\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \MSS_HPMS_READY_int\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVEARBITER_0 is

    port( masterAddrInProg                                   : out   std_logic_vector(3 downto 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS : in    std_logic_vector(1 to 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR  : in    std_logic_vector(27 downto 24);
          arbRegSMCurrentState_ns_i_0_0_0_a0_0               : in    std_logic_vector(1 to 1);
          SADDRSEL_0_0_0_1_0                                 : in    std_logic_vector(0 to 0);
          SADDRSEL_0_0_0_0                                   : in    std_logic_vector(0 to 0);
          HADDR_i_0                                          : in    std_logic_vector(5 downto 2);
          arbRegSMCurrentState_14                            : out   std_logic;
          arbRegSMCurrentState_13                            : out   std_logic;
          arbRegSMCurrentState_9                             : out   std_logic;
          arbRegSMCurrentState_5                             : out   std_logic;
          arbRegSMCurrentState_1                             : out   std_logic;
          MSS_READY                                          : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                       : in    std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY             : in    std_logic;
          N_321_2                                            : in    std_logic;
          N_359                                              : in    std_logic;
          N_344                                              : out   std_logic;
          N_208                                              : out   std_logic;
          d_masterRegAddrSel_0_1_i_a2_5_2_1_0                : in    std_logic;
          masterRegAddrSel                                   : in    std_logic;
          N_253                                              : in    std_logic;
          N_154_i_0                                          : out   std_logic;
          N_48_i_0                                           : out   std_logic;
          N_46_i_0                                           : out   std_logic;
          N_44_i_0                                           : out   std_logic;
          N_42_i_0                                           : out   std_logic;
          N_16_i_0                                           : out   std_logic
        );

end COREAHBLITE_SLAVEARBITER_0;

architecture DEF_ARCH of COREAHBLITE_SLAVEARBITER_0 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \arbRegSMCurrentState[1]_net_1\, VCC_net_1, N_126_i_0, 
        GND_net_1, \masterAddrInProg[3]\, N_96_i_0, 
        \arbRegSMCurrentState_14\, N_104_i_0, 
        \arbRegSMCurrentState_13\, N_106_i_0, 
        \arbRegSMCurrentState_9\, 
        \arbRegSMCurrentState_ns[5]_net_1\, 
        \arbRegSMCurrentState[9]_net_1\, N_114_i_0, 
        \masterAddrInProg[1]\, N_92_i_0, \arbRegSMCurrentState_5\, 
        \arbRegSMCurrentState_ns[9]_net_1\, 
        \arbRegSMCurrentState[5]_net_1\, N_120_i_0, 
        \masterAddrInProg[2]\, N_94_i_0, \arbRegSMCurrentState_1\, 
        \arbRegSMCurrentState_ns[13]_net_1\, N_104_i_1, \N_344\, 
        \N_208\, N_367, arbRegSMCurrentState_N_5_mux, 
        arbRegSMCurrentState_m2_0, \arbRegSMCurrentState_m2_1_0\, 
        \arbRegSMCurrentState_m2_0_0\, \HADDR_i_0_a1_0[5]\, 
        \arbRegSMCurrentState_ns_i_0_0_0_a1[1]_net_1\, 
        \arbRegSMCurrentState_ns_i_0_0_a2_c[1]\, 
        \arbRegSMCurrentState_ns_i_0_0_a2_0_1[1]_net_1\, 
        \arbRegSMCurrentState_ns_i_0_a2_1_0[0]\ : std_logic;

begin 

    masterAddrInProg(3) <= \masterAddrInProg[3]\;
    masterAddrInProg(2) <= \masterAddrInProg[2]\;
    masterAddrInProg(1) <= \masterAddrInProg[1]\;
    arbRegSMCurrentState_14 <= \arbRegSMCurrentState_14\;
    arbRegSMCurrentState_13 <= \arbRegSMCurrentState_13\;
    arbRegSMCurrentState_9 <= \arbRegSMCurrentState_9\;
    arbRegSMCurrentState_5 <= \arbRegSMCurrentState_5\;
    arbRegSMCurrentState_1 <= \arbRegSMCurrentState_1\;
    N_344 <= \N_344\;
    N_208 <= \N_208\;

    \arbRegSMCurrentState_RNO[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \masterAddrInProg[3]\, Y => N_126_i_0);
    
    \arbRegSMCurrentState_ns_i_0_0_0_a1[1]\ : CFG3
      generic map(INIT => x"45")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        N_359, C => \arbRegSMCurrentState_13\, Y => 
        \arbRegSMCurrentState_ns_i_0_0_0_a1[1]_net_1\);
    
    \arbRegSMCurrentState_ns[13]\ : CFG4
      generic map(INIT => x"ECEE")

      port map(A => arbRegSMCurrentState_m2_0, B => 
        \arbRegSMCurrentState[1]_net_1\, C => \N_208\, D => 
        \N_344\, Y => \arbRegSMCurrentState_ns[13]_net_1\);
    
    arbRegSMCurrentState_m2_0_a2 : CFG4
      generic map(INIT => x"00B0")

      port map(A => \arbRegSMCurrentState_5\, B => 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0, C => N_367, D => 
        N_359, Y => arbRegSMCurrentState_N_5_mux);
    
    \arbRegSMCurrentState_ns[9]\ : CFG4
      generic map(INIT => x"ECEE")

      port map(A => \arbRegSMCurrentState_m2_0_0\, B => 
        \arbRegSMCurrentState[5]_net_1\, C => \N_208\, D => 
        \N_344\, Y => \arbRegSMCurrentState_ns[9]_net_1\);
    
    \arbRegSMCurrentState[8]\ : SLE
      port map(D => N_92_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \masterAddrInProg[1]\);
    
    \arbRegSMCurrentState[10]\ : SLE
      port map(D => \arbRegSMCurrentState_ns[5]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_9\);
    
    \arbRegSMCurrentState_RNO_0[15]\ : CFG3
      generic map(INIT => x"51")

      port map(A => N_359, B => \N_344\, C => \N_208\, Y => 
        N_104_i_1);
    
    \arbRegSMCurrentState_RNINANK2[15]\ : CFG4
      generic map(INIT => x"3331")

      port map(A => \N_208\, B => 
        \arbRegSMCurrentState_ns_i_0_a2_1_0[0]\, C => 
        \arbRegSMCurrentState_14\, D => N_359, Y => N_16_i_0);
    
    \arbRegSMCurrentState_ns_a2_0_i_0_o2_RNI62N62[5]\ : CFG4
      generic map(INIT => x"1131")

      port map(A => \HADDR_i_0_a1_0[5]\, B => HADDR_i_0(5), C => 
        \N_344\, D => \N_208\, Y => N_48_i_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \arbRegSMCurrentState_RNO[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \masterAddrInProg[3]\, Y => N_96_i_0);
    
    \arbRegSMCurrentState_ns_a2_0_i_0_o2_RNI51N62[5]\ : CFG4
      generic map(INIT => x"1131")

      port map(A => \HADDR_i_0_a1_0[5]\, B => HADDR_i_0(4), C => 
        \N_344\, D => \N_208\, Y => N_46_i_0);
    
    \arbRegSMCurrentState[0]\ : SLE
      port map(D => N_96_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \masterAddrInProg[3]\);
    
    arbRegSMCurrentState_m2_1_0 : CFG2
      generic map(INIT => x"4")

      port map(A => N_359, B => \arbRegSMCurrentState_9\, Y => 
        \arbRegSMCurrentState_m2_1_0\);
    
    \arbRegSMCurrentState_RNO[15]\ : CFG4
      generic map(INIT => x"2223")

      port map(A => \arbRegSMCurrentState_14\, B => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, C => N_321_2, D
         => N_104_i_1, Y => N_104_i_0);
    
    \arbRegSMCurrentState_ns_i_0_0_a2_0_1[1]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => arbRegSMCurrentState_ns_i_0_0_0_a0_0(1), B
         => \arbRegSMCurrentState_ns_i_0_0_0_a1[1]_net_1\, C => 
        \N_208\, D => \arbRegSMCurrentState_ns_i_0_0_a2_c[1]\, Y
         => \arbRegSMCurrentState_ns_i_0_0_a2_0_1[1]_net_1\);
    
    \arbRegSMCurrentState_ns_a2_0_i_0_a2_1_RNIMG872[5]\ : CFG4
      generic map(INIT => x"8FCF")

      port map(A => N_321_2, B => SADDRSEL_0_0_0_1_0(0), C => 
        N_253, D => \N_344\, Y => 
        \arbRegSMCurrentState_ns_i_0_a2_1_0[0]\);
    
    \arbRegSMCurrentState_RNO[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \masterAddrInProg[1]\, Y => N_92_i_0);
    
    \arbRegSMCurrentState[14]\ : SLE
      port map(D => N_106_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_13\);
    
    arbRegSMCurrentState_m2_0_0 : CFG2
      generic map(INIT => x"4")

      port map(A => N_359, B => \arbRegSMCurrentState_5\, Y => 
        \arbRegSMCurrentState_m2_0_0\);
    
    \arbRegSMCurrentState[6]\ : SLE
      port map(D => \arbRegSMCurrentState_ns[9]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_5\);
    
    \arbRegSMCurrentState[1]\ : SLE
      port map(D => N_126_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[1]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \arbRegSMCurrentState_RNO[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \masterAddrInProg[2]\, Y => N_94_i_0);
    
    \arbRegSMCurrentState_ns_i_0_0_a2_c_0[1]\ : CFG4
      generic map(INIT => x"CFAA")

      port map(A => N_321_2, B => masterRegAddrSel, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), D
         => arbRegSMCurrentState_N_5_mux, Y => 
        \arbRegSMCurrentState_ns_i_0_0_a2_c[1]\);
    
    \arbRegSMCurrentState_RNO[14]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \N_208\, B => 
        \arbRegSMCurrentState_ns_i_0_0_a2_0_1[1]_net_1\, C => 
        N_367, D => N_359, Y => N_106_i_0);
    
    \arbRegSMCurrentState[9]\ : SLE
      port map(D => N_114_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[9]_net_1\);
    
    \arbRegSMCurrentState[4]\ : SLE
      port map(D => N_94_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \masterAddrInProg[2]\);
    
    \arbRegSMCurrentState_RNIAT3S1[15]\ : CFG4
      generic map(INIT => x"AEAF")

      port map(A => \arbRegSMCurrentState_14\, B => N_359, C => 
        SADDRSEL_0_0_0_0(0), D => \N_208\, Y => N_154_i_0);
    
    arbRegSMCurrentState_m2_0_1 : CFG2
      generic map(INIT => x"4")

      port map(A => N_359, B => \arbRegSMCurrentState_1\, Y => 
        arbRegSMCurrentState_m2_0);
    
    \arbRegSMCurrentState_ns_a2_0_i_0_a2_1[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), B
         => masterRegAddrSel, Y => \N_344\);
    
    \arbRegSMCurrentState[2]\ : SLE
      port map(D => \arbRegSMCurrentState_ns[13]_net_1\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_1\);
    
    \arbRegSMCurrentState_ns_a2_0_i_0_o2_RNI3VM62[5]\ : CFG4
      generic map(INIT => x"1131")

      port map(A => \HADDR_i_0_a1_0[5]\, B => HADDR_i_0(2), C => 
        \N_344\, D => \N_208\, Y => N_42_i_0);
    
    \arbRegSMCurrentState[5]\ : SLE
      port map(D => N_120_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[5]_net_1\);
    
    \arbRegSMCurrentState[15]\ : SLE
      port map(D => N_104_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => VCC_net_1, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_14\);
    
    \arbRegSMCurrentState_RNI54F8[15]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_359, B => \arbRegSMCurrentState_14\, Y => 
        \HADDR_i_0_a1_0[5]\);
    
    \arbRegSMCurrentState_ns_i_0_0_a2_1[1]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \arbRegSMCurrentState_14\, B => 
        \arbRegSMCurrentState_13\, Y => N_367);
    
    \arbRegSMCurrentState_ns[5]\ : CFG4
      generic map(INIT => x"ECEE")

      port map(A => \arbRegSMCurrentState_m2_1_0\, B => 
        \arbRegSMCurrentState[9]_net_1\, C => \N_208\, D => 
        \N_344\, Y => \arbRegSMCurrentState_ns[5]_net_1\);
    
    \arbRegSMCurrentState_RNO[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \masterAddrInProg[2]\, Y => N_120_i_0);
    
    \arbRegSMCurrentState_ns_a2_0_i_0_o2[5]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(26), B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(24), 
        C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(27), D
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(25), 
        Y => \N_208\);
    
    \arbRegSMCurrentState_ns_a2_0_i_0_o2_RNI40N62[5]\ : CFG4
      generic map(INIT => x"1131")

      port map(A => \HADDR_i_0_a1_0[5]\, B => HADDR_i_0(3), C => 
        \N_344\, D => \N_208\, Y => N_44_i_0);
    
    \arbRegSMCurrentState_RNO[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \masterAddrInProg[1]\, Y => N_114_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVESTAGE_1 is

    port( masterAddrInProg                                     : out   std_logic_vector(3 downto 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0);
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          regHADDR                                             : in    std_logic_vector(5 downto 2);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1);
          arbRegSMCurrentState_ns_i_0_0_0_a0_0                 : in    std_logic_vector(1 to 1);
          SADDRSEL_0_0_0_1_0                                   : in    std_logic_vector(0 to 0);
          SADDRSEL_0_0_0_0                                     : in    std_logic_vector(0 to 0);
          masterDataInProg_0                                   : out   std_logic;
          arbRegSMCurrentState_13                              : out   std_logic;
          arbRegSMCurrentState_12                              : out   std_logic;
          arbRegSMCurrentState_8                               : out   std_logic;
          arbRegSMCurrentState_4                               : out   std_logic;
          arbRegSMCurrentState_0                               : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic;
          MSS_READY                                            : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic;
          N_321_2                                              : in    std_logic;
          masterRegAddrSel                                     : in    std_logic;
          N_359                                                : in    std_logic;
          N_344                                                : out   std_logic;
          N_208                                                : out   std_logic;
          d_masterRegAddrSel_0_1_i_a2_5_2_1_0                  : in    std_logic;
          N_253                                                : in    std_logic;
          N_48_i_0                                             : out   std_logic;
          N_46_i_0                                             : out   std_logic;
          N_44_i_0                                             : out   std_logic;
          N_42_i_0                                             : out   std_logic;
          N_16_i_0                                             : out   std_logic
        );

end COREAHBLITE_SLAVESTAGE_1;

architecture DEF_ARCH of COREAHBLITE_SLAVESTAGE_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVEARBITER_0
    port( masterAddrInProg                                   : out   std_logic_vector(3 downto 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS : in    std_logic_vector(1 to 1) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR  : in    std_logic_vector(27 downto 24) := (others => 'U');
          arbRegSMCurrentState_ns_i_0_0_0_a0_0               : in    std_logic_vector(1 to 1) := (others => 'U');
          SADDRSEL_0_0_0_1_0                                 : in    std_logic_vector(0 to 0) := (others => 'U');
          SADDRSEL_0_0_0_0                                   : in    std_logic_vector(0 to 0) := (others => 'U');
          HADDR_i_0                                          : in    std_logic_vector(5 downto 2) := (others => 'U');
          arbRegSMCurrentState_14                            : out   std_logic;
          arbRegSMCurrentState_13                            : out   std_logic;
          arbRegSMCurrentState_9                             : out   std_logic;
          arbRegSMCurrentState_5                             : out   std_logic;
          arbRegSMCurrentState_1                             : out   std_logic;
          MSS_READY                                          : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                       : in    std_logic := 'U';
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY             : in    std_logic := 'U';
          N_321_2                                            : in    std_logic := 'U';
          N_359                                              : in    std_logic := 'U';
          N_344                                              : out   std_logic;
          N_208                                              : out   std_logic;
          d_masterRegAddrSel_0_1_i_a2_5_2_1_0                : in    std_logic := 'U';
          masterRegAddrSel                                   : in    std_logic := 'U';
          N_253                                              : in    std_logic := 'U';
          N_154_i_0                                          : out   std_logic;
          N_48_i_0                                           : out   std_logic;
          N_46_i_0                                           : out   std_logic;
          N_44_i_0                                           : out   std_logic;
          N_42_i_0                                           : out   std_logic;
          N_16_i_0                                           : out   std_logic
        );
  end component;

    signal \masterDataInProg[3]_net_1\, VCC_net_1, 
        \masterAddrInProg[3]\, GND_net_1, \masterDataInProg_0\, 
        N_154_i_0, \masterDataInProg[1]_net_1\, 
        \masterAddrInProg[1]\, \masterDataInProg[2]_net_1\, 
        \masterAddrInProg[2]\, \hwdata10\, \HADDR_i_0[5]_net_1\, 
        \HADDR_i_0[3]_net_1\, \HADDR_i_0[2]_net_1\, 
        \HADDR_i_0[4]_net_1\ : std_logic;

    for all : COREAHBLITE_SLAVEARBITER_0
	Use entity work.COREAHBLITE_SLAVEARBITER_0(DEF_ARCH);
begin 

    masterAddrInProg(3) <= \masterAddrInProg[3]\;
    masterAddrInProg(2) <= \masterAddrInProg[2]\;
    masterAddrInProg(1) <= \masterAddrInProg[1]\;
    masterDataInProg_0 <= \masterDataInProg_0\;

    \masterDataInProg[3]\ : SLE
      port map(D => \masterAddrInProg[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \masterDataInProg[3]_net_1\);
    
    hwdata10_RNI2UPH_18 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(22));
    
    hwdata10_RNI2UPH_20 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(20));
    
    hwdata10_RNI2UPH_11 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(29));
    
    hwdata10_RNI2UPH_22 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(18));
    
    hwdata10_RNI2UPH_23 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(17));
    
    hwdata10_RNI2UPH_0 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(8));
    
    hwdata10_RNI2UPH_10 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(30));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \masterDataInProg[2]\ : SLE
      port map(D => \masterAddrInProg[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \masterDataInProg[2]_net_1\);
    
    hwdata10_RNI2UPH_26 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(14));
    
    hwdata10_RNI2UPH_12 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(28));
    
    hwdata10_RNI2UPH_3 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(5));
    
    \HADDR_i_0[4]\ : CFG4
      generic map(INIT => x"AFBB")

      port map(A => N_321_2, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, C
         => regHADDR(4), D => masterRegAddrSel, Y => 
        \HADDR_i_0[4]_net_1\);
    
    hwdata10_RNI2UPH_13 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(27));
    
    hwdata10_RNI2UPH_5 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(3));
    
    hwdata10_RNI2UPH_25 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(15));
    
    hwdata10_RNI2UPH_24 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(16));
    
    hwdata10_RNI2UPH_16 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(24));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \HADDR_i_0[2]\ : CFG4
      generic map(INIT => x"AFBB")

      port map(A => N_321_2, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, C
         => regHADDR(2), D => masterRegAddrSel, Y => 
        \HADDR_i_0[2]_net_1\);
    
    \masterDataInProg[1]\ : SLE
      port map(D => \masterAddrInProg[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \masterDataInProg[1]_net_1\);
    
    \masterDataInProg[0]\ : SLE
      port map(D => N_154_i_0, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \masterDataInProg_0\);
    
    hwdata10_RNI2UPH_2 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(6));
    
    hwdata10_RNI2UPH_29 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(11));
    
    \HADDR_i_0[3]\ : CFG4
      generic map(INIT => x"AFBB")

      port map(A => N_321_2, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, C
         => regHADDR(3), D => masterRegAddrSel, Y => 
        \HADDR_i_0[3]_net_1\);
    
    hwdata10_RNI2UPH_15 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(25));
    
    hwdata10_RNI2UPH_14 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(26));
    
    hwdata10_RNI2UPH_8 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(0));
    
    hwdata10_RNI2UPH_7 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(1));
    
    hwdata10_RNI2UPH_1 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(7));
    
    hwdata10_RNI2UPH_27 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(13));
    
    hwdata10_RNI2UPH_19 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(21));
    
    slave_arbiter : COREAHBLITE_SLAVEARBITER_0
      port map(masterAddrInProg(3) => \masterAddrInProg[3]\, 
        masterAddrInProg(2) => \masterAddrInProg[2]\, 
        masterAddrInProg(1) => \masterAddrInProg[1]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(27) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(26) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(25) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(24) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1) => 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1), 
        SADDRSEL_0_0_0_1_0(0) => SADDRSEL_0_0_0_1_0(0), 
        SADDRSEL_0_0_0_0(0) => SADDRSEL_0_0_0_0(0), HADDR_i_0(5)
         => \HADDR_i_0[5]_net_1\, HADDR_i_0(4) => 
        \HADDR_i_0[4]_net_1\, HADDR_i_0(3) => 
        \HADDR_i_0[3]_net_1\, HADDR_i_0(2) => 
        \HADDR_i_0[2]_net_1\, arbRegSMCurrentState_14 => 
        arbRegSMCurrentState_13, arbRegSMCurrentState_13 => 
        arbRegSMCurrentState_12, arbRegSMCurrentState_9 => 
        arbRegSMCurrentState_8, arbRegSMCurrentState_5 => 
        arbRegSMCurrentState_4, arbRegSMCurrentState_1 => 
        arbRegSMCurrentState_0, MSS_READY => MSS_READY, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, N_321_2 => 
        N_321_2, N_359 => N_359, N_344 => N_344, N_208 => N_208, 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0 => 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0, masterRegAddrSel => 
        masterRegAddrSel, N_253 => N_253, N_154_i_0 => N_154_i_0, 
        N_48_i_0 => N_48_i_0, N_46_i_0 => N_46_i_0, N_44_i_0 => 
        N_44_i_0, N_42_i_0 => N_42_i_0, N_16_i_0 => N_16_i_0);
    
    hwdata10 : CFG4
      generic map(INIT => x"0100")

      port map(A => \masterDataInProg[3]_net_1\, B => 
        \masterDataInProg[2]_net_1\, C => 
        \masterDataInProg[1]_net_1\, D => \masterDataInProg_0\, Y
         => \hwdata10\);
    
    hwdata10_RNI2UPH_17 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(23));
    
    hwdata10_RNI2UPH_4 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(4));
    
    \HADDR_i_0[5]\ : CFG4
      generic map(INIT => x"AFBB")

      port map(A => N_321_2, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, C
         => regHADDR(5), D => masterRegAddrSel, Y => 
        \HADDR_i_0[5]_net_1\);
    
    hwdata10_RNI2UPH_28 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(12));
    
    hwdata10_RNI2UPH_30 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(10));
    
    hwdata10_RNI2UPH_21 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(19));
    
    hwdata10_RNI2UPH_6 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(2));
    
    hwdata10_RNI2UPH_9 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(31));
    
    hwdata10_RNI2UPH : CFG2
      generic map(INIT => x"8")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), B
         => \hwdata10\, Y => AHB_slave_dummy_0_mem_wdata(9));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_DEFAULTSLAVESM_0 is

    port( xhdl1222                     : in    std_logic_vector(0 to 0);
          SDATASELInt_12               : in    std_logic;
          SDATASELInt_1                : in    std_logic;
          SDATASELInt_10               : in    std_logic;
          SDATASELInt_5                : in    std_logic;
          SDATASELInt_4                : in    std_logic;
          SDATASELInt_3                : in    std_logic;
          SDATASELInt_2                : in    std_logic;
          SDATASELInt_14               : in    std_logic;
          SDATASELInt_13               : in    std_logic;
          SDATASELInt_8                : in    std_logic;
          SDATASELInt_0                : in    std_logic;
          defSlaveSMCurrentState       : out   std_logic;
          MSS_READY                    : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK : in    std_logic;
          N_357                        : out   std_logic;
          HREADY_M_iv_i_i_1_1          : in    std_logic;
          N_358                        : out   std_logic;
          N_453_tz                     : in    std_logic;
          HREADY_M_iv_i_i_1            : out   std_logic;
          N_356                        : out   std_logic;
          N_353                        : out   std_logic;
          N_352                        : out   std_logic;
          N_354                        : in    std_logic;
          N_355                        : out   std_logic
        );

end COREAHBLITE_DEFAULTSLAVESM_0;

architecture DEF_ARCH of COREAHBLITE_DEFAULTSLAVESM_0 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal defSlaveSMCurrentState_net_1, VCC_net_1, N_38_i_0, 
        GND_net_1, \N_357\, \N_358\, \N_353\, \N_352\, \N_355\
         : std_logic;

begin 

    defSlaveSMCurrentState <= defSlaveSMCurrentState_net_1;
    N_357 <= \N_357\;
    N_358 <= \N_358\;
    N_353 <= \N_353\;
    N_352 <= \N_352\;
    N_355 <= \N_355\;

    defSlaveSMNextState_i_a2_4 : CFG3
      generic map(INIT => x"01")

      port map(A => SDATASELInt_12, B => SDATASELInt_1, C => 
        SDATASELInt_10, Y => N_356);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    defSlaveSMNextState_i_a2_3 : CFG4
      generic map(INIT => x"0001")

      port map(A => SDATASELInt_5, B => SDATASELInt_4, C => 
        SDATASELInt_3, D => SDATASELInt_2, Y => \N_353\);
    
    defSlaveSMCurrentState_RNO : CFG3
      generic map(INIT => x"13")

      port map(A => \N_357\, B => defSlaveSMCurrentState_net_1, C
         => \N_355\, Y => N_38_i_0);
    
    \defSlaveSMCurrentState\ : SLE
      port map(D => N_38_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        defSlaveSMCurrentState_net_1);
    
    defSlaveSMCurrentState_RNIU1EG : CFG2
      generic map(INIT => x"1")

      port map(A => xhdl1222(0), B => 
        defSlaveSMCurrentState_net_1, Y => \N_358\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    defSlaveSMNextState_i_a2_1_RNICKFE1 : CFG4
      generic map(INIT => x"B030")

      port map(A => \N_357\, B => HREADY_M_iv_i_i_1_1, C => 
        \N_358\, D => N_453_tz, Y => HREADY_M_iv_i_i_1);
    
    defSlaveSMNextState_i_a2_2 : CFG4
      generic map(INIT => x"0001")

      port map(A => SDATASELInt_14, B => SDATASELInt_13, C => 
        SDATASELInt_8, D => SDATASELInt_0, Y => \N_352\);
    
    defSlaveSMNextState_i_a2_0 : CFG2
      generic map(INIT => x"8")

      port map(A => \N_352\, B => \N_353\, Y => \N_355\);
    
    defSlaveSMNextState_i_a2_1 : CFG4
      generic map(INIT => x"0010")

      port map(A => SDATASELInt_12, B => SDATASELInt_10, C => 
        N_354, D => SDATASELInt_1, Y => \N_357\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MASTERSTAGE_2_1_0_1_0 is

    port( regHADDR                                             : out   std_logic_vector(5 downto 2);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1);
          masterDataInProg                                     : in    std_logic_vector(0 to 0);
          SADDRSEL_0_0_0_0                                     : out   std_logic_vector(0 to 0);
          SADDRSEL_0_0_0_1_0                                   : out   std_logic_vector(0 to 0);
          arbRegSMCurrentState_ns_i_0_0_0_a0_0                 : in    std_logic_vector(1 to 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          arbRegSMCurrentState_0                               : in    std_logic;
          arbRegSMCurrentState_8                               : in    std_logic;
          arbRegSMCurrentState_13                              : in    std_logic;
          arbRegSMCurrentState_12                              : in    std_logic;
          arbRegSMCurrentState_4                               : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic;
          MSS_READY                                            : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic;
          regHWRITE                                            : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic;
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_358                                                : out   std_logic;
          N_401                                                : out   std_logic;
          N_403                                                : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic;
          N_208                                                : in    std_logic;
          N_211                                                : out   std_logic;
          N_354                                                : out   std_logic;
          N_355                                                : out   std_logic;
          N_395                                                : out   std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          N_23_i_0                                             : out   std_logic;
          d_masterRegAddrSel_0_1_i_a2_5_2_1_0                  : out   std_logic;
          N_359                                                : out   std_logic;
          N_253                                                : out   std_logic;
          N_344                                                : in    std_logic;
          N_321_2                                              : out   std_logic;
          N_36_2                                               : in    std_logic
        );

end COREAHBLITE_MASTERSTAGE_2_1_0_1_0;

architecture DEF_ARCH of COREAHBLITE_MASTERSTAGE_2_1_0_1_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_DEFAULTSLAVESM_0
    port( xhdl1222                     : in    std_logic_vector(0 to 0) := (others => 'U');
          SDATASELInt_12               : in    std_logic := 'U';
          SDATASELInt_1                : in    std_logic := 'U';
          SDATASELInt_10               : in    std_logic := 'U';
          SDATASELInt_5                : in    std_logic := 'U';
          SDATASELInt_4                : in    std_logic := 'U';
          SDATASELInt_3                : in    std_logic := 'U';
          SDATASELInt_2                : in    std_logic := 'U';
          SDATASELInt_14               : in    std_logic := 'U';
          SDATASELInt_13               : in    std_logic := 'U';
          SDATASELInt_8                : in    std_logic := 'U';
          SDATASELInt_0                : in    std_logic := 'U';
          defSlaveSMCurrentState       : out   std_logic;
          MSS_READY                    : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK : in    std_logic := 'U';
          N_357                        : out   std_logic;
          HREADY_M_iv_i_i_1_1          : in    std_logic := 'U';
          N_358                        : out   std_logic;
          N_453_tz                     : in    std_logic := 'U';
          HREADY_M_iv_i_i_1            : out   std_logic;
          N_356                        : out   std_logic;
          N_353                        : out   std_logic;
          N_352                        : out   std_logic;
          N_354                        : in    std_logic := 'U';
          N_355                        : out   std_logic
        );
  end component;

    signal \SDATASELInt[1]_net_1\, VCC_net_1, \SADDRSEL[1]\, 
        N_21_i_0, GND_net_1, \SDATASELInt[2]_net_1\, 
        \SADDRSEL[2]\, \SDATASELInt[3]_net_1\, \SADDRSEL[3]\, 
        \SDATASELInt[4]_net_1\, \SADDRSEL[4]\, 
        \SDATASELInt[5]_net_1\, \SADDRSEL[5]\, 
        \SDATASELInt[6]_net_1\, \SADDRSEL[6]\, 
        \SDATASELInt[7]_net_1\, \SADDRSEL[7]\, 
        \SDATASELInt[8]_net_1\, \SADDRSEL[8]\, 
        \SDATASELInt[9]_net_1\, \SADDRSEL[9]\, 
        \SDATASELInt[10]_net_1\, \SADDRSEL[10]\, 
        \SDATASELInt[11]_net_1\, \SADDRSEL[11]\, 
        \SDATASELInt[12]_net_1\, \SADDRSEL[12]\, 
        \SDATASELInt[13]_net_1\, \SADDRSEL[13]\, 
        \SDATASELInt[14]_net_1\, \SADDRSEL[14]\, 
        \SDATASELInt[15]_net_1\, N_296, N_36_i_0, \xhdl1222[0]\, 
        \xhdl1221[0]\, regHWRITE_net_1, regHTRANS_net_1, 
        masterRegAddrSel_net_1, N_30_i_0, N_353, N_203, N_357, 
        \N_358\, \N_401\, N_352, N_202, \N_403\, N_36_i_1, 
        d_masterRegAddrSel_0_1_i_a2_5_out, 
        \d_masterRegAddrSel_0_1_i_2_0\, 
        \d_masterRegAddrSel_0_1_i_2_1\, \N_211\, \N_354\, \N_355\, 
        \N_395\, HREADY_M_iv_i_i_1_1, HREADY_M_iv_i_i_1, 
        \hready_m_xhdl339\, N_340, N_210, 
        \SADDRSEL_0_a2_0_a2_0_0[7]_net_1\, 
        \d_masterRegAddrSel_0_i_a2_0_0\, 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0_net_1, \N_359\, N_394, 
        N_360, \N_321_2\, N_189, defSlaveSMCurrentState, N_235, 
        \d_masterRegAddrSel_0_i_a0_1\, N_356, 
        \d_masterRegAddrSel_0_1_i_o2_0_0_d\, 
        \d_masterRegAddrSel_0_1_i_o2_0_0_c\, 
        \d_masterRegAddrSel_0_i_o2_0\, N_453_tz, N_397, N_281, 
        N_299, N_286, \d_masterRegAddrSel_0_i_3_0\, 
        \un1_hready_m_xhdl339_2_i_0_0_o2_0\, 
        \d_masterRegAddrSel_0_i_1_tz\, N_159, 
        \d_masterRegAddrSel_0_i_3_2\ : std_logic;

    for all : COREAHBLITE_DEFAULTSLAVESM_0
	Use entity work.COREAHBLITE_DEFAULTSLAVESM_0(DEF_ARCH);
begin 

    regHWRITE <= regHWRITE_net_1;
    regHTRANS <= regHTRANS_net_1;
    masterRegAddrSel <= masterRegAddrSel_net_1;
    N_358 <= \N_358\;
    N_401 <= \N_401\;
    N_403 <= \N_403\;
    N_211 <= \N_211\;
    N_354 <= \N_354\;
    N_355 <= \N_355\;
    N_395 <= \N_395\;
    hready_m_xhdl339 <= \hready_m_xhdl339\;
    d_masterRegAddrSel_0_1_i_a2_5_2_1_0 <= 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0_net_1;
    N_359 <= \N_359\;
    N_321_2 <= \N_321_2\;

    d_masterRegAddrSel_0_1_i_o2_2_RNI3IPJ : CFG4
      generic map(INIT => x"8000")

      port map(A => N_352, B => N_202, C => N_357, D => \N_358\, 
        Y => \N_403\);
    
    \SADDRSEL_0_a2_0_a2[2]\ : CFG3
      generic map(INIT => x"08")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, B
         => N_394, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, Y
         => \SADDRSEL[2]\);
    
    d_masterRegAddrSel_0_i_o2_2 : CFG4
      generic map(INIT => x"CFCE")

      port map(A => arbRegSMCurrentState_ns_i_0_0_0_a0_0(1), B
         => \d_masterRegAddrSel_0_i_o2_0\, C => N_208, D => 
        d_masterRegAddrSel_0_1_i_a2_5_out, Y => N_159);
    
    d_masterRegAddrSel_0_1_i_o2_3_RNI5IPJ : CFG4
      generic map(INIT => x"8000")

      port map(A => N_353, B => N_203, C => N_357, D => \N_358\, 
        Y => \N_401\);
    
    \SADDRSEL_0_a2_0_a2[6]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => N_344, D => \SADDRSEL_0_a2_0_a2_0_0[7]_net_1\, Y => 
        \SADDRSEL[6]\);
    
    d_masterRegAddrSel_0_i_o2_0 : CFG4
      generic map(INIT => x"FF60")

      port map(A => \SDATASELInt[13]_net_1\, B => 
        \SDATASELInt[2]_net_1\, C => \N_358\, D => N_340, Y => 
        N_210);
    
    d_masterRegAddrSel_0_i_a2_6 : CFG4
      generic map(INIT => x"0010")

      port map(A => \SDATASELInt[2]_net_1\, B => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, C => 
        \xhdl1222[0]\, D => \SDATASELInt[13]_net_1\, Y => N_340);
    
    \SADDRSEL_0_a2_0_a2[14]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        D => N_360, Y => \SADDRSEL[14]\);
    
    d_masterRegAddrSel_0_i_o2_1 : CFG4
      generic map(INIT => x"0246")

      port map(A => \xhdl1222[0]\, B => \SDATASELInt[11]_net_1\, 
        C => masterDataInProg(0), D => defSlaveSMCurrentState, Y
         => N_235);
    
    un1_hready_m_xhdl339_2_i_0_0_a2_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => \N_211\, B => \N_354\, C => N_353, D => N_352, 
        Y => N_397);
    
    d_masterRegAddrSel_0_1_i_o2_0_0_c : CFG4
      generic map(INIT => x"222F")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \N_321_2\, C => \SDATASELInt[13]_net_1\, D => 
        \SDATASELInt[2]_net_1\, Y => 
        \d_masterRegAddrSel_0_1_i_o2_0_0_c\);
    
    d_masterRegAddrSel_0_1_i_a2_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => \SDATASELInt[11]_net_1\, B => \N_354\, C => 
        \N_355\, D => N_210, Y => N_286);
    
    \masterRegAddrSel\ : SLE
      port map(D => N_30_i_0, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        masterRegAddrSel_net_1);
    
    \SADDRSEL_0_0_a2_1[15]\ : CFG2
      generic map(INIT => x"8")

      port map(A => masterRegAddrSel_net_1, B => regHTRANS_net_1, 
        Y => \N_359\);
    
    \regHTRANS\ : SLE
      port map(D => VCC_net_1, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_36_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHTRANS_net_1);
    
    hready_m_xhdl339_0_a5_0_a2_RNIM4RH2 : CFG4
      generic map(INIT => x"080F")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        masterDataInProg(0), C => HREADY_M_iv_i_i_1, D => 
        \hready_m_xhdl339\, Y => N_23_i_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \SADDRSEL_0_a2_2_a2[9]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        D => N_360, Y => \SADDRSEL[9]\);
    
    \SADDRSEL_0_a2_1_a2[11]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        D => N_360, Y => \SADDRSEL[11]\);
    
    d_masterRegAddrSel_0_1_i_2_1 : CFG4
      generic map(INIT => x"ECCC")

      port map(A => \d_masterRegAddrSel_0_1_i_o2_0_0_d\, B => 
        N_36_2, C => N_235, D => 
        \d_masterRegAddrSel_0_1_i_o2_0_0_c\, Y => 
        \d_masterRegAddrSel_0_1_i_2_1\);
    
    d_masterRegAddrSel_0_i_a2_13 : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt[12]_net_1\, B => 
        \SDATASELInt[10]_net_1\, C => \SDATASELInt[8]_net_1\, D
         => \SDATASELInt[7]_net_1\, Y => \N_354\);
    
    d_masterRegAddrSel_0_i_1_tz : CFG3
      generic map(INIT => x"F8")

      port map(A => \N_358\, B => \N_395\, C => \N_403\, Y => 
        \d_masterRegAddrSel_0_i_1_tz\);
    
    \SADDRSEL_0_a2_2_a2[8]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        D => N_360, Y => \SADDRSEL[8]\);
    
    d_masterRegAddrSel_0_i_o2_0_0 : CFG3
      generic map(INIT => x"C4")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        \N_359\, C => \N_321_2\, Y => 
        \d_masterRegAddrSel_0_i_o2_0\);
    
    \d_masterRegAddrSel_0_1_i_a2_5_2_1_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => arbRegSMCurrentState_0, B => 
        arbRegSMCurrentState_8, Y => 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0_net_1);
    
    un1_hready_m_xhdl339_2_i_0_0_o2_0_RNI23MO : CFG4
      generic map(INIT => x"007F")

      port map(A => \N_211\, B => \N_354\, C => \N_355\, D => 
        \N_395\, Y => HREADY_M_iv_i_i_1_1);
    
    d_masterRegAddrSel_0_1_i_o2_3 : CFG4
      generic map(INIT => x"0116")

      port map(A => \SDATASELInt[15]_net_1\, B => 
        \SDATASELInt[14]_net_1\, C => \SDATASELInt[9]_net_1\, D
         => \SDATASELInt[1]_net_1\, Y => N_203);
    
    \regHADDR[5]\ : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => N_36_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(5));
    
    \SDATASELInt[4]\ : SLE
      port map(D => \SADDRSEL[4]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[4]_net_1\);
    
    \regHADDR[2]\ : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => N_36_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(2));
    
    d_masterRegAddrSel_0_1_i_a2_5_s : CFG3
      generic map(INIT => x"08")

      port map(A => \N_321_2\, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), C
         => masterRegAddrSel_net_1, Y => 
        d_masterRegAddrSel_0_1_i_a2_5_out);
    
    \SDATASELInt[15]\ : SLE
      port map(D => N_296, CLK => sha256_system_sb_0_FIC_0_CLK, 
        EN => N_21_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[15]_net_1\);
    
    d_masterRegAddrSel_0_1_i_o2_2 : CFG4
      generic map(INIT => x"0116")

      port map(A => \SDATASELInt[6]_net_1\, B => 
        \SDATASELInt[5]_net_1\, C => \SDATASELInt[4]_net_1\, D
         => \SDATASELInt[3]_net_1\, Y => N_202);
    
    \SDATASELInt[14]\ : SLE
      port map(D => \SADDRSEL[14]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[14]_net_1\);
    
    d_masterRegAddrSel_0_i_3_2 : CFG4
      generic map(INIT => x"CFCE")

      port map(A => \d_masterRegAddrSel_0_i_1_tz\, B => 
        \d_masterRegAddrSel_0_i_3_0\, C => masterRegAddrSel_net_1, 
        D => \N_401\, Y => \d_masterRegAddrSel_0_i_3_2\);
    
    \SDATASELInt[2]\ : SLE
      port map(D => \SADDRSEL[2]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[2]_net_1\);
    
    \SADDRSEL_0_a2_0_a2[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, B
         => N_394, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, Y
         => \SADDRSEL[3]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GATEDHWRITE_i_m3_i_m2 : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, C => 
        regHWRITE_net_1, Y => N_253);
    
    \SADDRSEL_0_a2_0_a2_0_0[7]\ : CFG2
      generic map(INIT => x"4")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        Y => \SADDRSEL_0_a2_0_a2_0_0[7]_net_1\);
    
    d_masterRegAddrSel_0_i_a0_1 : CFG4
      generic map(INIT => x"0004")

      port map(A => masterRegAddrSel_net_1, B => N_235, C => 
        \SDATASELInt[13]_net_1\, D => \SDATASELInt[2]_net_1\, Y
         => \d_masterRegAddrSel_0_i_a0_1\);
    
    \SADDRSEL_0_0_a2_1_RNISSES[15]\ : CFG3
      generic map(INIT => x"51")

      port map(A => arbRegSMCurrentState_13, B => \N_359\, C => 
        \N_321_2\, Y => SADDRSEL_0_0_0_1_0(0));
    
    \SADDRSEL_0_0_a2_1_RNI93LE1[15]\ : CFG4
      generic map(INIT => x"AAFB")

      port map(A => \N_321_2\, B => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), C
         => masterRegAddrSel_net_1, D => \N_359\, Y => 
        SADDRSEL_0_0_0_0(0));
    
    \SDATASELInt[13]\ : SLE
      port map(D => \SADDRSEL[13]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[13]_net_1\);
    
    \SADDRSEL_0_a2_0_a2[5]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => N_344, D => \SADDRSEL_0_a2_0_a2_0_0[7]_net_1\, Y => 
        \SADDRSEL[5]\);
    
    \regHWRITE\ : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => N_36_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHWRITE_net_1);
    
    d_masterRegAddrSel_0_1_i_2_0_RNI9AIT : CFG4
      generic map(INIT => x"0010")

      port map(A => \d_masterRegAddrSel_0_1_i_2_0\, B => 
        masterRegAddrSel_net_1, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), D
         => \d_masterRegAddrSel_0_1_i_2_1\, Y => N_36_i_1);
    
    hready_m_xhdl339_0_a5_0_a2 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_356, B => \xhdl1222[0]\, C => \N_355\, D
         => \N_354\, Y => \hready_m_xhdl339\);
    
    d_masterRegAddrSel_0_1_i_2_0 : CFG3
      generic map(INIT => x"EC")

      port map(A => \N_395\, B => N_286, C => \N_358\, Y => 
        \d_masterRegAddrSel_0_1_i_2_0\);
    
    \SDATASELInt[9]\ : SLE
      port map(D => \SADDRSEL[9]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[9]_net_1\);
    
    \SDATASELInt[1]\ : SLE
      port map(D => \SADDRSEL[1]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[1]_net_1\);
    
    \SDATASELInt[12]\ : SLE
      port map(D => \SADDRSEL[12]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[12]_net_1\);
    
    \SDATASELInt[0]\ : SLE
      port map(D => \xhdl1221[0]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \xhdl1222[0]\);
    
    \SADDRSEL_0_a2_0_a2_0[3]\ : CFG3
      generic map(INIT => x"04")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => N_344, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, Y
         => N_394);
    
    d_masterRegAddrSel_0_i_a2_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => \d_masterRegAddrSel_0_i_a2_0_0\, B => \N_354\, 
        C => \N_355\, D => N_210, Y => N_281);
    
    \SDATASELInt[5]\ : SLE
      port map(D => \SADDRSEL[5]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[5]_net_1\);
    
    \SADDRSEL_0_a2_0_a2[7]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => N_344, D => \SADDRSEL_0_a2_0_a2_0_0[7]_net_1\, Y => 
        \SADDRSEL[7]\);
    
    d_masterRegAddrSel_0_i_a2_0_0 : CFG2
      generic map(INIT => x"1")

      port map(A => masterRegAddrSel_net_1, B => 
        \SDATASELInt[11]_net_1\, Y => 
        \d_masterRegAddrSel_0_i_a2_0_0\);
    
    un1_hready_m_xhdl339_2_i_0_0_o2_0_0 : CFG3
      generic map(INIT => x"EC")

      port map(A => N_453_tz, B => \N_395\, C => N_357, Y => 
        \un1_hready_m_xhdl339_2_i_0_0_o2_0\);
    
    un1_hready_m_xhdl339_2_i_0_0_a2 : CFG3
      generic map(INIT => x"32")

      port map(A => \un1_hready_m_xhdl339_2_i_0_0_o2_0\, B => 
        \xhdl1222[0]\, C => N_397, Y => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0));
    
    \regHADDR[3]\ : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => N_36_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(3));
    
    \SDATASELInt[3]\ : SLE
      port map(D => \SADDRSEL[3]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[3]_net_1\);
    
    d_masterRegAddrSel_0_1_i_a2_5_2_1_0_RNINOVJ : CFG4
      generic map(INIT => x"0004")

      port map(A => arbRegSMCurrentState_13, B => 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0_net_1, C => 
        arbRegSMCurrentState_12, D => arbRegSMCurrentState_4, Y
         => \N_321_2\);
    
    hready_m_xhdl339_0_a5_0_a2_RNIUBPK : CFG2
      generic map(INIT => x"2")

      port map(A => \hready_m_xhdl339\, B => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, Y => N_299);
    
    \SDATASELInt[7]\ : SLE
      port map(D => \SADDRSEL[7]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[7]_net_1\);
    
    d_masterRegAddrSel_0_1_i_o2_0_0_d : CFG4
      generic map(INIT => x"A0EC")

      port map(A => \N_354\, B => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, C => \N_355\, D
         => \N_321_2\, Y => \d_masterRegAddrSel_0_1_i_o2_0_0_d\);
    
    \SADDRSEL_0_0_a2_0[15]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        D => N_360, Y => N_296);
    
    un1_hready_m_xhdl339_2_i_0_0_a2_2_RNIV1FO1 : CFG4
      generic map(INIT => x"0313")

      port map(A => \un1_hready_m_xhdl339_2_i_0_0_o2_0\, B => 
        N_299, C => \N_358\, D => N_397, Y => N_21_i_0);
    
    \SDATASELInt[6]\ : SLE
      port map(D => \SADDRSEL[6]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[6]_net_1\);
    
    masterRegAddrSel_RNO : CFG2
      generic map(INIT => x"2")

      port map(A => N_159, B => \d_masterRegAddrSel_0_i_3_2\, Y
         => N_30_i_0);
    
    d_masterRegAddrSel_0_1_i_a2_5_s_RNIIQ6H1 : CFG4
      generic map(INIT => x"00C4")

      port map(A => sha256_system_sb_0_AMBA_SLAVE_0_HREADY, B => 
        N_36_i_1, C => d_masterRegAddrSel_0_1_i_a2_5_out, D => 
        N_208, Y => N_36_i_0);
    
    \SADDRSEL_0_a2_2_a2[10]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        D => N_360, Y => \SADDRSEL[10]\);
    
    d_masterRegAddrSel_0_i_3_0 : CFG4
      generic map(INIT => x"F8F0")

      port map(A => \d_masterRegAddrSel_0_i_a0_1\, B => \N_354\, 
        C => N_281, D => \N_355\, Y => 
        \d_masterRegAddrSel_0_i_3_0\);
    
    \SADDRSEL_0_a2_1_a2_1[11]\ : CFG3
      generic map(INIT => x"20")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, B
         => masterRegAddrSel_net_1, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), Y
         => N_360);
    
    \SADDRSEL_0_a2_0_a2[1]\ : CFG3
      generic map(INIT => x"40")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, B
         => N_394, C => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, Y
         => \SADDRSEL[1]\);
    
    \SDATASELInt[11]\ : SLE
      port map(D => \SADDRSEL[11]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[11]_net_1\);
    
    d_masterRegAddrSel_0_1_i_a2_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_353, B => N_352, C => N_189, D => N_356, Y
         => \N_395\);
    
    \SADDRSEL_0_a2_1_a2[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => N_344, D => \SADDRSEL_0_a2_0_a2_0_0[7]_net_1\, Y => 
        \SADDRSEL[4]\);
    
    \SADDRSEL_0_a2_1_a2[12]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        D => N_360, Y => \SADDRSEL[12]\);
    
    d_masterRegAddrSel_0_1_i_o2_1 : CFG4
      generic map(INIT => x"0116")

      port map(A => \SDATASELInt[12]_net_1\, B => 
        \SDATASELInt[10]_net_1\, C => \SDATASELInt[8]_net_1\, D
         => \SDATASELInt[7]_net_1\, Y => N_189);
    
    \SDATASELInt[8]\ : SLE
      port map(D => \SADDRSEL[8]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[8]_net_1\);
    
    d_masterRegAddrSel_0_1_i_o2_2_RNICUV3 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_203, B => N_202, C => N_353, D => N_352, Y
         => N_453_tz);
    
    \SADDRSEL_0_0[0]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \N_359\, B => N_344, C => N_208, Y => 
        \xhdl1221[0]\);
    
    \regHADDR[4]\ : SLE
      port map(D => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, CLK
         => sha256_system_sb_0_FIC_0_CLK, EN => N_36_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(4));
    
    \SDATASELInt[10]\ : SLE
      port map(D => \SADDRSEL[10]\, CLK => 
        sha256_system_sb_0_FIC_0_CLK, EN => N_21_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[10]_net_1\);
    
    \SADDRSEL_0_a2_0_a2[13]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, B
         => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        C => sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        D => N_360, Y => \SADDRSEL[13]\);
    
    un1_hready_m_xhdl339_2_i_0_0_o2_0 : CFG3
      generic map(INIT => x"16")

      port map(A => \SDATASELInt[13]_net_1\, B => 
        \SDATASELInt[2]_net_1\, C => \SDATASELInt[11]_net_1\, Y
         => \N_211\);
    
    default_slave_sm : COREAHBLITE_DEFAULTSLAVESM_0
      port map(xhdl1222(0) => \xhdl1222[0]\, SDATASELInt_12 => 
        \SDATASELInt[13]_net_1\, SDATASELInt_1 => 
        \SDATASELInt[2]_net_1\, SDATASELInt_10 => 
        \SDATASELInt[11]_net_1\, SDATASELInt_5 => 
        \SDATASELInt[6]_net_1\, SDATASELInt_4 => 
        \SDATASELInt[5]_net_1\, SDATASELInt_3 => 
        \SDATASELInt[4]_net_1\, SDATASELInt_2 => 
        \SDATASELInt[3]_net_1\, SDATASELInt_14 => 
        \SDATASELInt[15]_net_1\, SDATASELInt_13 => 
        \SDATASELInt[14]_net_1\, SDATASELInt_8 => 
        \SDATASELInt[9]_net_1\, SDATASELInt_0 => 
        \SDATASELInt[1]_net_1\, defSlaveSMCurrentState => 
        defSlaveSMCurrentState, MSS_READY => MSS_READY, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, N_357 => N_357, 
        HREADY_M_iv_i_i_1_1 => HREADY_M_iv_i_i_1_1, N_358 => 
        \N_358\, N_453_tz => N_453_tz, HREADY_M_iv_i_i_1 => 
        HREADY_M_iv_i_i_1, N_356 => N_356, N_353 => N_353, N_352
         => N_352, N_354 => \N_354\, N_355 => \N_355\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MATRIX4X16 is

    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1);
          arbRegSMCurrentState_ns_i_0_0_0_a0_0                 : in    std_logic_vector(1 to 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          masterAddrInProg                                     : out   std_logic_vector(3 downto 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0);
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          arbRegSMCurrentState_13                              : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic;
          MSS_READY                                            : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic;
          regHWRITE                                            : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic;
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_358                                                : out   std_logic;
          N_401                                                : out   std_logic;
          N_403                                                : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic;
          N_208                                                : out   std_logic;
          N_211                                                : out   std_logic;
          N_354                                                : out   std_logic;
          N_355                                                : out   std_logic;
          N_395                                                : out   std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          N_23_i_0                                             : out   std_logic;
          N_359                                                : out   std_logic;
          N_253                                                : out   std_logic;
          N_344                                                : out   std_logic;
          N_321_2                                              : out   std_logic;
          N_36_2                                               : in    std_logic;
          N_48_i_0                                             : out   std_logic;
          N_46_i_0                                             : out   std_logic;
          N_44_i_0                                             : out   std_logic;
          N_42_i_0                                             : out   std_logic;
          N_16_i_0                                             : out   std_logic
        );

end COREAHBLITE_MATRIX4X16;

architecture DEF_ARCH of COREAHBLITE_MATRIX4X16 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVESTAGE_1
    port( masterAddrInProg                                     : out   std_logic_vector(3 downto 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0) := (others => 'U');
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          regHADDR                                             : in    std_logic_vector(5 downto 2) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1) := (others => 'U');
          arbRegSMCurrentState_ns_i_0_0_0_a0_0                 : in    std_logic_vector(1 to 1) := (others => 'U');
          SADDRSEL_0_0_0_1_0                                   : in    std_logic_vector(0 to 0) := (others => 'U');
          SADDRSEL_0_0_0_0                                     : in    std_logic_vector(0 to 0) := (others => 'U');
          masterDataInProg_0                                   : out   std_logic;
          arbRegSMCurrentState_13                              : out   std_logic;
          arbRegSMCurrentState_12                              : out   std_logic;
          arbRegSMCurrentState_8                               : out   std_logic;
          arbRegSMCurrentState_4                               : out   std_logic;
          arbRegSMCurrentState_0                               : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic := 'U';
          MSS_READY                                            : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic := 'U';
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic := 'U';
          N_321_2                                              : in    std_logic := 'U';
          masterRegAddrSel                                     : in    std_logic := 'U';
          N_359                                                : in    std_logic := 'U';
          N_344                                                : out   std_logic;
          N_208                                                : out   std_logic;
          d_masterRegAddrSel_0_1_i_a2_5_2_1_0                  : in    std_logic := 'U';
          N_253                                                : in    std_logic := 'U';
          N_48_i_0                                             : out   std_logic;
          N_46_i_0                                             : out   std_logic;
          N_44_i_0                                             : out   std_logic;
          N_42_i_0                                             : out   std_logic;
          N_16_i_0                                             : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MASTERSTAGE_2_1_0_1_0
    port( regHADDR                                             : out   std_logic_vector(5 downto 2);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1) := (others => 'U');
          masterDataInProg                                     : in    std_logic_vector(0 to 0) := (others => 'U');
          SADDRSEL_0_0_0_0                                     : out   std_logic_vector(0 to 0);
          SADDRSEL_0_0_0_1_0                                   : out   std_logic_vector(0 to 0);
          arbRegSMCurrentState_ns_i_0_0_0_a0_0                 : in    std_logic_vector(1 to 1) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          arbRegSMCurrentState_0                               : in    std_logic := 'U';
          arbRegSMCurrentState_8                               : in    std_logic := 'U';
          arbRegSMCurrentState_13                              : in    std_logic := 'U';
          arbRegSMCurrentState_12                              : in    std_logic := 'U';
          arbRegSMCurrentState_4                               : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic := 'U';
          MSS_READY                                            : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic := 'U';
          regHWRITE                                            : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_358                                                : out   std_logic;
          N_401                                                : out   std_logic;
          N_403                                                : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic := 'U';
          N_208                                                : in    std_logic := 'U';
          N_211                                                : out   std_logic;
          N_354                                                : out   std_logic;
          N_355                                                : out   std_logic;
          N_395                                                : out   std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          N_23_i_0                                             : out   std_logic;
          d_masterRegAddrSel_0_1_i_a2_5_2_1_0                  : out   std_logic;
          N_359                                                : out   std_logic;
          N_253                                                : out   std_logic;
          N_344                                                : in    std_logic := 'U';
          N_321_2                                              : out   std_logic;
          N_36_2                                               : in    std_logic := 'U'
        );
  end component;

    signal \regHADDR[2]\, \regHADDR[3]\, \regHADDR[4]\, 
        \regHADDR[5]\, \masterDataInProg[0]\, 
        \arbRegSMCurrentState[2]\, \arbRegSMCurrentState[10]\, 
        \arbRegSMCurrentState_13\, \arbRegSMCurrentState[14]\, 
        \arbRegSMCurrentState[6]\, \SADDRSEL_0_0_0_0[0]\, 
        \SADDRSEL_0_0_0_1_0[0]\, \masterRegAddrSel\, \N_208\, 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0, \N_359\, \N_253\, 
        \N_344\, \N_321_2\, GND_net_1, VCC_net_1 : std_logic;

    for all : COREAHBLITE_SLAVESTAGE_1
	Use entity work.COREAHBLITE_SLAVESTAGE_1(DEF_ARCH);
    for all : COREAHBLITE_MASTERSTAGE_2_1_0_1_0
	Use entity work.COREAHBLITE_MASTERSTAGE_2_1_0_1_0(DEF_ARCH);
begin 

    arbRegSMCurrentState_13 <= \arbRegSMCurrentState_13\;
    masterRegAddrSel <= \masterRegAddrSel\;
    N_208 <= \N_208\;
    N_359 <= \N_359\;
    N_253 <= \N_253\;
    N_344 <= \N_344\;
    N_321_2 <= \N_321_2\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    slavestage_0 : COREAHBLITE_SLAVESTAGE_1
      port map(masterAddrInProg(3) => masterAddrInProg(3), 
        masterAddrInProg(2) => masterAddrInProg(2), 
        masterAddrInProg(1) => masterAddrInProg(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        AHB_slave_dummy_0_mem_wdata(31) => 
        AHB_slave_dummy_0_mem_wdata(31), 
        AHB_slave_dummy_0_mem_wdata(30) => 
        AHB_slave_dummy_0_mem_wdata(30), 
        AHB_slave_dummy_0_mem_wdata(29) => 
        AHB_slave_dummy_0_mem_wdata(29), 
        AHB_slave_dummy_0_mem_wdata(28) => 
        AHB_slave_dummy_0_mem_wdata(28), 
        AHB_slave_dummy_0_mem_wdata(27) => 
        AHB_slave_dummy_0_mem_wdata(27), 
        AHB_slave_dummy_0_mem_wdata(26) => 
        AHB_slave_dummy_0_mem_wdata(26), 
        AHB_slave_dummy_0_mem_wdata(25) => 
        AHB_slave_dummy_0_mem_wdata(25), 
        AHB_slave_dummy_0_mem_wdata(24) => 
        AHB_slave_dummy_0_mem_wdata(24), 
        AHB_slave_dummy_0_mem_wdata(23) => 
        AHB_slave_dummy_0_mem_wdata(23), 
        AHB_slave_dummy_0_mem_wdata(22) => 
        AHB_slave_dummy_0_mem_wdata(22), 
        AHB_slave_dummy_0_mem_wdata(21) => 
        AHB_slave_dummy_0_mem_wdata(21), 
        AHB_slave_dummy_0_mem_wdata(20) => 
        AHB_slave_dummy_0_mem_wdata(20), 
        AHB_slave_dummy_0_mem_wdata(19) => 
        AHB_slave_dummy_0_mem_wdata(19), 
        AHB_slave_dummy_0_mem_wdata(18) => 
        AHB_slave_dummy_0_mem_wdata(18), 
        AHB_slave_dummy_0_mem_wdata(17) => 
        AHB_slave_dummy_0_mem_wdata(17), 
        AHB_slave_dummy_0_mem_wdata(16) => 
        AHB_slave_dummy_0_mem_wdata(16), 
        AHB_slave_dummy_0_mem_wdata(15) => 
        AHB_slave_dummy_0_mem_wdata(15), 
        AHB_slave_dummy_0_mem_wdata(14) => 
        AHB_slave_dummy_0_mem_wdata(14), 
        AHB_slave_dummy_0_mem_wdata(13) => 
        AHB_slave_dummy_0_mem_wdata(13), 
        AHB_slave_dummy_0_mem_wdata(12) => 
        AHB_slave_dummy_0_mem_wdata(12), 
        AHB_slave_dummy_0_mem_wdata(11) => 
        AHB_slave_dummy_0_mem_wdata(11), 
        AHB_slave_dummy_0_mem_wdata(10) => 
        AHB_slave_dummy_0_mem_wdata(10), 
        AHB_slave_dummy_0_mem_wdata(9) => 
        AHB_slave_dummy_0_mem_wdata(9), 
        AHB_slave_dummy_0_mem_wdata(8) => 
        AHB_slave_dummy_0_mem_wdata(8), 
        AHB_slave_dummy_0_mem_wdata(7) => 
        AHB_slave_dummy_0_mem_wdata(7), 
        AHB_slave_dummy_0_mem_wdata(6) => 
        AHB_slave_dummy_0_mem_wdata(6), 
        AHB_slave_dummy_0_mem_wdata(5) => 
        AHB_slave_dummy_0_mem_wdata(5), 
        AHB_slave_dummy_0_mem_wdata(4) => 
        AHB_slave_dummy_0_mem_wdata(4), 
        AHB_slave_dummy_0_mem_wdata(3) => 
        AHB_slave_dummy_0_mem_wdata(3), 
        AHB_slave_dummy_0_mem_wdata(2) => 
        AHB_slave_dummy_0_mem_wdata(2), 
        AHB_slave_dummy_0_mem_wdata(1) => 
        AHB_slave_dummy_0_mem_wdata(1), 
        AHB_slave_dummy_0_mem_wdata(0) => 
        AHB_slave_dummy_0_mem_wdata(0), regHADDR(5) => 
        \regHADDR[5]\, regHADDR(4) => \regHADDR[4]\, regHADDR(3)
         => \regHADDR[3]\, regHADDR(2) => \regHADDR[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1) => 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1), 
        SADDRSEL_0_0_0_1_0(0) => \SADDRSEL_0_0_0_1_0[0]\, 
        SADDRSEL_0_0_0_0(0) => \SADDRSEL_0_0_0_0[0]\, 
        masterDataInProg_0 => \masterDataInProg[0]\, 
        arbRegSMCurrentState_13 => \arbRegSMCurrentState_13\, 
        arbRegSMCurrentState_12 => \arbRegSMCurrentState[14]\, 
        arbRegSMCurrentState_8 => \arbRegSMCurrentState[10]\, 
        arbRegSMCurrentState_4 => \arbRegSMCurrentState[6]\, 
        arbRegSMCurrentState_0 => \arbRegSMCurrentState[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, 
        MSS_READY => MSS_READY, sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, N_321_2 => 
        \N_321_2\, masterRegAddrSel => \masterRegAddrSel\, N_359
         => \N_359\, N_344 => \N_344\, N_208 => \N_208\, 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0 => 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0, N_253 => \N_253\, 
        N_48_i_0 => N_48_i_0, N_46_i_0 => N_46_i_0, N_44_i_0 => 
        N_44_i_0, N_42_i_0 => N_42_i_0, N_16_i_0 => N_16_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    masterstage_0 : COREAHBLITE_MASTERSTAGE_2_1_0_1_0
      port map(regHADDR(5) => \regHADDR[5]\, regHADDR(4) => 
        \regHADDR[4]\, regHADDR(3) => \regHADDR[3]\, regHADDR(2)
         => \regHADDR[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        masterDataInProg(0) => \masterDataInProg[0]\, 
        SADDRSEL_0_0_0_0(0) => \SADDRSEL_0_0_0_0[0]\, 
        SADDRSEL_0_0_0_1_0(0) => \SADDRSEL_0_0_0_1_0[0]\, 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1) => 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        arbRegSMCurrentState_0 => \arbRegSMCurrentState[2]\, 
        arbRegSMCurrentState_8 => \arbRegSMCurrentState[10]\, 
        arbRegSMCurrentState_13 => \arbRegSMCurrentState_13\, 
        arbRegSMCurrentState_12 => \arbRegSMCurrentState[14]\, 
        arbRegSMCurrentState_4 => \arbRegSMCurrentState[6]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        MSS_READY => MSS_READY, sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, regHWRITE => regHWRITE, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        regHTRANS => regHTRANS, masterRegAddrSel => 
        \masterRegAddrSel\, N_358 => N_358, N_401 => N_401, N_403
         => N_403, sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, N_208 => \N_208\, 
        N_211 => N_211, N_354 => N_354, N_355 => N_355, N_395 => 
        N_395, hready_m_xhdl339 => hready_m_xhdl339, N_23_i_0 => 
        N_23_i_0, d_masterRegAddrSel_0_1_i_a2_5_2_1_0 => 
        d_masterRegAddrSel_0_1_i_a2_5_2_1_0, N_359 => \N_359\, 
        N_253 => \N_253\, N_344 => \N_344\, N_321_2 => \N_321_2\, 
        N_36_2 => N_36_2);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLite is

    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1);
          arbRegSMCurrentState                                 : out   std_logic_vector(15 to 15);
          arbRegSMCurrentState_ns_i_0_0_0_a0_0                 : in    std_logic_vector(1 to 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          masterAddrInProg                                     : out   std_logic_vector(3 downto 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0);
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic;
          MSS_READY                                            : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic;
          regHWRITE                                            : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic;
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_358                                                : out   std_logic;
          N_401                                                : out   std_logic;
          N_403                                                : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic;
          N_208                                                : out   std_logic;
          N_211                                                : out   std_logic;
          N_354                                                : out   std_logic;
          N_355                                                : out   std_logic;
          N_395                                                : out   std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          N_23_i_0                                             : out   std_logic;
          N_359                                                : out   std_logic;
          N_253                                                : out   std_logic;
          N_344                                                : out   std_logic;
          N_321_2                                              : out   std_logic;
          N_36_2                                               : in    std_logic;
          N_48_i_0                                             : out   std_logic;
          N_46_i_0                                             : out   std_logic;
          N_44_i_0                                             : out   std_logic;
          N_42_i_0                                             : out   std_logic;
          N_16_i_0                                             : out   std_logic
        );

end CoreAHBLite;

architecture DEF_ARCH of CoreAHBLite is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MATRIX4X16
    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1) := (others => 'U');
          arbRegSMCurrentState_ns_i_0_0_0_a0_0                 : in    std_logic_vector(1 to 1) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          masterAddrInProg                                     : out   std_logic_vector(3 downto 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0) := (others => 'U');
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          arbRegSMCurrentState_13                              : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic := 'U';
          MSS_READY                                            : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic := 'U';
          regHWRITE                                            : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_358                                                : out   std_logic;
          N_401                                                : out   std_logic;
          N_403                                                : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic := 'U';
          N_208                                                : out   std_logic;
          N_211                                                : out   std_logic;
          N_354                                                : out   std_logic;
          N_355                                                : out   std_logic;
          N_395                                                : out   std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          N_23_i_0                                             : out   std_logic;
          N_359                                                : out   std_logic;
          N_253                                                : out   std_logic;
          N_344                                                : out   std_logic;
          N_321_2                                              : out   std_logic;
          N_36_2                                               : in    std_logic := 'U';
          N_48_i_0                                             : out   std_logic;
          N_46_i_0                                             : out   std_logic;
          N_44_i_0                                             : out   std_logic;
          N_42_i_0                                             : out   std_logic;
          N_16_i_0                                             : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : COREAHBLITE_MATRIX4X16
	Use entity work.COREAHBLITE_MATRIX4X16(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    matrix4x16 : COREAHBLITE_MATRIX4X16
      port map(
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1) => 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        masterAddrInProg(3) => masterAddrInProg(3), 
        masterAddrInProg(2) => masterAddrInProg(2), 
        masterAddrInProg(1) => masterAddrInProg(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        AHB_slave_dummy_0_mem_wdata(31) => 
        AHB_slave_dummy_0_mem_wdata(31), 
        AHB_slave_dummy_0_mem_wdata(30) => 
        AHB_slave_dummy_0_mem_wdata(30), 
        AHB_slave_dummy_0_mem_wdata(29) => 
        AHB_slave_dummy_0_mem_wdata(29), 
        AHB_slave_dummy_0_mem_wdata(28) => 
        AHB_slave_dummy_0_mem_wdata(28), 
        AHB_slave_dummy_0_mem_wdata(27) => 
        AHB_slave_dummy_0_mem_wdata(27), 
        AHB_slave_dummy_0_mem_wdata(26) => 
        AHB_slave_dummy_0_mem_wdata(26), 
        AHB_slave_dummy_0_mem_wdata(25) => 
        AHB_slave_dummy_0_mem_wdata(25), 
        AHB_slave_dummy_0_mem_wdata(24) => 
        AHB_slave_dummy_0_mem_wdata(24), 
        AHB_slave_dummy_0_mem_wdata(23) => 
        AHB_slave_dummy_0_mem_wdata(23), 
        AHB_slave_dummy_0_mem_wdata(22) => 
        AHB_slave_dummy_0_mem_wdata(22), 
        AHB_slave_dummy_0_mem_wdata(21) => 
        AHB_slave_dummy_0_mem_wdata(21), 
        AHB_slave_dummy_0_mem_wdata(20) => 
        AHB_slave_dummy_0_mem_wdata(20), 
        AHB_slave_dummy_0_mem_wdata(19) => 
        AHB_slave_dummy_0_mem_wdata(19), 
        AHB_slave_dummy_0_mem_wdata(18) => 
        AHB_slave_dummy_0_mem_wdata(18), 
        AHB_slave_dummy_0_mem_wdata(17) => 
        AHB_slave_dummy_0_mem_wdata(17), 
        AHB_slave_dummy_0_mem_wdata(16) => 
        AHB_slave_dummy_0_mem_wdata(16), 
        AHB_slave_dummy_0_mem_wdata(15) => 
        AHB_slave_dummy_0_mem_wdata(15), 
        AHB_slave_dummy_0_mem_wdata(14) => 
        AHB_slave_dummy_0_mem_wdata(14), 
        AHB_slave_dummy_0_mem_wdata(13) => 
        AHB_slave_dummy_0_mem_wdata(13), 
        AHB_slave_dummy_0_mem_wdata(12) => 
        AHB_slave_dummy_0_mem_wdata(12), 
        AHB_slave_dummy_0_mem_wdata(11) => 
        AHB_slave_dummy_0_mem_wdata(11), 
        AHB_slave_dummy_0_mem_wdata(10) => 
        AHB_slave_dummy_0_mem_wdata(10), 
        AHB_slave_dummy_0_mem_wdata(9) => 
        AHB_slave_dummy_0_mem_wdata(9), 
        AHB_slave_dummy_0_mem_wdata(8) => 
        AHB_slave_dummy_0_mem_wdata(8), 
        AHB_slave_dummy_0_mem_wdata(7) => 
        AHB_slave_dummy_0_mem_wdata(7), 
        AHB_slave_dummy_0_mem_wdata(6) => 
        AHB_slave_dummy_0_mem_wdata(6), 
        AHB_slave_dummy_0_mem_wdata(5) => 
        AHB_slave_dummy_0_mem_wdata(5), 
        AHB_slave_dummy_0_mem_wdata(4) => 
        AHB_slave_dummy_0_mem_wdata(4), 
        AHB_slave_dummy_0_mem_wdata(3) => 
        AHB_slave_dummy_0_mem_wdata(3), 
        AHB_slave_dummy_0_mem_wdata(2) => 
        AHB_slave_dummy_0_mem_wdata(2), 
        AHB_slave_dummy_0_mem_wdata(1) => 
        AHB_slave_dummy_0_mem_wdata(1), 
        AHB_slave_dummy_0_mem_wdata(0) => 
        AHB_slave_dummy_0_mem_wdata(0), arbRegSMCurrentState_13
         => arbRegSMCurrentState(15), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        MSS_READY => MSS_READY, sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, regHWRITE => regHWRITE, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        regHTRANS => regHTRANS, masterRegAddrSel => 
        masterRegAddrSel, N_358 => N_358, N_401 => N_401, N_403
         => N_403, sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, N_208 => N_208, 
        N_211 => N_211, N_354 => N_354, N_355 => N_355, N_395 => 
        N_395, hready_m_xhdl339 => hready_m_xhdl339, N_23_i_0 => 
        N_23_i_0, N_359 => N_359, N_253 => N_253, N_344 => N_344, 
        N_321_2 => N_321_2, N_36_2 => N_36_2, N_48_i_0 => 
        N_48_i_0, N_46_i_0 => N_46_i_0, N_44_i_0 => N_44_i_0, 
        N_42_i_0 => N_42_i_0, N_16_i_0 => N_16_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_system_sb_CCC_0_FCCC is

    port( sha256_system_sb_0_FIC_0_CLK                       : out   std_logic;
          FIC_0_LOCK                                         : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic
        );

end sha256_system_sb_CCC_0_FCCC;

architecture DEF_ARCH of sha256_system_sb_CCC_0_FCCC is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => sha256_system_sb_0_FIC_0_CLK);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007FB8000044D74000318C6318C1F18C61EC0404040400301",
         VCOFREQUENCY => 800.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => FIC_0_LOCK, 
        BUSY => OPEN, CLK0 => VCC_net_1, CLK1 => VCC_net_1, CLK2
         => VCC_net_1, CLK3 => VCC_net_1, NGMUX0_SEL => GND_net_1, 
        NGMUX1_SEL => GND_net_1, NGMUX2_SEL => GND_net_1, 
        NGMUX3_SEL => GND_net_1, NGMUX0_HOLD_N => VCC_net_1, 
        NGMUX1_HOLD_N => VCC_net_1, NGMUX2_HOLD_N => VCC_net_1, 
        NGMUX3_HOLD_N => VCC_net_1, NGMUX0_ARST_N => VCC_net_1, 
        NGMUX1_ARST_N => VCC_net_1, NGMUX2_ARST_N => VCC_net_1, 
        NGMUX3_ARST_N => VCC_net_1, PLL_BYPASS_N => VCC_net_1, 
        PLL_ARST_N => VCC_net_1, PLL_POWERDOWN_N => VCC_net_1, 
        GPD0_ARST_N => VCC_net_1, GPD1_ARST_N => VCC_net_1, 
        GPD2_ARST_N => VCC_net_1, GPD3_ARST_N => VCC_net_1, 
        PRESET_N => GND_net_1, PCLK => VCC_net_1, PSEL => 
        VCC_net_1, PENABLE => VCC_net_1, PWRITE => VCC_net_1, 
        PADDR(7) => VCC_net_1, PADDR(6) => VCC_net_1, PADDR(5)
         => VCC_net_1, PADDR(4) => VCC_net_1, PADDR(3) => 
        VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7) => VCC_net_1, 
        PWDATA(6) => VCC_net_1, PWDATA(5) => VCC_net_1, PWDATA(4)
         => VCC_net_1, PWDATA(3) => VCC_net_1, PWDATA(2) => 
        VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0) => VCC_net_1, 
        CLK0_PAD => GND_net_1, CLK1_PAD => GND_net_1, CLK2_PAD
         => GND_net_1, CLK3_PAD => GND_net_1, GL0 => GL0_net, GL1
         => OPEN, GL2 => OPEN, GL3 => OPEN, RCOSC_25_50MHZ => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        RCOSC_1MHZ => GND_net_1, XTLOSC => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_system_sb is

    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : inout std_logic_vector(1 to 1) := (others => 'Z');
          arbRegSMCurrentState                                 : out   std_logic_vector(15 to 15);
          masterAddrInProg                                     : out   std_logic_vector(3 downto 1);
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : inout std_logic := 'Z';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : inout std_logic := 'Z';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : inout std_logic := 'Z';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : inout std_logic := 'Z';
          data_out_9_0_29                                      : in    std_logic;
          data_out_9_0_31                                      : in    std_logic;
          data_out_9_0_1                                       : in    std_logic;
          data_out_9_0_0                                       : in    std_logic;
          sha256_system_sb_0_POWER_ON_RESET_N                  : out   std_logic;
          DEVRST_N                                             : in    std_logic;
          sha256_system_sb_0_FIC_0_CLK                         : out   std_logic;
          regHWRITE                                            : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : inout std_logic := 'Z';
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_358                                                : out   std_logic;
          N_401                                                : out   std_logic;
          N_403                                                : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic;
          N_208                                                : out   std_logic;
          N_211                                                : out   std_logic;
          N_354                                                : out   std_logic;
          N_355                                                : out   std_logic;
          N_395                                                : out   std_logic;
          N_359                                                : out   std_logic;
          N_253                                                : out   std_logic;
          N_344                                                : out   std_logic;
          N_321_2                                              : out   std_logic;
          N_36_2                                               : in    std_logic;
          N_48_i_0                                             : out   std_logic;
          N_46_i_0                                             : out   std_logic;
          N_44_i_0                                             : out   std_logic;
          N_42_i_0                                             : out   std_logic;
          N_16_i_0                                             : out   std_logic;
          N_1256                                               : in    std_logic;
          data_out_sn_N_12_mux                                 : in    std_logic;
          N_1323                                               : in    std_logic;
          N_1257                                               : in    std_logic;
          N_1324                                               : in    std_logic;
          N_1258                                               : in    std_logic;
          N_1325                                               : in    std_logic;
          N_1259                                               : in    std_logic;
          N_1326                                               : in    std_logic;
          N_1260                                               : in    std_logic;
          N_1327                                               : in    std_logic;
          N_1261                                               : in    std_logic;
          N_1328                                               : in    std_logic;
          N_1262                                               : in    std_logic;
          N_1329                                               : in    std_logic;
          N_1263                                               : in    std_logic;
          N_1330                                               : in    std_logic;
          N_1264                                               : in    std_logic;
          N_1331                                               : in    std_logic;
          N_1265                                               : in    std_logic;
          N_1332                                               : in    std_logic;
          N_1266                                               : in    std_logic;
          N_1333                                               : in    std_logic;
          N_1267                                               : in    std_logic;
          N_1334                                               : in    std_logic;
          N_1268                                               : in    std_logic;
          N_1335                                               : in    std_logic;
          N_1269                                               : in    std_logic;
          N_1336                                               : in    std_logic;
          N_1270                                               : in    std_logic;
          N_1337                                               : in    std_logic;
          N_1271                                               : in    std_logic;
          N_1338                                               : in    std_logic;
          N_1272                                               : in    std_logic;
          N_1339                                               : in    std_logic;
          N_1273                                               : in    std_logic;
          N_1340                                               : in    std_logic;
          N_1274                                               : in    std_logic;
          N_1341                                               : in    std_logic;
          N_1275                                               : in    std_logic;
          N_1342                                               : in    std_logic;
          N_1276                                               : in    std_logic;
          N_1343                                               : in    std_logic;
          N_1277                                               : in    std_logic;
          N_1344                                               : in    std_logic;
          N_1278                                               : in    std_logic;
          N_1345                                               : in    std_logic;
          N_1279                                               : in    std_logic;
          N_1346                                               : in    std_logic;
          N_1280                                               : in    std_logic;
          N_1347                                               : in    std_logic;
          N_1281                                               : in    std_logic;
          N_1348                                               : in    std_logic;
          N_1282                                               : in    std_logic;
          N_1349                                               : in    std_logic;
          N_1284                                               : in    std_logic;
          N_1351                                               : in    std_logic;
          N_1446                                               : in    std_logic;
          N_1423_3                                             : in    std_logic;
          N_53                                                 : in    std_logic;
          N_1457                                               : in    std_logic;
          N_1458                                               : in    std_logic;
          GPIO_2_M2F_c                                         : out   std_logic;
          GPIO_1_M2F_c                                         : out   std_logic;
          GPIO_0_M2F_c                                         : out   std_logic
        );

end sha256_system_sb;

architecture DEF_ARCH of sha256_system_sb is 

  component sha256_system_sb_MSS
    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : inout   std_logic_vector(1 to 1);
          arbRegSMCurrentState_ns_i_0_0_0_a0_0                 : out   std_logic_vector(1 to 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : out   std_logic_vector(31 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : in    std_logic_vector(0 to 0) := (others => 'U');
          data_out_9_0_29                                      : in    std_logic := 'U';
          data_out_9_0_31                                      : in    std_logic := 'U';
          data_out_9_0_1                                       : in    std_logic := 'U';
          data_out_9_0_0                                       : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_26 : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_27 : out   std_logic;
          masterRegAddrSel                                     : in    std_logic := 'U';
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic := 'U';
          N_1256                                               : in    std_logic := 'U';
          data_out_sn_N_12_mux                                 : in    std_logic := 'U';
          N_1323                                               : in    std_logic := 'U';
          hready_m_xhdl339                                     : in    std_logic := 'U';
          N_1257                                               : in    std_logic := 'U';
          N_1324                                               : in    std_logic := 'U';
          N_1258                                               : in    std_logic := 'U';
          N_1325                                               : in    std_logic := 'U';
          N_1259                                               : in    std_logic := 'U';
          N_1326                                               : in    std_logic := 'U';
          N_1260                                               : in    std_logic := 'U';
          N_1327                                               : in    std_logic := 'U';
          N_1261                                               : in    std_logic := 'U';
          N_1328                                               : in    std_logic := 'U';
          N_1262                                               : in    std_logic := 'U';
          N_1329                                               : in    std_logic := 'U';
          N_1263                                               : in    std_logic := 'U';
          N_1330                                               : in    std_logic := 'U';
          N_1264                                               : in    std_logic := 'U';
          N_1331                                               : in    std_logic := 'U';
          N_1265                                               : in    std_logic := 'U';
          N_1332                                               : in    std_logic := 'U';
          N_1266                                               : in    std_logic := 'U';
          N_1333                                               : in    std_logic := 'U';
          N_1267                                               : in    std_logic := 'U';
          N_1334                                               : in    std_logic := 'U';
          N_1268                                               : in    std_logic := 'U';
          N_1335                                               : in    std_logic := 'U';
          N_1269                                               : in    std_logic := 'U';
          N_1336                                               : in    std_logic := 'U';
          N_1270                                               : in    std_logic := 'U';
          N_1337                                               : in    std_logic := 'U';
          N_1271                                               : in    std_logic := 'U';
          N_1338                                               : in    std_logic := 'U';
          N_1272                                               : in    std_logic := 'U';
          N_1339                                               : in    std_logic := 'U';
          N_1273                                               : in    std_logic := 'U';
          N_1340                                               : in    std_logic := 'U';
          N_1274                                               : in    std_logic := 'U';
          N_1341                                               : in    std_logic := 'U';
          N_1275                                               : in    std_logic := 'U';
          N_1342                                               : in    std_logic := 'U';
          N_1276                                               : in    std_logic := 'U';
          N_1343                                               : in    std_logic := 'U';
          N_1277                                               : in    std_logic := 'U';
          N_1344                                               : in    std_logic := 'U';
          N_1278                                               : in    std_logic := 'U';
          N_1345                                               : in    std_logic := 'U';
          N_1279                                               : in    std_logic := 'U';
          N_1346                                               : in    std_logic := 'U';
          N_1280                                               : in    std_logic := 'U';
          N_1347                                               : in    std_logic := 'U';
          N_1281                                               : in    std_logic := 'U';
          N_1348                                               : in    std_logic := 'U';
          N_1282                                               : in    std_logic := 'U';
          N_1349                                               : in    std_logic := 'U';
          N_1284                                               : in    std_logic := 'U';
          N_1351                                               : in    std_logic := 'U';
          N_1446                                               : in    std_logic := 'U';
          N_1423_3                                             : in    std_logic := 'U';
          N_53                                                 : in    std_logic := 'U';
          N_1457                                               : in    std_logic := 'U';
          N_1458                                               : in    std_logic := 'U';
          GPIO_2_M2F_c                                         : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N      : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : out   std_logic;
          sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F           : out   std_logic;
          GPIO_1_M2F_c                                         : out   std_logic;
          GPIO_0_M2F_c                                         : out   std_logic;
          N_23_i_0                                             : in    std_logic := 'U';
          FIC_0_LOCK                                           : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic := 'U'
        );
  end component;

  component sha256_system_sb_FABOSC_0_OSC
    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );
  end component;

  component CoreResetP
    port( MSS_READY                                       : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK                    : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic := 'U';
          sha256_system_sb_0_POWER_ON_RESET_N             : in    std_logic := 'U'
        );
  end component;

  component CoreAHBLite
    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1) := (others => 'U');
          arbRegSMCurrentState                                 : out   std_logic_vector(15 to 15);
          arbRegSMCurrentState_ns_i_0_0_0_a0_0                 : in    std_logic_vector(1 to 1) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          masterAddrInProg                                     : out   std_logic_vector(3 downto 1);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0) := (others => 'U');
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : in    std_logic := 'U';
          MSS_READY                                            : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : in    std_logic := 'U';
          regHWRITE                                            : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_358                                                : out   std_logic;
          N_401                                                : out   std_logic;
          N_403                                                : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic := 'U';
          N_208                                                : out   std_logic;
          N_211                                                : out   std_logic;
          N_354                                                : out   std_logic;
          N_355                                                : out   std_logic;
          N_395                                                : out   std_logic;
          hready_m_xhdl339                                     : out   std_logic;
          N_23_i_0                                             : out   std_logic;
          N_359                                                : out   std_logic;
          N_253                                                : out   std_logic;
          N_344                                                : out   std_logic;
          N_321_2                                              : out   std_logic;
          N_36_2                                               : in    std_logic := 'U';
          N_48_i_0                                             : out   std_logic;
          N_46_i_0                                             : out   std_logic;
          N_44_i_0                                             : out   std_logic;
          N_42_i_0                                             : out   std_logic;
          N_16_i_0                                             : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component sha256_system_sb_CCC_0_FCCC
    port( sha256_system_sb_0_FIC_0_CLK                       : out   std_logic;
          FIC_0_LOCK                                         : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

    signal \sha256_system_sb_0_POWER_ON_RESET_N\, \SYSRESET_POR\, 
        \sha256_system_sb_0_FIC_0_CLK\, FIC_0_LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        \arbRegSMCurrentState_ns_i_0_0_0_a0_0[1]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        MSS_READY, \masterRegAddrSel\, hready_m_xhdl339, N_23_i_0, 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        GND_net_1, VCC_net_1 : std_logic;

    for all : sha256_system_sb_MSS
	Use entity work.sha256_system_sb_MSS(DEF_ARCH);
    for all : sha256_system_sb_FABOSC_0_OSC
	Use entity work.sha256_system_sb_FABOSC_0_OSC(DEF_ARCH);
    for all : CoreResetP
	Use entity work.CoreResetP(DEF_ARCH);
    for all : CoreAHBLite
	Use entity work.CoreAHBLite(DEF_ARCH);
    for all : sha256_system_sb_CCC_0_FCCC
	Use entity work.sha256_system_sb_CCC_0_FCCC(DEF_ARCH);
begin 

    sha256_system_sb_0_POWER_ON_RESET_N <= 
        \sha256_system_sb_0_POWER_ON_RESET_N\;
    sha256_system_sb_0_FIC_0_CLK <= 
        \sha256_system_sb_0_FIC_0_CLK\;
    masterRegAddrSel <= \masterRegAddrSel\;

    sha256_system_sb_MSS_0 : sha256_system_sb_MSS
      port map(
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1) => 
        \arbRegSMCurrentState_ns_i_0_0_0_a0_0[1]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        data_out_9_0_29 => data_out_9_0_29, data_out_9_0_31 => 
        data_out_9_0_31, data_out_9_0_1 => data_out_9_0_1, 
        data_out_9_0_0 => data_out_9_0_0, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_26 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_27 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, 
        masterRegAddrSel => \masterRegAddrSel\, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, N_1256 => N_1256, 
        data_out_sn_N_12_mux => data_out_sn_N_12_mux, N_1323 => 
        N_1323, hready_m_xhdl339 => hready_m_xhdl339, N_1257 => 
        N_1257, N_1324 => N_1324, N_1258 => N_1258, N_1325 => 
        N_1325, N_1259 => N_1259, N_1326 => N_1326, N_1260 => 
        N_1260, N_1327 => N_1327, N_1261 => N_1261, N_1328 => 
        N_1328, N_1262 => N_1262, N_1329 => N_1329, N_1263 => 
        N_1263, N_1330 => N_1330, N_1264 => N_1264, N_1331 => 
        N_1331, N_1265 => N_1265, N_1332 => N_1332, N_1266 => 
        N_1266, N_1333 => N_1333, N_1267 => N_1267, N_1334 => 
        N_1334, N_1268 => N_1268, N_1335 => N_1335, N_1269 => 
        N_1269, N_1336 => N_1336, N_1270 => N_1270, N_1337 => 
        N_1337, N_1271 => N_1271, N_1338 => N_1338, N_1272 => 
        N_1272, N_1339 => N_1339, N_1273 => N_1273, N_1340 => 
        N_1340, N_1274 => N_1274, N_1341 => N_1341, N_1275 => 
        N_1275, N_1342 => N_1342, N_1276 => N_1276, N_1343 => 
        N_1343, N_1277 => N_1277, N_1344 => N_1344, N_1278 => 
        N_1278, N_1345 => N_1345, N_1279 => N_1279, N_1346 => 
        N_1346, N_1280 => N_1280, N_1347 => N_1347, N_1281 => 
        N_1281, N_1348 => N_1348, N_1282 => N_1282, N_1349 => 
        N_1349, N_1284 => N_1284, N_1351 => N_1351, N_1446 => 
        N_1446, N_1423_3 => N_1423_3, N_53 => N_53, N_1457 => 
        N_1457, N_1458 => N_1458, GPIO_2_M2F_c => GPIO_2_M2F_c, 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, GPIO_1_M2F_c
         => GPIO_1_M2F_c, GPIO_0_M2F_c => GPIO_0_M2F_c, N_23_i_0
         => N_23_i_0, FIC_0_LOCK => FIC_0_LOCK, 
        sha256_system_sb_0_FIC_0_CLK => 
        \sha256_system_sb_0_FIC_0_CLK\);
    
    FABOSC_0 : sha256_system_sb_FABOSC_0_OSC
      port map(FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
         => FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    CORERESETP_0 : CoreResetP
      port map(MSS_READY => MSS_READY, 
        sha256_system_sb_0_FIC_0_CLK => 
        \sha256_system_sb_0_FIC_0_CLK\, 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        sha256_system_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        sha256_system_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        sha256_system_sb_0_POWER_ON_RESET_N => 
        \sha256_system_sb_0_POWER_ON_RESET_N\);
    
    CoreAHBLite_0 : CoreAHBLite
      port map(
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        arbRegSMCurrentState(15) => arbRegSMCurrentState(15), 
        arbRegSMCurrentState_ns_i_0_0_0_a0_0(1) => 
        \arbRegSMCurrentState_ns_i_0_0_0_a0_0[1]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        masterAddrInProg(3) => masterAddrInProg(3), 
        masterAddrInProg(2) => masterAddrInProg(2), 
        masterAddrInProg(1) => masterAddrInProg(1), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0) => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        AHB_slave_dummy_0_mem_wdata(31) => 
        AHB_slave_dummy_0_mem_wdata(31), 
        AHB_slave_dummy_0_mem_wdata(30) => 
        AHB_slave_dummy_0_mem_wdata(30), 
        AHB_slave_dummy_0_mem_wdata(29) => 
        AHB_slave_dummy_0_mem_wdata(29), 
        AHB_slave_dummy_0_mem_wdata(28) => 
        AHB_slave_dummy_0_mem_wdata(28), 
        AHB_slave_dummy_0_mem_wdata(27) => 
        AHB_slave_dummy_0_mem_wdata(27), 
        AHB_slave_dummy_0_mem_wdata(26) => 
        AHB_slave_dummy_0_mem_wdata(26), 
        AHB_slave_dummy_0_mem_wdata(25) => 
        AHB_slave_dummy_0_mem_wdata(25), 
        AHB_slave_dummy_0_mem_wdata(24) => 
        AHB_slave_dummy_0_mem_wdata(24), 
        AHB_slave_dummy_0_mem_wdata(23) => 
        AHB_slave_dummy_0_mem_wdata(23), 
        AHB_slave_dummy_0_mem_wdata(22) => 
        AHB_slave_dummy_0_mem_wdata(22), 
        AHB_slave_dummy_0_mem_wdata(21) => 
        AHB_slave_dummy_0_mem_wdata(21), 
        AHB_slave_dummy_0_mem_wdata(20) => 
        AHB_slave_dummy_0_mem_wdata(20), 
        AHB_slave_dummy_0_mem_wdata(19) => 
        AHB_slave_dummy_0_mem_wdata(19), 
        AHB_slave_dummy_0_mem_wdata(18) => 
        AHB_slave_dummy_0_mem_wdata(18), 
        AHB_slave_dummy_0_mem_wdata(17) => 
        AHB_slave_dummy_0_mem_wdata(17), 
        AHB_slave_dummy_0_mem_wdata(16) => 
        AHB_slave_dummy_0_mem_wdata(16), 
        AHB_slave_dummy_0_mem_wdata(15) => 
        AHB_slave_dummy_0_mem_wdata(15), 
        AHB_slave_dummy_0_mem_wdata(14) => 
        AHB_slave_dummy_0_mem_wdata(14), 
        AHB_slave_dummy_0_mem_wdata(13) => 
        AHB_slave_dummy_0_mem_wdata(13), 
        AHB_slave_dummy_0_mem_wdata(12) => 
        AHB_slave_dummy_0_mem_wdata(12), 
        AHB_slave_dummy_0_mem_wdata(11) => 
        AHB_slave_dummy_0_mem_wdata(11), 
        AHB_slave_dummy_0_mem_wdata(10) => 
        AHB_slave_dummy_0_mem_wdata(10), 
        AHB_slave_dummy_0_mem_wdata(9) => 
        AHB_slave_dummy_0_mem_wdata(9), 
        AHB_slave_dummy_0_mem_wdata(8) => 
        AHB_slave_dummy_0_mem_wdata(8), 
        AHB_slave_dummy_0_mem_wdata(7) => 
        AHB_slave_dummy_0_mem_wdata(7), 
        AHB_slave_dummy_0_mem_wdata(6) => 
        AHB_slave_dummy_0_mem_wdata(6), 
        AHB_slave_dummy_0_mem_wdata(5) => 
        AHB_slave_dummy_0_mem_wdata(5), 
        AHB_slave_dummy_0_mem_wdata(4) => 
        AHB_slave_dummy_0_mem_wdata(4), 
        AHB_slave_dummy_0_mem_wdata(3) => 
        AHB_slave_dummy_0_mem_wdata(3), 
        AHB_slave_dummy_0_mem_wdata(2) => 
        AHB_slave_dummy_0_mem_wdata(2), 
        AHB_slave_dummy_0_mem_wdata(1) => 
        AHB_slave_dummy_0_mem_wdata(1), 
        AHB_slave_dummy_0_mem_wdata(0) => 
        AHB_slave_dummy_0_mem_wdata(0), 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3 => 
        \sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22, 
        MSS_READY => MSS_READY, sha256_system_sb_0_FIC_0_CLK => 
        \sha256_system_sb_0_FIC_0_CLK\, regHWRITE => regHWRITE, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE => 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        regHTRANS => regHTRANS, masterRegAddrSel => 
        \masterRegAddrSel\, N_358 => N_358, N_401 => N_401, N_403
         => N_403, sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, N_208 => N_208, 
        N_211 => N_211, N_354 => N_354, N_355 => N_355, N_395 => 
        N_395, hready_m_xhdl339 => hready_m_xhdl339, N_23_i_0 => 
        N_23_i_0, N_359 => N_359, N_253 => N_253, N_344 => N_344, 
        N_321_2 => N_321_2, N_36_2 => N_36_2, N_48_i_0 => 
        N_48_i_0, N_46_i_0 => N_46_i_0, N_44_i_0 => N_44_i_0, 
        N_42_i_0 => N_42_i_0, N_16_i_0 => N_16_i_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    SYSRESET_POR_RNI03O8 : CLKINT
      port map(A => \SYSRESET_POR\, Y => 
        \sha256_system_sb_0_POWER_ON_RESET_N\);
    
    CCC_0 : sha256_system_sb_CCC_0_FCCC
      port map(sha256_system_sb_0_FIC_0_CLK => 
        \sha256_system_sb_0_FIC_0_CLK\, FIC_0_LOCK => FIC_0_LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => \SYSRESET_POR\, DEVRST_N => 
        DEVRST_N);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_system is

    port( DEVRST_N   : in    std_logic;
          GPIO_0_M2F : out   std_logic;
          GPIO_1_M2F : out   std_logic;
          GPIO_2_M2F : out   std_logic
        );

end sha256_system;

architecture DEF_ARCH of sha256_system is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component reg_8x32
    port( raddr_in_net_0                      : in    std_logic_vector(3 downto 0) := (others => 'U');
          waddr_in_net_0                      : in    std_logic_vector(3 downto 0) := (others => 'U');
          AHB_slave_dummy_0_mem_wdata         : in    std_logic_vector(31 downto 0) := (others => 'U');
          data_out_9_0_29                     : out   std_logic;
          data_out_9_0_1                      : out   std_logic;
          data_out_9_0_0                      : out   std_logic;
          data_out_9_0_31                     : out   std_logic;
          sha256_system_sb_0_FIC_0_CLK        : in    std_logic := 'U';
          sha256_system_sb_0_POWER_ON_RESET_N : in    std_logic := 'U';
          N_1323                              : out   std_logic;
          N_1328                              : out   std_logic;
          N_1330                              : out   std_logic;
          N_1331                              : out   std_logic;
          N_1332                              : out   std_logic;
          N_1324                              : out   std_logic;
          N_1325                              : out   std_logic;
          N_1326                              : out   std_logic;
          N_1329                              : out   std_logic;
          N_1333                              : out   std_logic;
          N_1334                              : out   std_logic;
          N_1335                              : out   std_logic;
          N_1336                              : out   std_logic;
          N_1337                              : out   std_logic;
          N_1338                              : out   std_logic;
          N_1339                              : out   std_logic;
          N_1340                              : out   std_logic;
          N_1341                              : out   std_logic;
          N_1342                              : out   std_logic;
          N_1343                              : out   std_logic;
          N_1344                              : out   std_logic;
          N_1345                              : out   std_logic;
          N_1327                              : out   std_logic;
          N_1346                              : out   std_logic;
          N_1347                              : out   std_logic;
          N_1348                              : out   std_logic;
          N_1349                              : out   std_logic;
          N_1351                              : out   std_logic;
          N_1270                              : out   std_logic;
          N_1256                              : out   std_logic;
          N_1261                              : out   std_logic;
          N_1263                              : out   std_logic;
          N_1265                              : out   std_logic;
          N_1257                              : out   std_logic;
          N_1258                              : out   std_logic;
          N_1259                              : out   std_logic;
          N_1262                              : out   std_logic;
          N_1264                              : out   std_logic;
          N_1266                              : out   std_logic;
          N_1267                              : out   std_logic;
          N_1268                              : out   std_logic;
          N_1269                              : out   std_logic;
          N_1271                              : out   std_logic;
          N_1272                              : out   std_logic;
          N_1273                              : out   std_logic;
          N_1274                              : out   std_logic;
          N_1275                              : out   std_logic;
          N_1276                              : out   std_logic;
          N_1277                              : out   std_logic;
          N_1278                              : out   std_logic;
          N_1260                              : out   std_logic;
          N_1279                              : out   std_logic;
          N_1280                              : out   std_logic;
          N_1281                              : out   std_logic;
          N_1282                              : out   std_logic;
          N_1284                              : out   std_logic;
          AHB_slave_dummy_0_read_en           : in    std_logic := 'U';
          AHB_slave_dummy_0_write_en          : in    std_logic := 'U';
          N_1446                              : out   std_logic;
          N_53                                : out   std_logic;
          N_1458                              : out   std_logic;
          N_1457                              : out   std_logic;
          data_out_sn_N_12_mux                : out   std_logic;
          N_1423_3                            : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AHB_slave_dummy
    port( waddr_in_net_0                                     : out   std_logic_vector(3 downto 0);
          raddr_in_net_0                                     : out   std_logic_vector(3 downto 0);
          arbRegSMCurrentState                               : in    std_logic_vector(15 to 15) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR  : in    std_logic_vector(27 downto 24) := (others => 'U');
          masterAddrInProg                                   : in    std_logic_vector(3 downto 1) := (others => 'U');
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS : in    std_logic_vector(1 to 1) := (others => 'U');
          sha256_system_sb_0_POWER_ON_RESET_N                : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                       : in    std_logic := 'U';
          N_42_i_0                                           : in    std_logic := 'U';
          N_44_i_0                                           : in    std_logic := 'U';
          N_46_i_0                                           : in    std_logic := 'U';
          N_48_i_0                                           : in    std_logic := 'U';
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY             : out   std_logic;
          AHB_slave_dummy_0_write_en                         : out   std_logic;
          AHB_slave_dummy_0_read_en                          : out   std_logic;
          N_16_i_0                                           : in    std_logic := 'U';
          masterRegAddrSel                                   : in    std_logic := 'U';
          regHTRANS                                          : in    std_logic := 'U';
          N_359                                              : in    std_logic := 'U';
          N_344                                              : in    std_logic := 'U';
          N_253                                              : in    std_logic := 'U';
          N_321_2                                            : in    std_logic := 'U';
          N_354                                              : in    std_logic := 'U';
          N_355                                              : in    std_logic := 'U';
          N_358                                              : in    std_logic := 'U';
          N_211                                              : in    std_logic := 'U';
          N_395                                              : in    std_logic := 'U';
          N_403                                              : in    std_logic := 'U';
          N_401                                              : in    std_logic := 'U';
          N_208                                              : in    std_logic := 'U';
          regHWRITE                                          : in    std_logic := 'U';
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE : in    std_logic := 'U';
          N_36_2                                             : out   std_logic
        );
  end component;

  component sha256_system_sb
    port( sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : inout   std_logic_vector(1 to 1);
          arbRegSMCurrentState                                 : out   std_logic_vector(15 to 15);
          masterAddrInProg                                     : out   std_logic_vector(3 downto 1);
          AHB_slave_dummy_0_mem_wdata                          : out   std_logic_vector(31 downto 0);
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 : inout   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 : inout   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 : inout   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 : inout   std_logic;
          data_out_9_0_29                                      : in    std_logic := 'U';
          data_out_9_0_31                                      : in    std_logic := 'U';
          data_out_9_0_1                                       : in    std_logic := 'U';
          data_out_9_0_0                                       : in    std_logic := 'U';
          sha256_system_sb_0_POWER_ON_RESET_N                  : out   std_logic;
          DEVRST_N                                             : in    std_logic := 'U';
          sha256_system_sb_0_FIC_0_CLK                         : out   std_logic;
          regHWRITE                                            : out   std_logic;
          sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : inout   std_logic;
          regHTRANS                                            : out   std_logic;
          masterRegAddrSel                                     : out   std_logic;
          N_358                                                : out   std_logic;
          N_401                                                : out   std_logic;
          N_403                                                : out   std_logic;
          sha256_system_sb_0_AMBA_SLAVE_0_HREADY               : in    std_logic := 'U';
          N_208                                                : out   std_logic;
          N_211                                                : out   std_logic;
          N_354                                                : out   std_logic;
          N_355                                                : out   std_logic;
          N_395                                                : out   std_logic;
          N_359                                                : out   std_logic;
          N_253                                                : out   std_logic;
          N_344                                                : out   std_logic;
          N_321_2                                              : out   std_logic;
          N_36_2                                               : in    std_logic := 'U';
          N_48_i_0                                             : out   std_logic;
          N_46_i_0                                             : out   std_logic;
          N_44_i_0                                             : out   std_logic;
          N_42_i_0                                             : out   std_logic;
          N_16_i_0                                             : out   std_logic;
          N_1256                                               : in    std_logic := 'U';
          data_out_sn_N_12_mux                                 : in    std_logic := 'U';
          N_1323                                               : in    std_logic := 'U';
          N_1257                                               : in    std_logic := 'U';
          N_1324                                               : in    std_logic := 'U';
          N_1258                                               : in    std_logic := 'U';
          N_1325                                               : in    std_logic := 'U';
          N_1259                                               : in    std_logic := 'U';
          N_1326                                               : in    std_logic := 'U';
          N_1260                                               : in    std_logic := 'U';
          N_1327                                               : in    std_logic := 'U';
          N_1261                                               : in    std_logic := 'U';
          N_1328                                               : in    std_logic := 'U';
          N_1262                                               : in    std_logic := 'U';
          N_1329                                               : in    std_logic := 'U';
          N_1263                                               : in    std_logic := 'U';
          N_1330                                               : in    std_logic := 'U';
          N_1264                                               : in    std_logic := 'U';
          N_1331                                               : in    std_logic := 'U';
          N_1265                                               : in    std_logic := 'U';
          N_1332                                               : in    std_logic := 'U';
          N_1266                                               : in    std_logic := 'U';
          N_1333                                               : in    std_logic := 'U';
          N_1267                                               : in    std_logic := 'U';
          N_1334                                               : in    std_logic := 'U';
          N_1268                                               : in    std_logic := 'U';
          N_1335                                               : in    std_logic := 'U';
          N_1269                                               : in    std_logic := 'U';
          N_1336                                               : in    std_logic := 'U';
          N_1270                                               : in    std_logic := 'U';
          N_1337                                               : in    std_logic := 'U';
          N_1271                                               : in    std_logic := 'U';
          N_1338                                               : in    std_logic := 'U';
          N_1272                                               : in    std_logic := 'U';
          N_1339                                               : in    std_logic := 'U';
          N_1273                                               : in    std_logic := 'U';
          N_1340                                               : in    std_logic := 'U';
          N_1274                                               : in    std_logic := 'U';
          N_1341                                               : in    std_logic := 'U';
          N_1275                                               : in    std_logic := 'U';
          N_1342                                               : in    std_logic := 'U';
          N_1276                                               : in    std_logic := 'U';
          N_1343                                               : in    std_logic := 'U';
          N_1277                                               : in    std_logic := 'U';
          N_1344                                               : in    std_logic := 'U';
          N_1278                                               : in    std_logic := 'U';
          N_1345                                               : in    std_logic := 'U';
          N_1279                                               : in    std_logic := 'U';
          N_1346                                               : in    std_logic := 'U';
          N_1280                                               : in    std_logic := 'U';
          N_1347                                               : in    std_logic := 'U';
          N_1281                                               : in    std_logic := 'U';
          N_1348                                               : in    std_logic := 'U';
          N_1282                                               : in    std_logic := 'U';
          N_1349                                               : in    std_logic := 'U';
          N_1284                                               : in    std_logic := 'U';
          N_1351                                               : in    std_logic := 'U';
          N_1446                                               : in    std_logic := 'U';
          N_1423_3                                             : in    std_logic := 'U';
          N_53                                                 : in    std_logic := 'U';
          N_1457                                               : in    std_logic := 'U';
          N_1458                                               : in    std_logic := 'U';
          GPIO_2_M2F_c                                         : out   std_logic;
          GPIO_1_M2F_c                                         : out   std_logic;
          GPIO_0_M2F_c                                         : out   std_logic
        );
  end component;

    signal sha256_system_sb_0_FIC_0_CLK, 
        sha256_system_sb_0_POWER_ON_RESET_N, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, 
        \waddr_in_net_0[0]\, \waddr_in_net_0[1]\, 
        \waddr_in_net_0[2]\, \waddr_in_net_0[3]\, 
        \raddr_in_net_0[0]\, \raddr_in_net_0[1]\, 
        \raddr_in_net_0[2]\, \raddr_in_net_0[3]\, 
        AHB_slave_dummy_0_write_en, AHB_slave_dummy_0_read_en, 
        GND_net_1, VCC_net_1, 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[24]\, 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[25]\, 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[26]\, 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[27]\, 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.masterAddrInProg[1]\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.masterAddrInProg[2]\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.masterAddrInProg[3]\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.masterRegAddrSel\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.regHTRANS\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.regHWRITE\, 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.slave_arbiter.arbRegSMCurrentState[15]\, 
        GPIO_0_M2F_c, GPIO_1_M2F_c, GPIO_2_M2F_c, 
        \AHB_slave_dummy_0_mem_wdata[0]\, 
        \AHB_slave_dummy_0_mem_wdata[1]\, 
        \reg_2x32_0.data_out_sn_N_12_mux\, \reg_2x32_0.N_1423_3\, 
        \reg_2x32_0.N_1457\, \reg_2x32_0.N_1458\, 
        \AHB_slave_dummy_0_mem_wdata[29]\, 
        \AHB_slave_dummy_0_mem_wdata[22]\, \reg_2x32_0.N_53\, 
        \AHB_slave_dummy_0_mem_wdata[31]\, N_359, N_36_2, N_253, 
        N_403, N_401, N_344, N_358, N_354, N_355, N_208, N_395, 
        N_211, \AHB_slave_dummy_0_mem_wdata[2]\, 
        \AHB_slave_dummy_0_mem_wdata[3]\, 
        \AHB_slave_dummy_0_mem_wdata[4]\, 
        \AHB_slave_dummy_0_mem_wdata[5]\, 
        \AHB_slave_dummy_0_mem_wdata[6]\, 
        \AHB_slave_dummy_0_mem_wdata[7]\, 
        \AHB_slave_dummy_0_mem_wdata[8]\, 
        \AHB_slave_dummy_0_mem_wdata[9]\, 
        \AHB_slave_dummy_0_mem_wdata[10]\, 
        \AHB_slave_dummy_0_mem_wdata[11]\, 
        \AHB_slave_dummy_0_mem_wdata[12]\, 
        \AHB_slave_dummy_0_mem_wdata[13]\, 
        \AHB_slave_dummy_0_mem_wdata[14]\, 
        \AHB_slave_dummy_0_mem_wdata[15]\, 
        \AHB_slave_dummy_0_mem_wdata[16]\, 
        \AHB_slave_dummy_0_mem_wdata[17]\, 
        \AHB_slave_dummy_0_mem_wdata[18]\, 
        \AHB_slave_dummy_0_mem_wdata[19]\, 
        \AHB_slave_dummy_0_mem_wdata[20]\, 
        \AHB_slave_dummy_0_mem_wdata[21]\, 
        \AHB_slave_dummy_0_mem_wdata[23]\, 
        \AHB_slave_dummy_0_mem_wdata[24]\, 
        \AHB_slave_dummy_0_mem_wdata[25]\, 
        \AHB_slave_dummy_0_mem_wdata[26]\, 
        \AHB_slave_dummy_0_mem_wdata[27]\, 
        \AHB_slave_dummy_0_mem_wdata[28]\, 
        \AHB_slave_dummy_0_mem_wdata[30]\, \reg_2x32_0.N_1270\, 
        \reg_2x32_0.N_1256\, \reg_2x32_0.N_1261\, 
        \reg_2x32_0.N_1323\, \reg_2x32_0.N_1328\, 
        \reg_2x32_0.N_1263\, \reg_2x32_0.N_1330\, 
        \reg_2x32_0.N_1331\, \reg_2x32_0.N_1265\, 
        \reg_2x32_0.N_1332\, \reg_2x32_0.N_1257\, 
        \reg_2x32_0.N_1324\, \reg_2x32_0.N_1258\, 
        \reg_2x32_0.N_1325\, \reg_2x32_0.N_1259\, 
        \reg_2x32_0.N_1326\, \reg_2x32_0.N_1262\, 
        \reg_2x32_0.N_1329\, \reg_2x32_0.N_1264\, 
        \reg_2x32_0.N_1266\, \reg_2x32_0.N_1333\, 
        \reg_2x32_0.N_1267\, \reg_2x32_0.N_1334\, 
        \reg_2x32_0.N_1268\, \reg_2x32_0.N_1335\, 
        \reg_2x32_0.N_1269\, \reg_2x32_0.N_1336\, 
        \reg_2x32_0.N_1337\, \reg_2x32_0.N_1271\, 
        \reg_2x32_0.N_1338\, \reg_2x32_0.N_1272\, 
        \reg_2x32_0.N_1339\, \reg_2x32_0.N_1273\, 
        \reg_2x32_0.N_1340\, \reg_2x32_0.N_1274\, 
        \reg_2x32_0.N_1341\, \reg_2x32_0.N_1275\, 
        \reg_2x32_0.N_1342\, \reg_2x32_0.N_1276\, 
        \reg_2x32_0.N_1343\, \reg_2x32_0.N_1277\, 
        \reg_2x32_0.N_1344\, \reg_2x32_0.N_1278\, 
        \reg_2x32_0.N_1345\, \reg_2x32_0.N_1260\, 
        \reg_2x32_0.N_1279\, \reg_2x32_0.N_1327\, 
        \reg_2x32_0.N_1346\, \reg_2x32_0.N_1280\, 
        \reg_2x32_0.N_1347\, \reg_2x32_0.N_1281\, 
        \reg_2x32_0.N_1282\, \reg_2x32_0.N_1348\, 
        \reg_2x32_0.N_1349\, \reg_2x32_0.N_1446\, 
        \reg_2x32_0.N_1284\, \reg_2x32_0.N_1351\, N_321_2, 
        \reg_2x32_0.data_out_9_0[31]\, 
        \reg_2x32_0.data_out_9_0[0]\, 
        \reg_2x32_0.data_out_9_0[1]\, 
        \reg_2x32_0.data_out_9_0[29]\, N_16_i_0, N_48_i_0, 
        N_46_i_0, N_44_i_0, N_42_i_0 : std_logic;

    for all : reg_8x32
	Use entity work.reg_8x32(DEF_ARCH);
    for all : AHB_slave_dummy
	Use entity work.AHB_slave_dummy(DEF_ARCH);
    for all : sha256_system_sb
	Use entity work.sha256_system_sb(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    GPIO_2_M2F_obuf : OUTBUF
      port map(D => GPIO_2_M2F_c, PAD => GPIO_2_M2F);
    
    reg_2x32_0 : reg_8x32
      port map(raddr_in_net_0(3) => \raddr_in_net_0[3]\, 
        raddr_in_net_0(2) => \raddr_in_net_0[2]\, 
        raddr_in_net_0(1) => \raddr_in_net_0[1]\, 
        raddr_in_net_0(0) => \raddr_in_net_0[0]\, 
        waddr_in_net_0(3) => \waddr_in_net_0[3]\, 
        waddr_in_net_0(2) => \waddr_in_net_0[2]\, 
        waddr_in_net_0(1) => \waddr_in_net_0[1]\, 
        waddr_in_net_0(0) => \waddr_in_net_0[0]\, 
        AHB_slave_dummy_0_mem_wdata(31) => 
        \AHB_slave_dummy_0_mem_wdata[31]\, 
        AHB_slave_dummy_0_mem_wdata(30) => 
        \AHB_slave_dummy_0_mem_wdata[30]\, 
        AHB_slave_dummy_0_mem_wdata(29) => 
        \AHB_slave_dummy_0_mem_wdata[29]\, 
        AHB_slave_dummy_0_mem_wdata(28) => 
        \AHB_slave_dummy_0_mem_wdata[28]\, 
        AHB_slave_dummy_0_mem_wdata(27) => 
        \AHB_slave_dummy_0_mem_wdata[27]\, 
        AHB_slave_dummy_0_mem_wdata(26) => 
        \AHB_slave_dummy_0_mem_wdata[26]\, 
        AHB_slave_dummy_0_mem_wdata(25) => 
        \AHB_slave_dummy_0_mem_wdata[25]\, 
        AHB_slave_dummy_0_mem_wdata(24) => 
        \AHB_slave_dummy_0_mem_wdata[24]\, 
        AHB_slave_dummy_0_mem_wdata(23) => 
        \AHB_slave_dummy_0_mem_wdata[23]\, 
        AHB_slave_dummy_0_mem_wdata(22) => 
        \AHB_slave_dummy_0_mem_wdata[22]\, 
        AHB_slave_dummy_0_mem_wdata(21) => 
        \AHB_slave_dummy_0_mem_wdata[21]\, 
        AHB_slave_dummy_0_mem_wdata(20) => 
        \AHB_slave_dummy_0_mem_wdata[20]\, 
        AHB_slave_dummy_0_mem_wdata(19) => 
        \AHB_slave_dummy_0_mem_wdata[19]\, 
        AHB_slave_dummy_0_mem_wdata(18) => 
        \AHB_slave_dummy_0_mem_wdata[18]\, 
        AHB_slave_dummy_0_mem_wdata(17) => 
        \AHB_slave_dummy_0_mem_wdata[17]\, 
        AHB_slave_dummy_0_mem_wdata(16) => 
        \AHB_slave_dummy_0_mem_wdata[16]\, 
        AHB_slave_dummy_0_mem_wdata(15) => 
        \AHB_slave_dummy_0_mem_wdata[15]\, 
        AHB_slave_dummy_0_mem_wdata(14) => 
        \AHB_slave_dummy_0_mem_wdata[14]\, 
        AHB_slave_dummy_0_mem_wdata(13) => 
        \AHB_slave_dummy_0_mem_wdata[13]\, 
        AHB_slave_dummy_0_mem_wdata(12) => 
        \AHB_slave_dummy_0_mem_wdata[12]\, 
        AHB_slave_dummy_0_mem_wdata(11) => 
        \AHB_slave_dummy_0_mem_wdata[11]\, 
        AHB_slave_dummy_0_mem_wdata(10) => 
        \AHB_slave_dummy_0_mem_wdata[10]\, 
        AHB_slave_dummy_0_mem_wdata(9) => 
        \AHB_slave_dummy_0_mem_wdata[9]\, 
        AHB_slave_dummy_0_mem_wdata(8) => 
        \AHB_slave_dummy_0_mem_wdata[8]\, 
        AHB_slave_dummy_0_mem_wdata(7) => 
        \AHB_slave_dummy_0_mem_wdata[7]\, 
        AHB_slave_dummy_0_mem_wdata(6) => 
        \AHB_slave_dummy_0_mem_wdata[6]\, 
        AHB_slave_dummy_0_mem_wdata(5) => 
        \AHB_slave_dummy_0_mem_wdata[5]\, 
        AHB_slave_dummy_0_mem_wdata(4) => 
        \AHB_slave_dummy_0_mem_wdata[4]\, 
        AHB_slave_dummy_0_mem_wdata(3) => 
        \AHB_slave_dummy_0_mem_wdata[3]\, 
        AHB_slave_dummy_0_mem_wdata(2) => 
        \AHB_slave_dummy_0_mem_wdata[2]\, 
        AHB_slave_dummy_0_mem_wdata(1) => 
        \AHB_slave_dummy_0_mem_wdata[1]\, 
        AHB_slave_dummy_0_mem_wdata(0) => 
        \AHB_slave_dummy_0_mem_wdata[0]\, data_out_9_0_29 => 
        \reg_2x32_0.data_out_9_0[29]\, data_out_9_0_1 => 
        \reg_2x32_0.data_out_9_0[1]\, data_out_9_0_0 => 
        \reg_2x32_0.data_out_9_0[0]\, data_out_9_0_31 => 
        \reg_2x32_0.data_out_9_0[31]\, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, 
        sha256_system_sb_0_POWER_ON_RESET_N => 
        sha256_system_sb_0_POWER_ON_RESET_N, N_1323 => 
        \reg_2x32_0.N_1323\, N_1328 => \reg_2x32_0.N_1328\, 
        N_1330 => \reg_2x32_0.N_1330\, N_1331 => 
        \reg_2x32_0.N_1331\, N_1332 => \reg_2x32_0.N_1332\, 
        N_1324 => \reg_2x32_0.N_1324\, N_1325 => 
        \reg_2x32_0.N_1325\, N_1326 => \reg_2x32_0.N_1326\, 
        N_1329 => \reg_2x32_0.N_1329\, N_1333 => 
        \reg_2x32_0.N_1333\, N_1334 => \reg_2x32_0.N_1334\, 
        N_1335 => \reg_2x32_0.N_1335\, N_1336 => 
        \reg_2x32_0.N_1336\, N_1337 => \reg_2x32_0.N_1337\, 
        N_1338 => \reg_2x32_0.N_1338\, N_1339 => 
        \reg_2x32_0.N_1339\, N_1340 => \reg_2x32_0.N_1340\, 
        N_1341 => \reg_2x32_0.N_1341\, N_1342 => 
        \reg_2x32_0.N_1342\, N_1343 => \reg_2x32_0.N_1343\, 
        N_1344 => \reg_2x32_0.N_1344\, N_1345 => 
        \reg_2x32_0.N_1345\, N_1327 => \reg_2x32_0.N_1327\, 
        N_1346 => \reg_2x32_0.N_1346\, N_1347 => 
        \reg_2x32_0.N_1347\, N_1348 => \reg_2x32_0.N_1348\, 
        N_1349 => \reg_2x32_0.N_1349\, N_1351 => 
        \reg_2x32_0.N_1351\, N_1270 => \reg_2x32_0.N_1270\, 
        N_1256 => \reg_2x32_0.N_1256\, N_1261 => 
        \reg_2x32_0.N_1261\, N_1263 => \reg_2x32_0.N_1263\, 
        N_1265 => \reg_2x32_0.N_1265\, N_1257 => 
        \reg_2x32_0.N_1257\, N_1258 => \reg_2x32_0.N_1258\, 
        N_1259 => \reg_2x32_0.N_1259\, N_1262 => 
        \reg_2x32_0.N_1262\, N_1264 => \reg_2x32_0.N_1264\, 
        N_1266 => \reg_2x32_0.N_1266\, N_1267 => 
        \reg_2x32_0.N_1267\, N_1268 => \reg_2x32_0.N_1268\, 
        N_1269 => \reg_2x32_0.N_1269\, N_1271 => 
        \reg_2x32_0.N_1271\, N_1272 => \reg_2x32_0.N_1272\, 
        N_1273 => \reg_2x32_0.N_1273\, N_1274 => 
        \reg_2x32_0.N_1274\, N_1275 => \reg_2x32_0.N_1275\, 
        N_1276 => \reg_2x32_0.N_1276\, N_1277 => 
        \reg_2x32_0.N_1277\, N_1278 => \reg_2x32_0.N_1278\, 
        N_1260 => \reg_2x32_0.N_1260\, N_1279 => 
        \reg_2x32_0.N_1279\, N_1280 => \reg_2x32_0.N_1280\, 
        N_1281 => \reg_2x32_0.N_1281\, N_1282 => 
        \reg_2x32_0.N_1282\, N_1284 => \reg_2x32_0.N_1284\, 
        AHB_slave_dummy_0_read_en => AHB_slave_dummy_0_read_en, 
        AHB_slave_dummy_0_write_en => AHB_slave_dummy_0_write_en, 
        N_1446 => \reg_2x32_0.N_1446\, N_53 => \reg_2x32_0.N_53\, 
        N_1458 => \reg_2x32_0.N_1458\, N_1457 => 
        \reg_2x32_0.N_1457\, data_out_sn_N_12_mux => 
        \reg_2x32_0.data_out_sn_N_12_mux\, N_1423_3 => 
        \reg_2x32_0.N_1423_3\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    AHB_slave_dummy_0 : AHB_slave_dummy
      port map(waddr_in_net_0(3) => \waddr_in_net_0[3]\, 
        waddr_in_net_0(2) => \waddr_in_net_0[2]\, 
        waddr_in_net_0(1) => \waddr_in_net_0[1]\, 
        waddr_in_net_0(0) => \waddr_in_net_0[0]\, 
        raddr_in_net_0(3) => \raddr_in_net_0[3]\, 
        raddr_in_net_0(2) => \raddr_in_net_0[2]\, 
        raddr_in_net_0(1) => \raddr_in_net_0[1]\, 
        raddr_in_net_0(0) => \raddr_in_net_0[0]\, 
        arbRegSMCurrentState(15) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.slave_arbiter.arbRegSMCurrentState[15]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(27) => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[27]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(26) => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[26]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(25) => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[25]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(24) => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[24]\, 
        masterAddrInProg(3) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.masterAddrInProg[3]\, 
        masterAddrInProg(2) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.masterAddrInProg[2]\, 
        masterAddrInProg(1) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.masterAddrInProg[1]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        sha256_system_sb_0_POWER_ON_RESET_N => 
        sha256_system_sb_0_POWER_ON_RESET_N, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, N_42_i_0 => N_42_i_0, 
        N_44_i_0 => N_44_i_0, N_46_i_0 => N_46_i_0, N_48_i_0 => 
        N_48_i_0, sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, 
        AHB_slave_dummy_0_write_en => AHB_slave_dummy_0_write_en, 
        AHB_slave_dummy_0_read_en => AHB_slave_dummy_0_read_en, 
        N_16_i_0 => N_16_i_0, masterRegAddrSel => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.masterRegAddrSel\, 
        regHTRANS => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.regHTRANS\, 
        N_359 => N_359, N_344 => N_344, N_253 => N_253, N_321_2
         => N_321_2, N_354 => N_354, N_355 => N_355, N_358 => 
        N_358, N_211 => N_211, N_395 => N_395, N_403 => N_403, 
        N_401 => N_401, N_208 => N_208, regHWRITE => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.regHWRITE\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE\, 
        N_36_2 => N_36_2);
    
    GPIO_1_M2F_obuf : OUTBUF
      port map(D => GPIO_1_M2F_c, PAD => GPIO_1_M2F);
    
    sha256_system_sb_0 : sha256_system_sb
      port map(
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1) => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        arbRegSMCurrentState(15) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.slave_arbiter.arbRegSMCurrentState[15]\, 
        masterAddrInProg(3) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.masterAddrInProg[3]\, 
        masterAddrInProg(2) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.masterAddrInProg[2]\, 
        masterAddrInProg(1) => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.slavestage_0.masterAddrInProg[1]\, 
        AHB_slave_dummy_0_mem_wdata(31) => 
        \AHB_slave_dummy_0_mem_wdata[31]\, 
        AHB_slave_dummy_0_mem_wdata(30) => 
        \AHB_slave_dummy_0_mem_wdata[30]\, 
        AHB_slave_dummy_0_mem_wdata(29) => 
        \AHB_slave_dummy_0_mem_wdata[29]\, 
        AHB_slave_dummy_0_mem_wdata(28) => 
        \AHB_slave_dummy_0_mem_wdata[28]\, 
        AHB_slave_dummy_0_mem_wdata(27) => 
        \AHB_slave_dummy_0_mem_wdata[27]\, 
        AHB_slave_dummy_0_mem_wdata(26) => 
        \AHB_slave_dummy_0_mem_wdata[26]\, 
        AHB_slave_dummy_0_mem_wdata(25) => 
        \AHB_slave_dummy_0_mem_wdata[25]\, 
        AHB_slave_dummy_0_mem_wdata(24) => 
        \AHB_slave_dummy_0_mem_wdata[24]\, 
        AHB_slave_dummy_0_mem_wdata(23) => 
        \AHB_slave_dummy_0_mem_wdata[23]\, 
        AHB_slave_dummy_0_mem_wdata(22) => 
        \AHB_slave_dummy_0_mem_wdata[22]\, 
        AHB_slave_dummy_0_mem_wdata(21) => 
        \AHB_slave_dummy_0_mem_wdata[21]\, 
        AHB_slave_dummy_0_mem_wdata(20) => 
        \AHB_slave_dummy_0_mem_wdata[20]\, 
        AHB_slave_dummy_0_mem_wdata(19) => 
        \AHB_slave_dummy_0_mem_wdata[19]\, 
        AHB_slave_dummy_0_mem_wdata(18) => 
        \AHB_slave_dummy_0_mem_wdata[18]\, 
        AHB_slave_dummy_0_mem_wdata(17) => 
        \AHB_slave_dummy_0_mem_wdata[17]\, 
        AHB_slave_dummy_0_mem_wdata(16) => 
        \AHB_slave_dummy_0_mem_wdata[16]\, 
        AHB_slave_dummy_0_mem_wdata(15) => 
        \AHB_slave_dummy_0_mem_wdata[15]\, 
        AHB_slave_dummy_0_mem_wdata(14) => 
        \AHB_slave_dummy_0_mem_wdata[14]\, 
        AHB_slave_dummy_0_mem_wdata(13) => 
        \AHB_slave_dummy_0_mem_wdata[13]\, 
        AHB_slave_dummy_0_mem_wdata(12) => 
        \AHB_slave_dummy_0_mem_wdata[12]\, 
        AHB_slave_dummy_0_mem_wdata(11) => 
        \AHB_slave_dummy_0_mem_wdata[11]\, 
        AHB_slave_dummy_0_mem_wdata(10) => 
        \AHB_slave_dummy_0_mem_wdata[10]\, 
        AHB_slave_dummy_0_mem_wdata(9) => 
        \AHB_slave_dummy_0_mem_wdata[9]\, 
        AHB_slave_dummy_0_mem_wdata(8) => 
        \AHB_slave_dummy_0_mem_wdata[8]\, 
        AHB_slave_dummy_0_mem_wdata(7) => 
        \AHB_slave_dummy_0_mem_wdata[7]\, 
        AHB_slave_dummy_0_mem_wdata(6) => 
        \AHB_slave_dummy_0_mem_wdata[6]\, 
        AHB_slave_dummy_0_mem_wdata(5) => 
        \AHB_slave_dummy_0_mem_wdata[5]\, 
        AHB_slave_dummy_0_mem_wdata(4) => 
        \AHB_slave_dummy_0_mem_wdata[4]\, 
        AHB_slave_dummy_0_mem_wdata(3) => 
        \AHB_slave_dummy_0_mem_wdata[3]\, 
        AHB_slave_dummy_0_mem_wdata(2) => 
        \AHB_slave_dummy_0_mem_wdata[2]\, 
        AHB_slave_dummy_0_mem_wdata(1) => 
        \AHB_slave_dummy_0_mem_wdata[1]\, 
        AHB_slave_dummy_0_mem_wdata(0) => 
        \AHB_slave_dummy_0_mem_wdata[0]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_25 => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[27]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_24 => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[26]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_23 => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[25]\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_22 => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[24]\, 
        data_out_9_0_29 => \reg_2x32_0.data_out_9_0[29]\, 
        data_out_9_0_31 => \reg_2x32_0.data_out_9_0[31]\, 
        data_out_9_0_1 => \reg_2x32_0.data_out_9_0[1]\, 
        data_out_9_0_0 => \reg_2x32_0.data_out_9_0[0]\, 
        sha256_system_sb_0_POWER_ON_RESET_N => 
        sha256_system_sb_0_POWER_ON_RESET_N, DEVRST_N => DEVRST_N, 
        sha256_system_sb_0_FIC_0_CLK => 
        sha256_system_sb_0_FIC_0_CLK, regHWRITE => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.regHWRITE\, 
        sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE => 
        \sha256_system_sb_0.sha256_system_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE\, 
        regHTRANS => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.regHTRANS\, 
        masterRegAddrSel => 
        \sha256_system_sb_0.CoreAHBLite_0.matrix4x16.masterstage_0.masterRegAddrSel\, 
        N_358 => N_358, N_401 => N_401, N_403 => N_403, 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY => 
        sha256_system_sb_0_AMBA_SLAVE_0_HREADY, N_208 => N_208, 
        N_211 => N_211, N_354 => N_354, N_355 => N_355, N_395 => 
        N_395, N_359 => N_359, N_253 => N_253, N_344 => N_344, 
        N_321_2 => N_321_2, N_36_2 => N_36_2, N_48_i_0 => 
        N_48_i_0, N_46_i_0 => N_46_i_0, N_44_i_0 => N_44_i_0, 
        N_42_i_0 => N_42_i_0, N_16_i_0 => N_16_i_0, N_1256 => 
        \reg_2x32_0.N_1256\, data_out_sn_N_12_mux => 
        \reg_2x32_0.data_out_sn_N_12_mux\, N_1323 => 
        \reg_2x32_0.N_1323\, N_1257 => \reg_2x32_0.N_1257\, 
        N_1324 => \reg_2x32_0.N_1324\, N_1258 => 
        \reg_2x32_0.N_1258\, N_1325 => \reg_2x32_0.N_1325\, 
        N_1259 => \reg_2x32_0.N_1259\, N_1326 => 
        \reg_2x32_0.N_1326\, N_1260 => \reg_2x32_0.N_1260\, 
        N_1327 => \reg_2x32_0.N_1327\, N_1261 => 
        \reg_2x32_0.N_1261\, N_1328 => \reg_2x32_0.N_1328\, 
        N_1262 => \reg_2x32_0.N_1262\, N_1329 => 
        \reg_2x32_0.N_1329\, N_1263 => \reg_2x32_0.N_1263\, 
        N_1330 => \reg_2x32_0.N_1330\, N_1264 => 
        \reg_2x32_0.N_1264\, N_1331 => \reg_2x32_0.N_1331\, 
        N_1265 => \reg_2x32_0.N_1265\, N_1332 => 
        \reg_2x32_0.N_1332\, N_1266 => \reg_2x32_0.N_1266\, 
        N_1333 => \reg_2x32_0.N_1333\, N_1267 => 
        \reg_2x32_0.N_1267\, N_1334 => \reg_2x32_0.N_1334\, 
        N_1268 => \reg_2x32_0.N_1268\, N_1335 => 
        \reg_2x32_0.N_1335\, N_1269 => \reg_2x32_0.N_1269\, 
        N_1336 => \reg_2x32_0.N_1336\, N_1270 => 
        \reg_2x32_0.N_1270\, N_1337 => \reg_2x32_0.N_1337\, 
        N_1271 => \reg_2x32_0.N_1271\, N_1338 => 
        \reg_2x32_0.N_1338\, N_1272 => \reg_2x32_0.N_1272\, 
        N_1339 => \reg_2x32_0.N_1339\, N_1273 => 
        \reg_2x32_0.N_1273\, N_1340 => \reg_2x32_0.N_1340\, 
        N_1274 => \reg_2x32_0.N_1274\, N_1341 => 
        \reg_2x32_0.N_1341\, N_1275 => \reg_2x32_0.N_1275\, 
        N_1342 => \reg_2x32_0.N_1342\, N_1276 => 
        \reg_2x32_0.N_1276\, N_1343 => \reg_2x32_0.N_1343\, 
        N_1277 => \reg_2x32_0.N_1277\, N_1344 => 
        \reg_2x32_0.N_1344\, N_1278 => \reg_2x32_0.N_1278\, 
        N_1345 => \reg_2x32_0.N_1345\, N_1279 => 
        \reg_2x32_0.N_1279\, N_1346 => \reg_2x32_0.N_1346\, 
        N_1280 => \reg_2x32_0.N_1280\, N_1347 => 
        \reg_2x32_0.N_1347\, N_1281 => \reg_2x32_0.N_1281\, 
        N_1348 => \reg_2x32_0.N_1348\, N_1282 => 
        \reg_2x32_0.N_1282\, N_1349 => \reg_2x32_0.N_1349\, 
        N_1284 => \reg_2x32_0.N_1284\, N_1351 => 
        \reg_2x32_0.N_1351\, N_1446 => \reg_2x32_0.N_1446\, 
        N_1423_3 => \reg_2x32_0.N_1423_3\, N_53 => 
        \reg_2x32_0.N_53\, N_1457 => \reg_2x32_0.N_1457\, N_1458
         => \reg_2x32_0.N_1458\, GPIO_2_M2F_c => GPIO_2_M2F_c, 
        GPIO_1_M2F_c => GPIO_1_M2F_c, GPIO_0_M2F_c => 
        GPIO_0_M2F_c);
    
    GPIO_0_M2F_obuf : OUTBUF
      port map(D => GPIO_0_M2F_c, PAD => GPIO_0_M2F);
    

end DEF_ARCH; 
