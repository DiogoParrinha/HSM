-- Version: v11.7 SP1 11.7.1.14

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_FABOSC_0_OSC is

    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );

end CertificationSystem_sb_FABOSC_0_OSC;

architecture DEF_ARCH of CertificationSystem_sb_FABOSC_0_OSC is 

  component RCOSC_25_50MHZ
    generic (FREQUENCY:real := 50.0);

    port( CLKOUT : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    I_RCOSC_25_50MHZ : RCOSC_25_50MHZ
      generic map(FREQUENCY => 50.0)

      port map(CLKOUT => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreResetP is

    port( MSS_READY                                             : out   std_logic;
          FAB_CCC_GL0                                           : in    std_logic;
          POWER_ON_RESET_N                                      : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic
        );

end CoreResetP;

architecture DEF_ARCH of CoreResetP is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \MSS_HPMS_READY_int\, \mss_ready_select\, VCC_net_1, 
        \POWER_ON_RESET_N_clk_base\, 
        \un6_fic_2_apb_m_preset_n_clk_base\, GND_net_1, 
        \mss_ready_state\, \RESET_N_M2F_clk_base\, 
        \POWER_ON_RESET_N_q1\, \RESET_N_M2F_q1\, 
        \FIC_2_APB_M_PRESET_N_q1\, 
        \FIC_2_APB_M_PRESET_N_clk_base\, \MSS_HPMS_READY_int_3\
         : std_logic;

begin 


    RESET_N_M2F_clk_base : SLE
      port map(D => \RESET_N_M2F_q1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RESET_N_M2F_clk_base\);
    
    POWER_ON_RESET_N_clk_base : SLE
      port map(D => \POWER_ON_RESET_N_q1\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \POWER_ON_RESET_N_clk_base\);
    
    mss_ready_select : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        \un6_fic_2_apb_m_preset_n_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_select\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    mss_ready_state : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        \RESET_N_M2F_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_state\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    un6_fic_2_apb_m_preset_n_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \FIC_2_APB_M_PRESET_N_clk_base\, B => 
        \mss_ready_state\, Y => 
        \un6_fic_2_apb_m_preset_n_clk_base\);
    
    RESET_N_M2F_q1 : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RESET_N_M2F_q1\);
    
    FIC_2_APB_M_PRESET_N_clk_base : SLE
      port map(D => \FIC_2_APB_M_PRESET_N_q1\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \FIC_2_APB_M_PRESET_N_clk_base\);
    
    POWER_ON_RESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => POWER_ON_RESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \POWER_ON_RESET_N_q1\);
    
    MSS_HPMS_READY_int_RNIRS5B : CLKINT
      port map(A => \MSS_HPMS_READY_int\, Y => MSS_READY);
    
    FIC_2_APB_M_PRESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \FIC_2_APB_M_PRESET_N_q1\);
    
    MSS_HPMS_READY_int_3 : CFG3
      generic map(INIT => x"E0")

      port map(A => \RESET_N_M2F_clk_base\, B => 
        \mss_ready_select\, C => \FIC_2_APB_M_PRESET_N_clk_base\, 
        Y => \MSS_HPMS_READY_int_3\);
    
    MSS_HPMS_READY_int : SLE
      port map(D => \MSS_HPMS_READY_int_3\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => \POWER_ON_RESET_N_clk_base\, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \MSS_HPMS_READY_int\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVEARBITER_1 is

    port( xhdl1221_i_0                                             : in    std_logic_vector(3 to 3);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS : in    std_logic_vector(1 to 1);
          MASTERADDRINPROG_i_a2_0_a3_d_d                           : out   std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_0                             : out   std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_1_0                           : out   std_logic_vector(0 to 0);
          sAddrDec                                                 : in    std_logic_vector(3 to 3);
          arbRegSMCurrentState_13                                  : out   std_logic;
          arbRegSMCurrentState_12                                  : out   std_logic;
          arbRegSMCurrentState_0                                   : out   std_logic;
          M0GATEDHADDR_2                                           : in    std_logic;
          M0GATEDHADDR_0                                           : in    std_logic;
          MSS_READY                                                : in    std_logic;
          FAB_CCC_GL0                                              : in    std_logic;
          regHTRANS                                                : in    std_logic;
          masterRegAddrSel                                         : in    std_logic;
          un3_saddrdec_i_a2_3_0                                    : in    std_logic;
          M0GATEDHTRANS                                            : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                      : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HSELx_i_1_i_0                   : out   std_logic;
          M0GATEDHWRITE                                            : in    std_logic;
          N_7_i_0                                                  : out   std_logic;
          N_25_i_0                                                 : out   std_logic
        );

end COREAHBLITE_SLAVEARBITER_1;

architecture DEF_ARCH of COREAHBLITE_SLAVEARBITER_1 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \arbRegSMCurrentState_13\, VCC_net_1, N_104_i_0, 
        GND_net_1, \arbRegSMCurrentState_12\, N_105, 
        \arbRegSMCurrentState_0\, N_89, 
        \arbRegSMCurrentState_ns_i_a2_1_o4_0[0]_net_1\, 
        \MASTERADDRINPROG_i_a2_0_a3_d_0[0]_net_1\, 
        \MASTERADDRINPROG_i_a2_0_a3_1_0[0]\ : std_logic;

begin 

    MASTERADDRINPROG_i_a2_0_a3_1_0(0) <= 
        \MASTERADDRINPROG_i_a2_0_a3_1_0[0]\;
    arbRegSMCurrentState_13 <= \arbRegSMCurrentState_13\;
    arbRegSMCurrentState_12 <= \arbRegSMCurrentState_12\;
    arbRegSMCurrentState_0 <= \arbRegSMCurrentState_0\;

    \arbRegSMCurrentState_ns_i_a2_1_o4_0_RNIRFNJ4[0]\ : CFG4
      generic map(INIT => x"4454")

      port map(A => CoreAHBLite_0_AHBmslave3_HREADY_i_1, B => 
        \arbRegSMCurrentState_13\, C => sAddrDec(3), D => 
        \arbRegSMCurrentState_ns_i_a2_1_o4_0[0]_net_1\, Y => 
        N_25_i_0);
    
    \arbRegSMCurrentState_ns_i_a2_1_o4_0_RNIKAUO[0]\ : CFG3
      generic map(INIT => x"F4")

      port map(A => 
        \arbRegSMCurrentState_ns_i_a2_1_o4_0[0]_net_1\, B => 
        sAddrDec(3), C => \arbRegSMCurrentState_13\, Y => 
        CoreAHBLite_0_AHBmslave3_HSELx_i_1_i_0);
    
    \arbRegSMCurrentState[15]\ : SLE
      port map(D => N_104_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_13\);
    
    \MASTERADDRINPROG_i_a2_0_a3_d_0[0]\ : CFG4
      generic map(INIT => x"5155")

      port map(A => \arbRegSMCurrentState_13\, B => 
        un3_saddrdec_i_a2_3_0, C => M0GATEDHADDR_2, D => 
        M0GATEDHADDR_0, Y => 
        \MASTERADDRINPROG_i_a2_0_a3_d_0[0]_net_1\);
    
    \arbRegSMCurrentState_ns_i_a2_1_o2_0_RNIJL905[0]\ : CFG4
      generic map(INIT => x"FF13")

      port map(A => N_89, B => \arbRegSMCurrentState_13\, C => 
        M0GATEDHTRANS, D => CoreAHBLite_0_AHBmslave3_HREADY_i_1, 
        Y => \MASTERADDRINPROG_i_a2_0_a3_1_0[0]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \arbRegSMCurrentState_RNO[15]\ : CFG4
      generic map(INIT => x"88A8")

      port map(A => CoreAHBLite_0_AHBmslave3_HREADY_i_1, B => 
        \arbRegSMCurrentState_13\, C => sAddrDec(3), D => 
        \arbRegSMCurrentState_ns_i_a2_1_o4_0[0]_net_1\, Y => 
        N_104_i_0);
    
    \arbRegSMCurrentState[14]\ : SLE
      port map(D => N_105, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_12\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \arbRegSMCurrentState_ns_i_a2_1_o2_0[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \arbRegSMCurrentState_12\, B => 
        \arbRegSMCurrentState_0\, Y => N_89);
    
    \arbRegSMCurrentState_ns_i_a2_1_o4_0[0]\ : CFG4
      generic map(INIT => x"5F77")

      port map(A => N_89, B => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        C => regHTRANS, D => masterRegAddrSel, Y => 
        \arbRegSMCurrentState_ns_i_a2_1_o4_0[0]_net_1\);
    
    \arbRegSMCurrentState_ns_i_a2_1_o4_0_RNIO5DT[0]\ : CFG4
      generic map(INIT => x"B0A0")

      port map(A => \arbRegSMCurrentState_13\, B => 
        \arbRegSMCurrentState_ns_i_a2_1_o4_0[0]_net_1\, C => 
        M0GATEDHWRITE, D => sAddrDec(3), Y => N_7_i_0);
    
    \arbRegSMCurrentState[2]\ : SLE
      port map(D => GND_net_1, CLK => FAB_CCC_GL0, EN => 
        xhdl1221_i_0(3), ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_0\);
    
    \arbRegSMCurrentState_ns_i_i_m3[1]\ : CFG4
      generic map(INIT => x"3075")

      port map(A => \MASTERADDRINPROG_i_a2_0_a3_1_0[0]\, B => 
        xhdl1221_i_0(3), C => \arbRegSMCurrentState_12\, D => 
        \MASTERADDRINPROG_i_a2_0_a3_d_0[0]_net_1\, Y => N_105);
    
    \MASTERADDRINPROG_i_a2_0_a3_d_d[0]\ : CFG3
      generic map(INIT => x"45")

      port map(A => \arbRegSMCurrentState_13\, B => 
        M0GATEDHADDR_2, C => M0GATEDHADDR_0, Y => 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0));
    
    \MASTERADDRINPROG_i_a2_0_a3_0_0[0]\ : CFG4
      generic map(INIT => x"1F3F")

      port map(A => N_89, B => \arbRegSMCurrentState_13\, C => 
        M0GATEDHTRANS, D => un3_saddrdec_i_a2_3_0, Y => 
        MASTERADDRINPROG_i_a2_0_a3_0(0));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVESTAGE_0 is

    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA : in    std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave3_HWDATA                          : out   std_logic_vector(31 downto 0);
          sAddrDec                                                 : in    std_logic_vector(3 to 3);
          xhdl1249                                                 : out   std_logic_vector(0 to 0);
          xhdl1221_i_0                                             : in    std_logic_vector(3 to 3);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS : in    std_logic_vector(1 to 1);
          MASTERADDRINPROG_i_a2_0_a3_d_d                           : out   std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_0                             : out   std_logic_vector(0 to 0);
          arbRegSMCurrentState_13                                  : out   std_logic;
          arbRegSMCurrentState_12                                  : out   std_logic;
          arbRegSMCurrentState_0                                   : out   std_logic;
          M0GATEDHADDR_2                                           : in    std_logic;
          M0GATEDHADDR_0                                           : in    std_logic;
          hwdata10                                                 : out   std_logic;
          MSS_READY                                                : in    std_logic;
          FAB_CCC_GL0                                              : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                  : in    std_logic;
          M0GATEDHTRANS                                            : in    std_logic;
          regHTRANS                                                : in    std_logic;
          masterRegAddrSel                                         : in    std_logic;
          un3_saddrdec_i_a2_3_0                                    : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                      : in    std_logic;
          M0GATEDHWRITE                                            : in    std_logic;
          N_7_i_0                                                  : out   std_logic;
          N_25_i_0                                                 : out   std_logic
        );

end COREAHBLITE_SLAVESTAGE_0;

architecture DEF_ARCH of COREAHBLITE_SLAVESTAGE_0 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVEARBITER_1
    port( xhdl1221_i_0                                             : in    std_logic_vector(3 to 3) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS : in    std_logic_vector(1 to 1) := (others => 'U');
          MASTERADDRINPROG_i_a2_0_a3_d_d                           : out   std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_0                             : out   std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_1_0                           : out   std_logic_vector(0 to 0);
          sAddrDec                                                 : in    std_logic_vector(3 to 3) := (others => 'U');
          arbRegSMCurrentState_13                                  : out   std_logic;
          arbRegSMCurrentState_12                                  : out   std_logic;
          arbRegSMCurrentState_0                                   : out   std_logic;
          M0GATEDHADDR_2                                           : in    std_logic := 'U';
          M0GATEDHADDR_0                                           : in    std_logic := 'U';
          MSS_READY                                                : in    std_logic := 'U';
          FAB_CCC_GL0                                              : in    std_logic := 'U';
          regHTRANS                                                : in    std_logic := 'U';
          masterRegAddrSel                                         : in    std_logic := 'U';
          un3_saddrdec_i_a2_3_0                                    : in    std_logic := 'U';
          M0GATEDHTRANS                                            : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                      : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HSELx_i_1_i_0                   : out   std_logic;
          M0GATEDHWRITE                                            : in    std_logic := 'U';
          N_7_i_0                                                  : out   std_logic;
          N_25_i_0                                                 : out   std_logic
        );
  end component;

    signal \hwdata10\, VCC_net_1, 
        CoreAHBLite_0_AHBmslave3_HSELx_i_1_i_0, GND_net_1, 
        \MASTERADDRINPROG_i_a2_0_a3_1_0[0]\ : std_logic;

    for all : COREAHBLITE_SLAVEARBITER_1
	Use entity work.COREAHBLITE_SLAVEARBITER_1(DEF_ARCH);
begin 

    hwdata10 <= \hwdata10\;

    \masterDataInProg_RNICEPO_6[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(1));
    
    \masterDataInProg_RNICEPO_8[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(9));
    
    \masterDataInProg_RNICEPO_23[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(23));
    
    \masterDataInProg_RNICEPO_17[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(29));
    
    \masterDataInProg_RNICEPO_15[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(31));
    
    \masterDataInProg_RNICEPO_12[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(12));
    
    \masterDataInProg_RNICEPO_20[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(26));
    
    \masterDataInProg_RNICEPO_24[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(22));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \masterDataInProg_RNICEPO_21[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(25));
    
    \MADDRREADY_5_iv[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => sAddrDec(3), B => M0GATEDHTRANS, C => 
        \MASTERADDRINPROG_i_a2_0_a3_1_0[0]\, Y => xhdl1249(0));
    
    \masterDataInProg_RNICEPO[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(8));
    
    \masterDataInProg_RNICEPO_1[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(6));
    
    \masterDataInProg_RNICEPO_7[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(0));
    
    \masterDataInProg_RNICEPO_18[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(28));
    
    \masterDataInProg_RNICEPO_26[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(20));
    
    \masterDataInProg_RNICEPO_13[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(11));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \masterDataInProg_RNICEPO_30[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(16));
    
    \masterDataInProg[0]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave3_HSELx_i_1_i_0, CLK
         => FAB_CCC_GL0, EN => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \hwdata10\);
    
    \masterDataInProg_RNICEPO_29[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(17));
    
    \masterDataInProg_RNICEPO_10[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(14));
    
    \masterDataInProg_RNICEPO_14[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(10));
    
    \masterDataInProg_RNICEPO_3[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(4));
    
    \masterDataInProg_RNICEPO_11[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(13));
    
    \masterDataInProg_RNICEPO_9[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(15));
    
    \masterDataInProg_RNICEPO_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(3));
    
    \masterDataInProg_RNICEPO_27[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(19));
    
    \masterDataInProg_RNICEPO_25[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(21));
    
    \masterDataInProg_RNICEPO_22[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(24));
    
    slave_arbiter : COREAHBLITE_SLAVEARBITER_1
      port map(xhdl1221_i_0(3) => xhdl1221_i_0(3), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0) => 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0), 
        MASTERADDRINPROG_i_a2_0_a3_0(0) => 
        MASTERADDRINPROG_i_a2_0_a3_0(0), 
        MASTERADDRINPROG_i_a2_0_a3_1_0(0) => 
        \MASTERADDRINPROG_i_a2_0_a3_1_0[0]\, sAddrDec(3) => 
        sAddrDec(3), arbRegSMCurrentState_13 => 
        arbRegSMCurrentState_13, arbRegSMCurrentState_12 => 
        arbRegSMCurrentState_12, arbRegSMCurrentState_0 => 
        arbRegSMCurrentState_0, M0GATEDHADDR_2 => M0GATEDHADDR_2, 
        M0GATEDHADDR_0 => M0GATEDHADDR_0, MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, regHTRANS => regHTRANS, 
        masterRegAddrSel => masterRegAddrSel, 
        un3_saddrdec_i_a2_3_0 => un3_saddrdec_i_a2_3_0, 
        M0GATEDHTRANS => M0GATEDHTRANS, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, 
        CoreAHBLite_0_AHBmslave3_HSELx_i_1_i_0 => 
        CoreAHBLite_0_AHBmslave3_HSELx_i_1_i_0, M0GATEDHWRITE => 
        M0GATEDHWRITE, N_7_i_0 => N_7_i_0, N_25_i_0 => N_25_i_0);
    
    \masterDataInProg_RNICEPO_0[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(7));
    
    \masterDataInProg_RNICEPO_2[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(5));
    
    \masterDataInProg_RNICEPO_16[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(30));
    
    \masterDataInProg_RNICEPO_19[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(27));
    
    \masterDataInProg_RNICEPO_5[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(2));
    
    \masterDataInProg_RNICEPO_28[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        B => \hwdata10\, Y => CoreAHBLite_0_AHBmslave3_HWDATA(18));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_DEFAULTSLAVESM_0 is

    port( xhdl1250_i_m_1                      : in    std_logic_vector(0 to 0);
          SDATASELInt_7                       : in    std_logic;
          SDATASELInt_5                       : in    std_logic;
          SDATASELInt_4                       : in    std_logic;
          SDATASELInt_0                       : in    std_logic;
          defSlaveSMCurrentState              : out   std_logic;
          MSS_READY                           : in    std_logic;
          FAB_CCC_GL0                         : in    std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3_0   : in    std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3_1   : in    std_logic;
          defSlaveSMNextState_m_0_a3_0_0      : out   std_logic;
          HREADY_M_iv_i_0                     : out   std_logic;
          N_42_2                              : out   std_logic;
          N_63                                : in    std_logic;
          N_65                                : in    std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_2     : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_m_0 : in    std_logic;
          defSlaveSMNextState_m_0_a3_d        : out   std_logic;
          defSlaveSMNextState_m               : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3     : in    std_logic;
          N_114                               : in    std_logic;
          N_4_i_0                             : out   std_logic
        );

end COREAHBLITE_DEFAULTSLAVESM_0;

architecture DEF_ARCH of COREAHBLITE_DEFAULTSLAVESM_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal defSlaveSMCurrentState_net_1, VCC_net_1, N_9_i_0, 
        GND_net_1, \defSlaveSMNextState_m_0_a3_0_0\, \N_42_2\
         : std_logic;

begin 

    defSlaveSMCurrentState <= defSlaveSMCurrentState_net_1;
    defSlaveSMNextState_m_0_a3_0_0 <= 
        \defSlaveSMNextState_m_0_a3_0_0\;
    N_42_2 <= \N_42_2\;

    defSlaveSMNextState_i_a3_1 : CFG4
      generic map(INIT => x"0001")

      port map(A => SDATASELInt_7, B => SDATASELInt_5, C => 
        SDATASELInt_4, D => SDATASELInt_0, Y => \N_42_2\);
    
    defSlaveSMCurrentState_RNI6KMQJ : CFG4
      generic map(INIT => x"3332")

      port map(A => un1_hready_m_xhdl342_1_i_0_o3_3_0, B => 
        defSlaveSMCurrentState_net_1, C => 
        un1_hready_m_xhdl342_1_i_0_o3_2, D => 
        un1_hready_m_xhdl342_1_i_0_o3_3_1, Y => 
        defSlaveSMNextState_m);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    defSlaveSMCurrentState_RNI2QMTO : CFG4
      generic map(INIT => x"00AB")

      port map(A => defSlaveSMCurrentState_net_1, B => 
        un1_hready_m_xhdl342_1_i_0_o3_3_0, C => 
        un1_hready_m_xhdl342_1_i_0_o3_3_1, D => 
        \defSlaveSMNextState_m_0_a3_0_0\, Y => HREADY_M_iv_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    defSlaveSMCurrentState_RNIK4LSB : CFG3
      generic map(INIT => x"54")

      port map(A => defSlaveSMCurrentState_net_1, B => 
        un1_hready_m_xhdl342_1_i_0_o3_3_0, C => 
        un1_hready_m_xhdl342_1_i_0_o3_3_1, Y => 
        defSlaveSMNextState_m_0_a3_d);
    
    defSlaveSMCurrentState_RNIEP4SN : CFG4
      generic map(INIT => x"00AB")

      port map(A => defSlaveSMCurrentState_net_1, B => 
        un1_hready_m_xhdl342_1_i_0_o3_2, C => 
        un1_hready_m_xhdl342_1_i_0_o3_3, D => N_114, Y => N_4_i_0);
    
    defSlaveSMCurrentState_RNO : CFG4
      generic map(INIT => x"070F")

      port map(A => \N_42_2\, B => N_63, C => 
        defSlaveSMCurrentState_net_1, D => N_65, Y => N_9_i_0);
    
    defSlaveSMCurrentState_RNIEL11D : CFG4
      generic map(INIT => x"44F4")

      port map(A => defSlaveSMCurrentState_net_1, B => 
        un1_hready_m_xhdl342_1_i_0_o3_2, C => xhdl1250_i_m_1(0), 
        D => CoreAHBLite_0_AHBmslave3_HREADY_m_0, Y => 
        \defSlaveSMNextState_m_0_a3_0_0\);
    
    \defSlaveSMCurrentState\ : SLE
      port map(D => N_9_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        defSlaveSMCurrentState_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MASTERSTAGE_1_1_0_8_0 is

    port( xhdl1221_i_0                                               : out   std_logic_vector(3 to 3);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0);
          xhdl1249                                                   : in    std_logic_vector(0 to 0);
          xhdl1250_i_m_1                                             : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1);
          M0GATEDHSIZE                                               : out   std_logic_vector(1 downto 0);
          sAddrDec                                                   : out   std_logic_vector(3 to 3);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          arbRegSMCurrentState_0                                     : in    std_logic;
          arbRegSMCurrentState_12                                    : in    std_logic;
          arbRegSMCurrentState_13                                    : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28 : in    std_logic;
          M0GATEDHADDR_31                                            : out   std_logic;
          M0GATEDHADDR_29                                            : out   std_logic;
          M0GATEDHADDR_0                                             : out   std_logic;
          M0GATEDHADDR_1                                             : out   std_logic;
          M0GATEDHADDR_2                                             : out   std_logic;
          M0GATEDHADDR_3                                             : out   std_logic;
          M0GATEDHADDR_12                                            : out   std_logic;
          M0GATEDHADDR_13                                            : out   std_logic;
          M0GATEDHADDR_14                                            : out   std_logic;
          M0GATEDHADDR_15                                            : out   std_logic;
          M0GATEDHADDR_4                                             : out   std_logic;
          M0GATEDHADDR_5                                             : out   std_logic;
          M0GATEDHADDR_6                                             : out   std_logic;
          M0GATEDHADDR_7                                             : out   std_logic;
          M0GATEDHADDR_8                                             : out   std_logic;
          M0GATEDHADDR_9                                             : out   std_logic;
          M0GATEDHADDR_10                                            : out   std_logic;
          M0GATEDHADDR_11                                            : out   std_logic;
          MSS_READY                                                  : in    std_logic;
          FAB_CCC_GL0                                                : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic;
          regHTRANS                                                  : out   std_logic;
          masterRegAddrSel                                           : out   std_logic;
          hwdata10                                                   : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                        : in    std_logic;
          M0GATEDHTRANS                                              : out   std_logic;
          M0GATEDHWRITE                                              : out   std_logic;
          un3_saddrdec_i_a2_3_0                                      : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_2                            : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3                            : out   std_logic;
          defSlaveSMCurrentState                                     : out   std_logic;
          HREADY_M_iv_i_0                                            : out   std_logic;
          defSlaveSMNextState_m                                      : out   std_logic
        );

end COREAHBLITE_MASTERSTAGE_1_1_0_8_0;

architecture DEF_ARCH of COREAHBLITE_MASTERSTAGE_1_1_0_8_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_DEFAULTSLAVESM_0
    port( xhdl1250_i_m_1                      : in    std_logic_vector(0 to 0) := (others => 'U');
          SDATASELInt_7                       : in    std_logic := 'U';
          SDATASELInt_5                       : in    std_logic := 'U';
          SDATASELInt_4                       : in    std_logic := 'U';
          SDATASELInt_0                       : in    std_logic := 'U';
          defSlaveSMCurrentState              : out   std_logic;
          MSS_READY                           : in    std_logic := 'U';
          FAB_CCC_GL0                         : in    std_logic := 'U';
          un1_hready_m_xhdl342_1_i_0_o3_3_0   : in    std_logic := 'U';
          un1_hready_m_xhdl342_1_i_0_o3_3_1   : in    std_logic := 'U';
          defSlaveSMNextState_m_0_a3_0_0      : out   std_logic;
          HREADY_M_iv_i_0                     : out   std_logic;
          N_42_2                              : out   std_logic;
          N_63                                : in    std_logic := 'U';
          N_65                                : in    std_logic := 'U';
          un1_hready_m_xhdl342_1_i_0_o3_2     : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_m_0 : in    std_logic := 'U';
          defSlaveSMNextState_m_0_a3_d        : out   std_logic;
          defSlaveSMNextState_m               : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3     : in    std_logic := 'U';
          N_114                               : in    std_logic := 'U';
          N_4_i_0                             : out   std_logic
        );
  end component;

    signal \SDATASELInt[1]_net_1\, VCC_net_1, 
        \SADDRSEL[1]_net_1\, N_4_i_0, GND_net_1, 
        \SDATASELInt[2]_net_1\, \SADDRSEL[2]_net_1\, 
        \xhdl1222[3]\, \xhdl1221_i_0[3]\, \SDATASELInt[4]_net_1\, 
        \SADDRSEL[4]_net_1\, \SDATASELInt[5]_net_1\, 
        \SADDRSEL[5]_net_1\, \SDATASELInt[6]_net_1\, 
        \SADDRSEL[6]_net_1\, \SDATASELInt[7]_net_1\, 
        \SADDRSEL[7]_net_1\, \SDATASELInt[8]_net_1\, 
        \SADDRSEL[8]_net_1\, \SDATASELInt[9]_net_1\, 
        \SADDRSEL[9]_net_1\, \SDATASELInt[10]_net_1\, 
        \SADDRSEL[10]_net_1\, \SDATASELInt[11]_net_1\, 
        \SADDRSEL[11]_net_1\, \SDATASELInt[12]_net_1\, 
        \SADDRSEL[12]_net_1\, \SDATASELInt[13]_net_1\, 
        \SADDRSEL[13]_net_1\, \SDATASELInt[14]_net_1\, 
        \SADDRSEL[14]_net_1\, \SDATASELInt[15]_net_1\, 
        \SADDRSEL[15]_net_1\, \regHADDR[12]_net_1\, 
        \masterAddrClockEnable\, \regHADDR[13]_net_1\, 
        \regHADDR[14]_net_1\, \regHADDR[15]_net_1\, 
        \regHSIZE[0]_net_1\, \regHSIZE[1]_net_1\, 
        \SDATASELInt[0]_net_1\, \SADDRSEL[0]_net_1\, 
        \regHADDR[0]_net_1\, \regHADDR[1]_net_1\, 
        \regHADDR[2]_net_1\, \regHADDR[3]_net_1\, 
        \regHADDR[4]_net_1\, \regHADDR[5]_net_1\, 
        \regHADDR[6]_net_1\, \regHADDR[7]_net_1\, 
        \regHADDR[8]_net_1\, \regHADDR[9]_net_1\, 
        \regHADDR[10]_net_1\, \regHADDR[11]_net_1\, \regHWRITE\, 
        regHTRANS_net_1, masterRegAddrSel_net_1, 
        d_masterRegAddrSel, \MASTERADDRINPROG_i_a2_0_a3_c_c[0]\, 
        N_63, un1_hready_m_xhdl342_1_i_0_o3_3_0_1, 
        un1_hready_m_xhdl342_1_i_0_o3_3_0, N_19, N_14, N_42_2, 
        N_65, \un88_htrans\, CoreAHBLite_0_AHBmslave3_HREADY_m_0, 
        \xhdl1250_i_m_1[0]\, \M0GATEDHADDR[28]\, 
        \M0GATEDHADDR_31\, \M0GATEDHTRANS\, \SADDRSEL_1[0]_net_1\, 
        \M0GATEDHADDR[30]\, \M0GATEDHADDR_29\, 
        un1_hready_m_xhdl342_1_i_0_a7_1_0, 
        un1_hready_m_xhdl342_1_i_0_a7_3_0, 
        un1_hready_m_xhdl342_1_i_0_a7_0_0, 
        un1_hready_m_xhdl342_1_i_0_a7_2_0, \SADDRSEL_2[12]\, N_58, 
        N_59, un3_saddrdec_i_a2_3_0_net_1, \SADDRSEL_1[6]\, 
        \SADDRSEL_2[8]\, \SADDRSEL_1[9]\, \sAddrDec[3]\, N_41_2, 
        N_39_2, un1_hready_m_xhdl342_1_i_0_o3_3_1, 
        \un1_hready_m_xhdl342_1_i_0_o3_2\, N_114, 
        \un88_htrans_2_1\, \un1_hready_m_xhdl342_1_i_0_o3_3\, 
        \un88_htrans_2\, defSlaveSMNextState_m_0_a3_0_0, 
        defSlaveSMNextState_m_0_a3_d : std_logic;

    for all : COREAHBLITE_DEFAULTSLAVESM_0
	Use entity work.COREAHBLITE_DEFAULTSLAVESM_0(DEF_ARCH);
begin 

    xhdl1221_i_0(3) <= \xhdl1221_i_0[3]\;
    xhdl1250_i_m_1(0) <= \xhdl1250_i_m_1[0]\;
    sAddrDec(3) <= \sAddrDec[3]\;
    M0GATEDHADDR_31 <= \M0GATEDHADDR_31\;
    M0GATEDHADDR_29 <= \M0GATEDHADDR_29\;
    regHTRANS <= regHTRANS_net_1;
    masterRegAddrSel <= masterRegAddrSel_net_1;
    M0GATEDHTRANS <= \M0GATEDHTRANS\;
    un3_saddrdec_i_a2_3_0 <= un3_saddrdec_i_a2_3_0_net_1;
    un1_hready_m_xhdl342_1_i_0_o3_2 <= 
        \un1_hready_m_xhdl342_1_i_0_o3_2\;
    un1_hready_m_xhdl342_1_i_0_o3_3 <= 
        \un1_hready_m_xhdl342_1_i_0_o3_3\;

    \SADDRSEL[12]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        B => \M0GATEDHADDR[30]\, C => \M0GATEDHADDR_29\, D => 
        \SADDRSEL_2[12]\, Y => \SADDRSEL[12]_net_1\);
    
    \PREGATEDHADDR[11]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[11]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11, 
        Y => M0GATEDHADDR_11);
    
    \PREGATEDHADDR[12]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[12]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12, 
        Y => M0GATEDHADDR_12);
    
    \GATEDHSIZE[0]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHSIZE[0]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0), 
        Y => M0GATEDHSIZE(0));
    
    \PREGATEDHADDR[31]\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        B => masterRegAddrSel_net_1, Y => \M0GATEDHADDR_31\);
    
    un3_saddrdec_i_a2_3 : CFG4
      generic map(INIT => x"0040")

      port map(A => \M0GATEDHADDR[30]\, B => \M0GATEDHADDR[28]\, 
        C => \M0GATEDHADDR_29\, D => \M0GATEDHADDR_31\, Y => 
        \sAddrDec[3]\);
    
    \regHADDR[15]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[15]_net_1\);
    
    \SDATASELInt_RNI3I3J1_1[8]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt[15]_net_1\, B => 
        \SDATASELInt[13]_net_1\, C => \SDATASELInt[10]_net_1\, D
         => \SDATASELInt[8]_net_1\, Y => N_58);
    
    \SADDRSEL[13]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        B => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        C => \M0GATEDHADDR_29\, D => \SADDRSEL_1[9]\, Y => 
        \SADDRSEL[13]_net_1\);
    
    hready_m_xhdl347_1_0_0_a2_1_0_a2_RNIM5TB2_0 : CFG4
      generic map(INIT => x"0800")

      port map(A => N_58, B => N_42_2, C => \xhdl1222[3]\, D => 
        N_65, Y => N_39_2);
    
    \regHADDR[7]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[7]_net_1\);
    
    \SADDRSEL_i_o3[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sAddrDec[3]\, B => \M0GATEDHTRANS\, Y => 
        \xhdl1221_i_0[3]\);
    
    \SADDRSEL[1]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \M0GATEDHADDR_29\, B => \SADDRSEL_1[9]\, C
         => \M0GATEDHADDR[30]\, D => \M0GATEDHADDR_31\, Y => 
        \SADDRSEL[1]_net_1\);
    
    \PREGATEDHADDR[10]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[10]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10, 
        Y => M0GATEDHADDR_10);
    
    \SADDRSEL[9]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        B => \M0GATEDHADDR[30]\, C => \M0GATEDHADDR_31\, D => 
        \SADDRSEL_1[9]\, Y => \SADDRSEL[9]_net_1\);
    
    \PREGATEDHADDR[30]\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        B => masterRegAddrSel_net_1, Y => \M0GATEDHADDR[30]\);
    
    \PREGATEDHADDR[0]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[0]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        Y => M0GATEDHADDR_0);
    
    hready_m_xhdl342_0_a2_1_a2_RNIST1N3 : CFG3
      generic map(INIT => x"02")

      port map(A => N_63, B => 
        un1_hready_m_xhdl342_1_i_0_o3_3_0_1, C => \xhdl1222[3]\, 
        Y => un1_hready_m_xhdl342_1_i_0_o3_3_0);
    
    hready_m_xhdl347_1_0_0_a2_1_0_a2_RNI9FS33 : CFG4
      generic map(INIT => x"153F")

      port map(A => N_19, B => N_14, C => N_42_2, D => N_65, Y
         => un1_hready_m_xhdl342_1_i_0_o3_3_0_1);
    
    \regHADDR[9]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[9]_net_1\);
    
    \SADDRSEL[11]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        B => \M0GATEDHADDR[30]\, C => \M0GATEDHADDR_31\, D => 
        \SADDRSEL_1[9]\, Y => \SADDRSEL[11]_net_1\);
    
    \masterRegAddrSel\ : SLE
      port map(D => d_masterRegAddrSel, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        masterRegAddrSel_net_1);
    
    \regHTRANS\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHTRANS_net_1);
    
    hready_m_xhdl342_0_a2_1_a2_RNIED3LB : CFG2
      generic map(INIT => x"E")

      port map(A => un1_hready_m_xhdl342_1_i_0_o3_3_1, B => 
        un1_hready_m_xhdl342_1_i_0_o3_3_0, Y => 
        \un1_hready_m_xhdl342_1_i_0_o3_3\);
    
    \SADDRSEL_1[11]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \M0GATEDHTRANS\, B => \M0GATEDHADDR[28]\, Y
         => \SADDRSEL_1[9]\);
    
    GATEDHTRANS : CFG3
      generic map(INIT => x"B8")

      port map(A => regHTRANS_net_1, B => masterRegAddrSel_net_1, 
        C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        Y => \M0GATEDHTRANS\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \PREGATEDHADDR[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[5]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        Y => M0GATEDHADDR_5);
    
    \SADDRSEL[15]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        B => \M0GATEDHADDR[30]\, C => \M0GATEDHADDR_31\, D => 
        \SADDRSEL_1[9]\, Y => \SADDRSEL[15]_net_1\);
    
    \SADDRSEL_2[4]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \M0GATEDHADDR_29\, B => \M0GATEDHADDR[28]\, Y
         => \SADDRSEL_2[8]\);
    
    \SADDRSEL[0]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \M0GATEDHADDR_29\, B => \SADDRSEL_1[0]_net_1\, 
        C => \M0GATEDHADDR[30]\, Y => \SADDRSEL[0]_net_1\);
    
    hready_m_xhdl342_0_a2_1_a3_RNI85E14 : CFG2
      generic map(INIT => x"8")

      port map(A => \xhdl1250_i_m_1[0]\, B => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, Y => N_114);
    
    \un3_saddrdec_i_a2_3_0\ : CFG4
      generic map(INIT => x"8B88")

      port map(A => regHTRANS_net_1, B => masterRegAddrSel_net_1, 
        C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        Y => un3_saddrdec_i_a2_3_0_net_1);
    
    \SDATASELInt_RNIGU1I1[0]\ : CFG4
      generic map(INIT => x"0116")

      port map(A => \SDATASELInt[7]_net_1\, B => 
        \SDATASELInt[5]_net_1\, C => \SDATASELInt[4]_net_1\, D
         => \SDATASELInt[0]_net_1\, Y => N_19);
    
    \regHADDR[10]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[10]_net_1\);
    
    \SDATASELInt_RNIPBH51[1]\ : CFG3
      generic map(INIT => x"16")

      port map(A => \SDATASELInt[6]_net_1\, B => 
        \SDATASELInt[2]_net_1\, C => \SDATASELInt[1]_net_1\, Y
         => N_14);
    
    \SDATASELInt_RNI3I3J1[9]\ : CFG4
      generic map(INIT => x"0104")

      port map(A => \SDATASELInt[14]_net_1\, B => 
        \SDATASELInt[12]_net_1\, C => \SDATASELInt[11]_net_1\, D
         => \SDATASELInt[9]_net_1\, Y => 
        un1_hready_m_xhdl342_1_i_0_a7_0_0);
    
    \regHADDR[13]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[13]_net_1\);
    
    \PREGATEDHADDR[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[6]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        Y => M0GATEDHADDR_6);
    
    \regHADDR[12]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[12]_net_1\);
    
    \PREGATEDHADDR[15]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[15]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15, 
        Y => M0GATEDHADDR_15);
    
    hready_m_xhdl342_0_a2_1_a2_RNI0T4JJ : CFG3
      generic map(INIT => x"FE")

      port map(A => un1_hready_m_xhdl342_1_i_0_o3_3_1, B => 
        \un1_hready_m_xhdl342_1_i_0_o3_2\, C => 
        un1_hready_m_xhdl342_1_i_0_o3_3_0, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0));
    
    \regHADDR[5]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[5]_net_1\);
    
    \GATEDHSIZE[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHSIZE[1]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1), 
        Y => M0GATEDHSIZE(1));
    
    \SDATASELInt[4]\ : SLE
      port map(D => \SADDRSEL[4]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[4]_net_1\);
    
    \SADDRSEL[8]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        B => \M0GATEDHADDR[30]\, C => \M0GATEDHADDR_31\, D => 
        \SADDRSEL_2[8]\, Y => \SADDRSEL[8]_net_1\);
    
    \regHADDR[2]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[2]_net_1\);
    
    hready_m_xhdl347_1_0_0_a2_1_0_a2 : CFG3
      generic map(INIT => x"01")

      port map(A => \SDATASELInt[6]_net_1\, B => 
        \SDATASELInt[2]_net_1\, C => \SDATASELInt[1]_net_1\, Y
         => N_65);
    
    \SDATASELInt[15]\ : SLE
      port map(D => \SADDRSEL[15]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[15]_net_1\);
    
    \PREGATEDHADDR[13]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[13]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13, 
        Y => M0GATEDHADDR_13);
    
    \SADDRSEL[10]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \SADDRSEL_1[6]\, B => \M0GATEDHADDR[30]\, C
         => \SADDRSEL_2[12]\, Y => \SADDRSEL[10]_net_1\);
    
    \PREGATEDHADDR[28]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => regHTRANS_net_1, B => masterRegAddrSel_net_1, 
        C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        Y => \M0GATEDHADDR[28]\);
    
    \SDATASELInt[14]\ : SLE
      port map(D => \SADDRSEL[14]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[14]_net_1\);
    
    \SDATASELInt[2]\ : SLE
      port map(D => \SADDRSEL[2]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[2]_net_1\);
    
    \regHADDR[8]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[8]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SDATASELInt_RNIIF1U7_0[8]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_hready_m_xhdl342_1_i_0_a7_3_0, B => 
        un1_hready_m_xhdl342_1_i_0_a7_1_0, C => N_39_2, D => 
        N_41_2, Y => un1_hready_m_xhdl342_1_i_0_o3_3_1);
    
    \PREGATEDHADDR[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[7]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7, 
        Y => M0GATEDHADDR_7);
    
    un88_htrans_2 : CFG4
      generic map(INIT => x"0080")

      port map(A => \M0GATEDHADDR_29\, B => \un88_htrans_2_1\, C
         => un3_saddrdec_i_a2_3_0_net_1, D => \M0GATEDHADDR_31\, 
        Y => \un88_htrans_2\);
    
    \SDATASELInt_RNIIF1U7[8]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => un1_hready_m_xhdl342_1_i_0_a7_2_0, B => 
        un1_hready_m_xhdl342_1_i_0_a7_0_0, C => N_41_2, D => 
        N_39_2, Y => \un1_hready_m_xhdl342_1_i_0_o3_2\);
    
    \SADDRSEL[7]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        B => \M0GATEDHADDR[30]\, C => \M0GATEDHADDR_31\, D => 
        \SADDRSEL_1[9]\, Y => \SADDRSEL[7]_net_1\);
    
    masterAddrClockEnable : CFG4
      generic map(INIT => x"0004")

      port map(A => defSlaveSMNextState_m_0_a3_0_0, B => 
        \un88_htrans_2\, C => masterRegAddrSel_net_1, D => 
        defSlaveSMNextState_m_0_a3_d, Y => 
        \masterAddrClockEnable\);
    
    d_masterRegAddrSel_ns : CFG3
      generic map(INIT => x"E2")

      port map(A => \un88_htrans\, B => masterRegAddrSel_net_1, C
         => xhdl1249(0), Y => d_masterRegAddrSel);
    
    \SDATASELInt_RNILEPK4[3]\ : CFG3
      generic map(INIT => x"20")

      port map(A => hwdata10, B => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, C => \xhdl1222[3]\, 
        Y => CoreAHBLite_0_AHBmslave3_HREADY_m_0);
    
    \SDATASELInt_RNI3I3J1_0[8]\ : CFG4
      generic map(INIT => x"0006")

      port map(A => \SDATASELInt[15]_net_1\, B => 
        \SDATASELInt[13]_net_1\, C => \SDATASELInt[10]_net_1\, D
         => \SDATASELInt[8]_net_1\, Y => 
        un1_hready_m_xhdl342_1_i_0_a7_2_0);
    
    \regHADDR[6]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[6]_net_1\);
    
    \PREGATEDHADDR[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[4]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        Y => M0GATEDHADDR_4);
    
    GATEDHWRITE : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHWRITE\, B => masterRegAddrSel_net_1, C
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        Y => M0GATEDHWRITE);
    
    \SDATASELInt[13]\ : SLE
      port map(D => \SADDRSEL[13]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[13]_net_1\);
    
    regHWRITE : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHWRITE\);
    
    \regHSIZE[1]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1), 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHSIZE[1]_net_1\);
    
    un88_htrans_2_1_RNO : CFG3
      generic map(INIT => x"01")

      port map(A => arbRegSMCurrentState_0, B => 
        arbRegSMCurrentState_12, C => arbRegSMCurrentState_13, Y
         => \MASTERADDRINPROG_i_a2_0_a3_c_c[0]\);
    
    \SADDRSEL[4]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        B => \M0GATEDHADDR[30]\, C => \M0GATEDHADDR_31\, D => 
        \SADDRSEL_2[8]\, Y => \SADDRSEL[4]_net_1\);
    
    \SDATASELInt[9]\ : SLE
      port map(D => \SADDRSEL[9]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[9]_net_1\);
    
    \SDATASELInt[1]\ : SLE
      port map(D => \SADDRSEL[1]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[1]_net_1\);
    
    \SDATASELInt[12]\ : SLE
      port map(D => \SADDRSEL[12]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[12]_net_1\);
    
    \SDATASELInt[0]\ : SLE
      port map(D => \SADDRSEL[0]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[0]_net_1\);
    
    \regHADDR[11]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[11]_net_1\);
    
    \regHADDR[0]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[0]_net_1\);
    
    hready_m_xhdl342_0_a2_1_a3 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_42_2, B => N_63, C => \xhdl1222[3]\, D => 
        N_65, Y => \xhdl1250_i_m_1[0]\);
    
    \SADDRSEL[5]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        B => \M0GATEDHADDR[30]\, C => \M0GATEDHADDR_31\, D => 
        \SADDRSEL_1[9]\, Y => \SADDRSEL[5]_net_1\);
    
    \SDATASELInt[5]\ : SLE
      port map(D => \SADDRSEL[5]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[5]_net_1\);
    
    \PREGATEDHADDR[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[1]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        Y => M0GATEDHADDR_1);
    
    \SADDRSEL[6]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        B => \M0GATEDHADDR[30]\, C => \M0GATEDHADDR_31\, D => 
        \SADDRSEL_1[6]\, Y => \SADDRSEL[6]_net_1\);
    
    \regHADDR[3]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[3]_net_1\);
    
    \SDATASELInt_RNI3I3J1_1[9]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt[14]_net_1\, B => 
        \SDATASELInt[12]_net_1\, C => \SDATASELInt[11]_net_1\, D
         => \SDATASELInt[9]_net_1\, Y => N_59);
    
    \SADDRSEL[14]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        B => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        C => \M0GATEDHADDR[28]\, D => \SADDRSEL_1[6]\, Y => 
        \SADDRSEL[14]_net_1\);
    
    un88_htrans : CFG4
      generic map(INIT => x"1000")

      port map(A => defSlaveSMNextState_m_0_a3_d, B => 
        defSlaveSMNextState_m_0_a3_0_0, C => \un88_htrans_2_1\, D
         => \sAddrDec[3]\, Y => \un88_htrans\);
    
    \SDATASELInt[3]\ : SLE
      port map(D => \xhdl1221_i_0[3]\, CLK => FAB_CCC_GL0, EN => 
        N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \xhdl1222[3]\);
    
    un88_htrans_2_1 : CFG4
      generic map(INIT => x"E000")

      port map(A => \MASTERADDRINPROG_i_a2_0_a3_c_c[0]\, B => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        D => \M0GATEDHTRANS\, Y => \un88_htrans_2_1\);
    
    \regHADDR[1]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[1]_net_1\);
    
    \SDATASELInt[7]\ : SLE
      port map(D => \SADDRSEL[7]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[7]_net_1\);
    
    \SADDRSEL_1[0]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \M0GATEDHADDR[28]\, B => \M0GATEDHADDR_31\, C
         => \M0GATEDHTRANS\, Y => \SADDRSEL_1[0]_net_1\);
    
    \regHSIZE[0]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0), 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHSIZE[0]_net_1\);
    
    hready_m_xhdl347_1_0_0_a2_1_0_a2_RNIM5TB2 : CFG4
      generic map(INIT => x"0800")

      port map(A => N_59, B => N_42_2, C => \xhdl1222[3]\, D => 
        N_65, Y => N_41_2);
    
    \PREGATEDHADDR[9]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[9]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9, 
        Y => M0GATEDHADDR_9);
    
    \PREGATEDHADDR[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[2]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        Y => M0GATEDHADDR_2);
    
    \SADDRSEL_1[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \M0GATEDHTRANS\, B => \M0GATEDHADDR_29\, Y
         => \SADDRSEL_1[6]\);
    
    hready_m_xhdl342_0_a2_1_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => N_58, B => N_59, Y => N_63);
    
    \SDATASELInt[6]\ : SLE
      port map(D => \SADDRSEL[6]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[6]_net_1\);
    
    \SADDRSEL_2[10]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \M0GATEDHADDR_31\, B => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        Y => \SADDRSEL_2[12]\);
    
    \PREGATEDHADDR[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[3]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        Y => M0GATEDHADDR_3);
    
    \PREGATEDHADDR[29]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => regHTRANS_net_1, B => masterRegAddrSel_net_1, 
        C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        Y => \M0GATEDHADDR_29\);
    
    \PREGATEDHADDR[8]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[8]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        Y => M0GATEDHADDR_8);
    
    \regHADDR[14]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[14]_net_1\);
    
    \SADDRSEL[2]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \M0GATEDHADDR[28]\, B => \M0GATEDHADDR[30]\, 
        C => \M0GATEDHADDR_31\, D => \SADDRSEL_1[6]\, Y => 
        \SADDRSEL[2]_net_1\);
    
    \SDATASELInt_RNI3I3J1_0[9]\ : CFG4
      generic map(INIT => x"0012")

      port map(A => \SDATASELInt[14]_net_1\, B => 
        \SDATASELInt[12]_net_1\, C => \SDATASELInt[11]_net_1\, D
         => \SDATASELInt[9]_net_1\, Y => 
        un1_hready_m_xhdl342_1_i_0_a7_1_0);
    
    \SDATASELInt_RNI3I3J1[8]\ : CFG4
      generic map(INIT => x"0110")

      port map(A => \SDATASELInt[15]_net_1\, B => 
        \SDATASELInt[13]_net_1\, C => \SDATASELInt[10]_net_1\, D
         => \SDATASELInt[8]_net_1\, Y => 
        un1_hready_m_xhdl342_1_i_0_a7_3_0);
    
    \PREGATEDHADDR[14]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[14]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14, 
        Y => M0GATEDHADDR_14);
    
    \SDATASELInt[11]\ : SLE
      port map(D => \SADDRSEL[11]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[11]_net_1\);
    
    \SDATASELInt[8]\ : SLE
      port map(D => \SADDRSEL[8]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[8]_net_1\);
    
    \regHADDR[4]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        CLK => FAB_CCC_GL0, EN => \masterAddrClockEnable\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHADDR[4]_net_1\);
    
    \SDATASELInt[10]\ : SLE
      port map(D => \SADDRSEL[10]_net_1\, CLK => FAB_CCC_GL0, EN
         => N_4_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDATASELInt[10]_net_1\);
    
    default_slave_sm : COREAHBLITE_DEFAULTSLAVESM_0
      port map(xhdl1250_i_m_1(0) => \xhdl1250_i_m_1[0]\, 
        SDATASELInt_7 => \SDATASELInt[7]_net_1\, SDATASELInt_5
         => \SDATASELInt[5]_net_1\, SDATASELInt_4 => 
        \SDATASELInt[4]_net_1\, SDATASELInt_0 => 
        \SDATASELInt[0]_net_1\, defSlaveSMCurrentState => 
        defSlaveSMCurrentState, MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, 
        un1_hready_m_xhdl342_1_i_0_o3_3_0 => 
        un1_hready_m_xhdl342_1_i_0_o3_3_0, 
        un1_hready_m_xhdl342_1_i_0_o3_3_1 => 
        un1_hready_m_xhdl342_1_i_0_o3_3_1, 
        defSlaveSMNextState_m_0_a3_0_0 => 
        defSlaveSMNextState_m_0_a3_0_0, HREADY_M_iv_i_0 => 
        HREADY_M_iv_i_0, N_42_2 => N_42_2, N_63 => N_63, N_65 => 
        N_65, un1_hready_m_xhdl342_1_i_0_o3_2 => 
        \un1_hready_m_xhdl342_1_i_0_o3_2\, 
        CoreAHBLite_0_AHBmslave3_HREADY_m_0 => 
        CoreAHBLite_0_AHBmslave3_HREADY_m_0, 
        defSlaveSMNextState_m_0_a3_d => 
        defSlaveSMNextState_m_0_a3_d, defSlaveSMNextState_m => 
        defSlaveSMNextState_m, un1_hready_m_xhdl342_1_i_0_o3_3
         => \un1_hready_m_xhdl342_1_i_0_o3_3\, N_114 => N_114, 
        N_4_i_0 => N_4_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MATRIX4X16 is

    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0);
          xhdl1250_i_m_1                                             : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1);
          M0GATEDHSIZE                                               : out   std_logic_vector(1 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave3_HWDATA                            : out   std_logic_vector(31 downto 0);
          MASTERADDRINPROG_i_a2_0_a3_d_d                             : out   std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_0                               : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28 : in    std_logic;
          M0GATEDHADDR_0                                             : out   std_logic;
          M0GATEDHADDR_1                                             : out   std_logic;
          M0GATEDHADDR_2                                             : out   std_logic;
          M0GATEDHADDR_3                                             : out   std_logic;
          M0GATEDHADDR_12                                            : out   std_logic;
          M0GATEDHADDR_13                                            : out   std_logic;
          M0GATEDHADDR_14                                            : out   std_logic;
          M0GATEDHADDR_15                                            : out   std_logic;
          M0GATEDHADDR_4                                             : out   std_logic;
          M0GATEDHADDR_5                                             : out   std_logic;
          M0GATEDHADDR_6                                             : out   std_logic;
          M0GATEDHADDR_7                                             : out   std_logic;
          M0GATEDHADDR_8                                             : out   std_logic;
          M0GATEDHADDR_9                                             : out   std_logic;
          M0GATEDHADDR_10                                            : out   std_logic;
          M0GATEDHADDR_11                                            : out   std_logic;
          MSS_READY                                                  : in    std_logic;
          FAB_CCC_GL0                                                : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                        : in    std_logic;
          M0GATEDHWRITE                                              : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_2                            : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3                            : out   std_logic;
          defSlaveSMCurrentState                                     : out   std_logic;
          HREADY_M_iv_i_0                                            : out   std_logic;
          defSlaveSMNextState_m                                      : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                    : in    std_logic;
          N_7_i_0                                                    : out   std_logic;
          N_25_i_0                                                   : out   std_logic
        );

end COREAHBLITE_MATRIX4X16;

architecture DEF_ARCH of COREAHBLITE_MATRIX4X16 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVESTAGE_0
    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HWDATA                          : out   std_logic_vector(31 downto 0);
          sAddrDec                                                 : in    std_logic_vector(3 to 3) := (others => 'U');
          xhdl1249                                                 : out   std_logic_vector(0 to 0);
          xhdl1221_i_0                                             : in    std_logic_vector(3 to 3) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS : in    std_logic_vector(1 to 1) := (others => 'U');
          MASTERADDRINPROG_i_a2_0_a3_d_d                           : out   std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_0                             : out   std_logic_vector(0 to 0);
          arbRegSMCurrentState_13                                  : out   std_logic;
          arbRegSMCurrentState_12                                  : out   std_logic;
          arbRegSMCurrentState_0                                   : out   std_logic;
          M0GATEDHADDR_2                                           : in    std_logic := 'U';
          M0GATEDHADDR_0                                           : in    std_logic := 'U';
          hwdata10                                                 : out   std_logic;
          MSS_READY                                                : in    std_logic := 'U';
          FAB_CCC_GL0                                              : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                  : in    std_logic := 'U';
          M0GATEDHTRANS                                            : in    std_logic := 'U';
          regHTRANS                                                : in    std_logic := 'U';
          masterRegAddrSel                                         : in    std_logic := 'U';
          un3_saddrdec_i_a2_3_0                                    : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                      : in    std_logic := 'U';
          M0GATEDHWRITE                                            : in    std_logic := 'U';
          N_7_i_0                                                  : out   std_logic;
          N_25_i_0                                                 : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MASTERSTAGE_1_1_0_8_0
    port( xhdl1221_i_0                                               : out   std_logic_vector(3 to 3);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0) := (others => 'U');
          xhdl1249                                                   : in    std_logic_vector(0 to 0) := (others => 'U');
          xhdl1250_i_m_1                                             : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1) := (others => 'U');
          M0GATEDHSIZE                                               : out   std_logic_vector(1 downto 0);
          sAddrDec                                                   : out   std_logic_vector(3 to 3);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          arbRegSMCurrentState_0                                     : in    std_logic := 'U';
          arbRegSMCurrentState_12                                    : in    std_logic := 'U';
          arbRegSMCurrentState_13                                    : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28 : in    std_logic := 'U';
          M0GATEDHADDR_31                                            : out   std_logic;
          M0GATEDHADDR_29                                            : out   std_logic;
          M0GATEDHADDR_0                                             : out   std_logic;
          M0GATEDHADDR_1                                             : out   std_logic;
          M0GATEDHADDR_2                                             : out   std_logic;
          M0GATEDHADDR_3                                             : out   std_logic;
          M0GATEDHADDR_12                                            : out   std_logic;
          M0GATEDHADDR_13                                            : out   std_logic;
          M0GATEDHADDR_14                                            : out   std_logic;
          M0GATEDHADDR_15                                            : out   std_logic;
          M0GATEDHADDR_4                                             : out   std_logic;
          M0GATEDHADDR_5                                             : out   std_logic;
          M0GATEDHADDR_6                                             : out   std_logic;
          M0GATEDHADDR_7                                             : out   std_logic;
          M0GATEDHADDR_8                                             : out   std_logic;
          M0GATEDHADDR_9                                             : out   std_logic;
          M0GATEDHADDR_10                                            : out   std_logic;
          M0GATEDHADDR_11                                            : out   std_logic;
          MSS_READY                                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                                : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          regHTRANS                                                  : out   std_logic;
          masterRegAddrSel                                           : out   std_logic;
          hwdata10                                                   : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                        : in    std_logic := 'U';
          M0GATEDHTRANS                                              : out   std_logic;
          M0GATEDHWRITE                                              : out   std_logic;
          un3_saddrdec_i_a2_3_0                                      : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_2                            : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3                            : out   std_logic;
          defSlaveSMCurrentState                                     : out   std_logic;
          HREADY_M_iv_i_0                                            : out   std_logic;
          defSlaveSMNextState_m                                      : out   std_logic
        );
  end component;

    signal \xhdl1221_i_0[3]\, \arbRegSMCurrentState[2]\, 
        \arbRegSMCurrentState[14]\, \arbRegSMCurrentState[15]\, 
        \xhdl1249[0]\, \M0GATEDHADDR[31]\, \M0GATEDHADDR[29]\, 
        \sAddrDec[3]\, regHTRANS, masterRegAddrSel, hwdata10, 
        M0GATEDHTRANS, \M0GATEDHWRITE\, un3_saddrdec_i_a2_3_0, 
        GND_net_1, VCC_net_1 : std_logic;

    for all : COREAHBLITE_SLAVESTAGE_0
	Use entity work.COREAHBLITE_SLAVESTAGE_0(DEF_ARCH);
    for all : COREAHBLITE_MASTERSTAGE_1_1_0_8_0
	Use entity work.COREAHBLITE_MASTERSTAGE_1_1_0_8_0(DEF_ARCH);
begin 

    M0GATEDHWRITE <= \M0GATEDHWRITE\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    slavestage_3 : COREAHBLITE_SLAVESTAGE_0
      port map(
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        CoreAHBLite_0_AHBmslave3_HWDATA(31) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), 
        CoreAHBLite_0_AHBmslave3_HWDATA(30) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), 
        CoreAHBLite_0_AHBmslave3_HWDATA(29) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), 
        CoreAHBLite_0_AHBmslave3_HWDATA(28) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), 
        CoreAHBLite_0_AHBmslave3_HWDATA(27) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), 
        CoreAHBLite_0_AHBmslave3_HWDATA(26) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), 
        CoreAHBLite_0_AHBmslave3_HWDATA(25) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), 
        CoreAHBLite_0_AHBmslave3_HWDATA(24) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), 
        CoreAHBLite_0_AHBmslave3_HWDATA(23) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), 
        CoreAHBLite_0_AHBmslave3_HWDATA(22) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), 
        CoreAHBLite_0_AHBmslave3_HWDATA(21) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), 
        CoreAHBLite_0_AHBmslave3_HWDATA(20) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), 
        CoreAHBLite_0_AHBmslave3_HWDATA(19) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), 
        CoreAHBLite_0_AHBmslave3_HWDATA(18) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), 
        CoreAHBLite_0_AHBmslave3_HWDATA(17) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), 
        CoreAHBLite_0_AHBmslave3_HWDATA(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), 
        CoreAHBLite_0_AHBmslave3_HWDATA(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), 
        CoreAHBLite_0_AHBmslave3_HWDATA(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), 
        CoreAHBLite_0_AHBmslave3_HWDATA(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), 
        CoreAHBLite_0_AHBmslave3_HWDATA(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), 
        CoreAHBLite_0_AHBmslave3_HWDATA(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), 
        CoreAHBLite_0_AHBmslave3_HWDATA(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), 
        CoreAHBLite_0_AHBmslave3_HWDATA(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), 
        CoreAHBLite_0_AHBmslave3_HWDATA(8) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), 
        CoreAHBLite_0_AHBmslave3_HWDATA(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(7), 
        CoreAHBLite_0_AHBmslave3_HWDATA(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(6), 
        CoreAHBLite_0_AHBmslave3_HWDATA(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), 
        CoreAHBLite_0_AHBmslave3_HWDATA(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), 
        CoreAHBLite_0_AHBmslave3_HWDATA(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), 
        CoreAHBLite_0_AHBmslave3_HWDATA(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), 
        CoreAHBLite_0_AHBmslave3_HWDATA(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), 
        CoreAHBLite_0_AHBmslave3_HWDATA(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), sAddrDec(3) => 
        \sAddrDec[3]\, xhdl1249(0) => \xhdl1249[0]\, 
        xhdl1221_i_0(3) => \xhdl1221_i_0[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0) => 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0), 
        MASTERADDRINPROG_i_a2_0_a3_0(0) => 
        MASTERADDRINPROG_i_a2_0_a3_0(0), arbRegSMCurrentState_13
         => \arbRegSMCurrentState[15]\, arbRegSMCurrentState_12
         => \arbRegSMCurrentState[14]\, arbRegSMCurrentState_0
         => \arbRegSMCurrentState[2]\, M0GATEDHADDR_2 => 
        \M0GATEDHADDR[31]\, M0GATEDHADDR_0 => \M0GATEDHADDR[29]\, 
        hwdata10 => hwdata10, MSS_READY => MSS_READY, FAB_CCC_GL0
         => FAB_CCC_GL0, CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0
         => CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, 
        M0GATEDHTRANS => M0GATEDHTRANS, regHTRANS => regHTRANS, 
        masterRegAddrSel => masterRegAddrSel, 
        un3_saddrdec_i_a2_3_0 => un3_saddrdec_i_a2_3_0, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, M0GATEDHWRITE => 
        \M0GATEDHWRITE\, N_7_i_0 => N_7_i_0, N_25_i_0 => N_25_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    masterstage_0 : COREAHBLITE_MASTERSTAGE_1_1_0_8_0
      port map(xhdl1221_i_0(3) => \xhdl1221_i_0[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0), 
        xhdl1249(0) => \xhdl1249[0]\, xhdl1250_i_m_1(0) => 
        xhdl1250_i_m_1(0), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        M0GATEDHSIZE(1) => M0GATEDHSIZE(1), M0GATEDHSIZE(0) => 
        M0GATEDHSIZE(0), sAddrDec(3) => \sAddrDec[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        arbRegSMCurrentState_0 => \arbRegSMCurrentState[2]\, 
        arbRegSMCurrentState_12 => \arbRegSMCurrentState[14]\, 
        arbRegSMCurrentState_13 => \arbRegSMCurrentState[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        M0GATEDHADDR_31 => \M0GATEDHADDR[31]\, M0GATEDHADDR_29
         => \M0GATEDHADDR[29]\, M0GATEDHADDR_0 => M0GATEDHADDR_0, 
        M0GATEDHADDR_1 => M0GATEDHADDR_1, M0GATEDHADDR_2 => 
        M0GATEDHADDR_2, M0GATEDHADDR_3 => M0GATEDHADDR_3, 
        M0GATEDHADDR_12 => M0GATEDHADDR_12, M0GATEDHADDR_13 => 
        M0GATEDHADDR_13, M0GATEDHADDR_14 => M0GATEDHADDR_14, 
        M0GATEDHADDR_15 => M0GATEDHADDR_15, M0GATEDHADDR_4 => 
        M0GATEDHADDR_4, M0GATEDHADDR_5 => M0GATEDHADDR_5, 
        M0GATEDHADDR_6 => M0GATEDHADDR_6, M0GATEDHADDR_7 => 
        M0GATEDHADDR_7, M0GATEDHADDR_8 => M0GATEDHADDR_8, 
        M0GATEDHADDR_9 => M0GATEDHADDR_9, M0GATEDHADDR_10 => 
        M0GATEDHADDR_10, M0GATEDHADDR_11 => M0GATEDHADDR_11, 
        MSS_READY => MSS_READY, FAB_CCC_GL0 => FAB_CCC_GL0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        regHTRANS => regHTRANS, masterRegAddrSel => 
        masterRegAddrSel, hwdata10 => hwdata10, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, M0GATEDHTRANS => 
        M0GATEDHTRANS, M0GATEDHWRITE => \M0GATEDHWRITE\, 
        un3_saddrdec_i_a2_3_0 => un3_saddrdec_i_a2_3_0, 
        un1_hready_m_xhdl342_1_i_0_o3_2 => 
        un1_hready_m_xhdl342_1_i_0_o3_2, 
        un1_hready_m_xhdl342_1_i_0_o3_3 => 
        un1_hready_m_xhdl342_1_i_0_o3_3, defSlaveSMCurrentState
         => defSlaveSMCurrentState, HREADY_M_iv_i_0 => 
        HREADY_M_iv_i_0, defSlaveSMNextState_m => 
        defSlaveSMNextState_m);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLite is

    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0);
          xhdl1250_i_m_1                                             : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1);
          M0GATEDHSIZE                                               : out   std_logic_vector(1 downto 0);
          M0GATEDHADDR                                               : out   std_logic_vector(15 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave3_HWDATA                            : out   std_logic_vector(31 downto 0);
          MASTERADDRINPROG_i_a2_0_a3_d_d                             : out   std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_0                               : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28 : in    std_logic;
          MSS_READY                                                  : in    std_logic;
          FAB_CCC_GL0                                                : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                        : in    std_logic;
          M0GATEDHWRITE                                              : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_2                            : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3                            : out   std_logic;
          defSlaveSMCurrentState                                     : out   std_logic;
          HREADY_M_iv_i_0                                            : out   std_logic;
          defSlaveSMNextState_m                                      : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                    : in    std_logic;
          N_7_i_0                                                    : out   std_logic;
          N_25_i_0                                                   : out   std_logic
        );

end CoreAHBLite;

architecture DEF_ARCH of CoreAHBLite is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MATRIX4X16
    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0) := (others => 'U');
          xhdl1250_i_m_1                                             : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1) := (others => 'U');
          M0GATEDHSIZE                                               : out   std_logic_vector(1 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HWDATA                            : out   std_logic_vector(31 downto 0);
          MASTERADDRINPROG_i_a2_0_a3_d_d                             : out   std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_0                               : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28 : in    std_logic := 'U';
          M0GATEDHADDR_0                                             : out   std_logic;
          M0GATEDHADDR_1                                             : out   std_logic;
          M0GATEDHADDR_2                                             : out   std_logic;
          M0GATEDHADDR_3                                             : out   std_logic;
          M0GATEDHADDR_12                                            : out   std_logic;
          M0GATEDHADDR_13                                            : out   std_logic;
          M0GATEDHADDR_14                                            : out   std_logic;
          M0GATEDHADDR_15                                            : out   std_logic;
          M0GATEDHADDR_4                                             : out   std_logic;
          M0GATEDHADDR_5                                             : out   std_logic;
          M0GATEDHADDR_6                                             : out   std_logic;
          M0GATEDHADDR_7                                             : out   std_logic;
          M0GATEDHADDR_8                                             : out   std_logic;
          M0GATEDHADDR_9                                             : out   std_logic;
          M0GATEDHADDR_10                                            : out   std_logic;
          M0GATEDHADDR_11                                            : out   std_logic;
          MSS_READY                                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                                : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                        : in    std_logic := 'U';
          M0GATEDHWRITE                                              : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_2                            : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3                            : out   std_logic;
          defSlaveSMCurrentState                                     : out   std_logic;
          HREADY_M_iv_i_0                                            : out   std_logic;
          defSlaveSMNextState_m                                      : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                    : in    std_logic := 'U';
          N_7_i_0                                                    : out   std_logic;
          N_25_i_0                                                   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : COREAHBLITE_MATRIX4X16
	Use entity work.COREAHBLITE_MATRIX4X16(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    matrix4x16 : COREAHBLITE_MATRIX4X16
      port map(
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0), 
        xhdl1250_i_m_1(0) => xhdl1250_i_m_1(0), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        M0GATEDHSIZE(1) => M0GATEDHSIZE(1), M0GATEDHSIZE(0) => 
        M0GATEDHSIZE(0), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        CoreAHBLite_0_AHBmslave3_HWDATA(31) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), 
        CoreAHBLite_0_AHBmslave3_HWDATA(30) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), 
        CoreAHBLite_0_AHBmslave3_HWDATA(29) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), 
        CoreAHBLite_0_AHBmslave3_HWDATA(28) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), 
        CoreAHBLite_0_AHBmslave3_HWDATA(27) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), 
        CoreAHBLite_0_AHBmslave3_HWDATA(26) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), 
        CoreAHBLite_0_AHBmslave3_HWDATA(25) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), 
        CoreAHBLite_0_AHBmslave3_HWDATA(24) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), 
        CoreAHBLite_0_AHBmslave3_HWDATA(23) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), 
        CoreAHBLite_0_AHBmslave3_HWDATA(22) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), 
        CoreAHBLite_0_AHBmslave3_HWDATA(21) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), 
        CoreAHBLite_0_AHBmslave3_HWDATA(20) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), 
        CoreAHBLite_0_AHBmslave3_HWDATA(19) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), 
        CoreAHBLite_0_AHBmslave3_HWDATA(18) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), 
        CoreAHBLite_0_AHBmslave3_HWDATA(17) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), 
        CoreAHBLite_0_AHBmslave3_HWDATA(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), 
        CoreAHBLite_0_AHBmslave3_HWDATA(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), 
        CoreAHBLite_0_AHBmslave3_HWDATA(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), 
        CoreAHBLite_0_AHBmslave3_HWDATA(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), 
        CoreAHBLite_0_AHBmslave3_HWDATA(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), 
        CoreAHBLite_0_AHBmslave3_HWDATA(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), 
        CoreAHBLite_0_AHBmslave3_HWDATA(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), 
        CoreAHBLite_0_AHBmslave3_HWDATA(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), 
        CoreAHBLite_0_AHBmslave3_HWDATA(8) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), 
        CoreAHBLite_0_AHBmslave3_HWDATA(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(7), 
        CoreAHBLite_0_AHBmslave3_HWDATA(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(6), 
        CoreAHBLite_0_AHBmslave3_HWDATA(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), 
        CoreAHBLite_0_AHBmslave3_HWDATA(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), 
        CoreAHBLite_0_AHBmslave3_HWDATA(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), 
        CoreAHBLite_0_AHBmslave3_HWDATA(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), 
        CoreAHBLite_0_AHBmslave3_HWDATA(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), 
        CoreAHBLite_0_AHBmslave3_HWDATA(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0) => 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0), 
        MASTERADDRINPROG_i_a2_0_a3_0(0) => 
        MASTERADDRINPROG_i_a2_0_a3_0(0), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        M0GATEDHADDR_0 => M0GATEDHADDR(0), M0GATEDHADDR_1 => 
        M0GATEDHADDR(1), M0GATEDHADDR_2 => M0GATEDHADDR(2), 
        M0GATEDHADDR_3 => M0GATEDHADDR(3), M0GATEDHADDR_12 => 
        M0GATEDHADDR(12), M0GATEDHADDR_13 => M0GATEDHADDR(13), 
        M0GATEDHADDR_14 => M0GATEDHADDR(14), M0GATEDHADDR_15 => 
        M0GATEDHADDR(15), M0GATEDHADDR_4 => M0GATEDHADDR(4), 
        M0GATEDHADDR_5 => M0GATEDHADDR(5), M0GATEDHADDR_6 => 
        M0GATEDHADDR(6), M0GATEDHADDR_7 => M0GATEDHADDR(7), 
        M0GATEDHADDR_8 => M0GATEDHADDR(8), M0GATEDHADDR_9 => 
        M0GATEDHADDR(9), M0GATEDHADDR_10 => M0GATEDHADDR(10), 
        M0GATEDHADDR_11 => M0GATEDHADDR(11), MSS_READY => 
        MSS_READY, FAB_CCC_GL0 => FAB_CCC_GL0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, M0GATEDHWRITE => 
        M0GATEDHWRITE, un1_hready_m_xhdl342_1_i_0_o3_2 => 
        un1_hready_m_xhdl342_1_i_0_o3_2, 
        un1_hready_m_xhdl342_1_i_0_o3_3 => 
        un1_hready_m_xhdl342_1_i_0_o3_3, defSlaveSMCurrentState
         => defSlaveSMCurrentState, HREADY_M_iv_i_0 => 
        HREADY_M_iv_i_0, defSlaveSMNextState_m => 
        defSlaveSMNextState_m, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, N_7_i_0 => 
        N_7_i_0, N_25_i_0 => N_25_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_MSS is

    port( xhdl1250_i_m_1                                             : in    std_logic_vector(0 to 0);
          CoreAHBLite_0_AHBmslave3_HRDATA                            : in    std_logic_vector(31 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE    : out   std_logic_vector(1 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : out   std_logic_vector(1 to 1);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : out   std_logic_vector(31 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : in    std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31 : out   std_logic;
          SPI_0_SS0                                                  : inout std_logic := 'Z';
          SPI_0_DO                                                   : out   std_logic;
          SPI_0_DI                                                   : in    std_logic;
          SPI_0_CLK                                                  : inout std_logic := 'Z';
          MMUART_1_TXD                                               : out   std_logic;
          MMUART_1_RXD                                               : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N      : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F           : out   std_logic;
          GPIO_0_M2F_c                                               : out   std_logic;
          HREADY_M_iv_i_0                                            : in    std_logic;
          FAB_CCC_LOCK                                               : in    std_logic;
          FAB_CCC_GL0                                                : in    std_logic
        );

end CertificationSystem_sb_MSS;

architecture DEF_ARCH of CertificationSystem_sb_MSS is 

  component TRIBUFF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component MSS_075

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MGPIO0B_IN                              : in    std_logic := 'U';
          MGPIO10B_IN                             : in    std_logic := 'U';
          MGPIO1B_IN                              : in    std_logic := 'U';
          MGPIO25A_IN                             : in    std_logic := 'U';
          MGPIO26A_IN                             : in    std_logic := 'U';
          MGPIO27A_IN                             : in    std_logic := 'U';
          MGPIO28A_IN                             : in    std_logic := 'U';
          MGPIO29A_IN                             : in    std_logic := 'U';
          MGPIO2B_IN                              : in    std_logic := 'U';
          MGPIO30A_IN                             : in    std_logic := 'U';
          MGPIO31A_IN                             : in    std_logic := 'U';
          MGPIO3B_IN                              : in    std_logic := 'U';
          MGPIO4B_IN                              : in    std_logic := 'U';
          MGPIO5B_IN                              : in    std_logic := 'U';
          MGPIO6B_IN                              : in    std_logic := 'U';
          MGPIO7B_IN                              : in    std_logic := 'U';
          MGPIO8B_IN                              : in    std_logic := 'U';
          MGPIO9B_IN                              : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_CTS_MGPIO13B_IN                 : in    std_logic := 'U';
          MMUART1_DCD_MGPIO16B_IN                 : in    std_logic := 'U';
          MMUART1_DSR_MGPIO14B_IN                 : in    std_logic := 'U';
          MMUART1_DTR_MGPIO12B_IN                 : in    std_logic := 'U';
          MMUART1_RI_MGPIO15B_IN                  : in    std_logic := 'U';
          MMUART1_RTS_MGPIO11B_IN                 : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI0_SS4_MGPIO19A_IN                    : in    std_logic := 'U';
          SPI0_SS5_MGPIO20A_IN                    : in    std_logic := 'U';
          SPI0_SS6_MGPIO21A_IN                    : in    std_logic := 'U';
          SPI0_SS7_MGPIO22A_IN                    : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          USBD_DATA0_IN                           : in    std_logic := 'U';
          USBD_DATA1_IN                           : in    std_logic := 'U';
          USBD_DATA2_IN                           : in    std_logic := 'U';
          USBD_DATA3_IN                           : in    std_logic := 'U';
          USBD_DATA4_IN                           : in    std_logic := 'U';
          USBD_DATA5_IN                           : in    std_logic := 'U';
          USBD_DATA6_IN                           : in    std_logic := 'U';
          USBD_DATA7_MGPIO23B_IN                  : in    std_logic := 'U';
          USBD_DIR_IN                             : in    std_logic := 'U';
          USBD_NXT_IN                             : in    std_logic := 'U';
          USBD_STP_IN                             : in    std_logic := 'U';
          USBD_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MGPIO0B_OUT                             : out   std_logic;
          MGPIO10B_OUT                            : out   std_logic;
          MGPIO1B_OUT                             : out   std_logic;
          MGPIO25A_OUT                            : out   std_logic;
          MGPIO26A_OUT                            : out   std_logic;
          MGPIO27A_OUT                            : out   std_logic;
          MGPIO28A_OUT                            : out   std_logic;
          MGPIO29A_OUT                            : out   std_logic;
          MGPIO2B_OUT                             : out   std_logic;
          MGPIO30A_OUT                            : out   std_logic;
          MGPIO31A_OUT                            : out   std_logic;
          MGPIO3B_OUT                             : out   std_logic;
          MGPIO4B_OUT                             : out   std_logic;
          MGPIO5B_OUT                             : out   std_logic;
          MGPIO6B_OUT                             : out   std_logic;
          MGPIO7B_OUT                             : out   std_logic;
          MGPIO8B_OUT                             : out   std_logic;
          MGPIO9B_OUT                             : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_CTS_MGPIO13B_OUT                : out   std_logic;
          MMUART1_DCD_MGPIO16B_OUT                : out   std_logic;
          MMUART1_DSR_MGPIO14B_OUT                : out   std_logic;
          MMUART1_DTR_MGPIO12B_OUT                : out   std_logic;
          MMUART1_RI_MGPIO15B_OUT                 : out   std_logic;
          MMUART1_RTS_MGPIO11B_OUT                : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI0_SS4_MGPIO19A_OUT                   : out   std_logic;
          SPI0_SS5_MGPIO20A_OUT                   : out   std_logic;
          SPI0_SS6_MGPIO21A_OUT                   : out   std_logic;
          SPI0_SS7_MGPIO22A_OUT                   : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          USBD_DATA0_OUT                          : out   std_logic;
          USBD_DATA1_OUT                          : out   std_logic;
          USBD_DATA2_OUT                          : out   std_logic;
          USBD_DATA3_OUT                          : out   std_logic;
          USBD_DATA4_OUT                          : out   std_logic;
          USBD_DATA5_OUT                          : out   std_logic;
          USBD_DATA6_OUT                          : out   std_logic;
          USBD_DATA7_MGPIO23B_OUT                 : out   std_logic;
          USBD_DIR_OUT                            : out   std_logic;
          USBD_NXT_OUT                            : out   std_logic;
          USBD_STP_OUT                            : out   std_logic;
          USBD_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MGPIO0B_OE                              : out   std_logic;
          MGPIO10B_OE                             : out   std_logic;
          MGPIO1B_OE                              : out   std_logic;
          MGPIO25A_OE                             : out   std_logic;
          MGPIO26A_OE                             : out   std_logic;
          MGPIO27A_OE                             : out   std_logic;
          MGPIO28A_OE                             : out   std_logic;
          MGPIO29A_OE                             : out   std_logic;
          MGPIO2B_OE                              : out   std_logic;
          MGPIO30A_OE                             : out   std_logic;
          MGPIO31A_OE                             : out   std_logic;
          MGPIO3B_OE                              : out   std_logic;
          MGPIO4B_OE                              : out   std_logic;
          MGPIO5B_OE                              : out   std_logic;
          MGPIO6B_OE                              : out   std_logic;
          MGPIO7B_OE                              : out   std_logic;
          MGPIO8B_OE                              : out   std_logic;
          MGPIO9B_OE                              : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_CTS_MGPIO13B_OE                 : out   std_logic;
          MMUART1_DCD_MGPIO16B_OE                 : out   std_logic;
          MMUART1_DSR_MGPIO14B_OE                 : out   std_logic;
          MMUART1_DTR_MGPIO12B_OE                 : out   std_logic;
          MMUART1_RI_MGPIO15B_OE                  : out   std_logic;
          MMUART1_RTS_MGPIO11B_OE                 : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI0_SS4_MGPIO19A_OE                    : out   std_logic;
          SPI0_SS5_MGPIO20A_OE                    : out   std_logic;
          SPI0_SS6_MGPIO21A_OE                    : out   std_logic;
          SPI0_SS7_MGPIO22A_OE                    : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic;
          USBD_DATA0_OE                           : out   std_logic;
          USBD_DATA1_OE                           : out   std_logic;
          USBD_DATA2_OE                           : out   std_logic;
          USBD_DATA3_OE                           : out   std_logic;
          USBD_DATA4_OE                           : out   std_logic;
          USBD_DATA5_OE                           : out   std_logic;
          USBD_DATA6_OE                           : out   std_logic;
          USBD_DATA7_MGPIO23B_OE                  : out   std_logic;
          USBD_DIR_OE                             : out   std_logic;
          USBD_NXT_OE                             : out   std_logic;
          USBD_STP_OE                             : out   std_logic;
          USBD_XCLK_OE                            : out   std_logic
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

    signal SPI_0_SS0_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI_0_DI_PAD_Y, SPI_0_CLK_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        MMUART_1_RXD_PAD_Y, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[31]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[30]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[29]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[28]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[27]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[26]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[25]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[24]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[23]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[22]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[21]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[20]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[19]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[18]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[17]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[16]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[15]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[14]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[13]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[12]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[11]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[10]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[9]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[8]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[7]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[6]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[5]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[4]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[3]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[2]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[1]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[0]\, VCC_net_1, 
        GND_net_1 : std_logic;
    signal nc228, nc203, nc265, nc216, nc194, nc151, nc23, nc175, 
        nc250, nc58, nc116, nc74, nc133, nc238, nc167, nc84, nc39, 
        nc72, nc256, nc212, nc205, nc82, nc145, nc181, nc160, 
        nc57, nc156, nc280, nc125, nc211, nc73, nc107, nc66, nc83, 
        nc9, nc252, nc171, nc54, nc286, nc307, nc135, nc41, nc100, 
        nc270, nc52, nc251, nc186, nc29, nc269, nc118, nc60, 
        nc141, nc311, nc276, nc193, nc214, nc298, nc282, nc240, 
        nc45, nc53, nc121, nc176, nc220, nc158, nc281, nc209, 
        nc246, nc162, nc11, nc272, nc131, nc254, nc267, nc96, 
        nc79, nc226, nc146, nc230, nc89, nc119, nc48, nc271, 
        nc213, nc300, nc126, nc195, nc188, nc242, nc15, nc308, 
        nc236, nc102, nc304, nc3, nc207, nc47, nc90, nc284, nc222, 
        nc159, nc136, nc241, nc253, nc178, nc306, nc215, nc59, 
        nc221, nc232, nc274, nc18, nc44, nc117, nc189, nc164, 
        nc148, nc42, nc231, nc191, nc255, nc283, nc317, nc290, 
        nc17, nc2, nc302, nc110, nc128, nc244, nc321, nc43, nc179, 
        nc157, nc36, nc224, nc296, nc273, nc61, nc104, nc138, 
        nc14, nc285, nc303, nc150, nc196, nc234, nc149, nc12, 
        nc219, nc30, nc243, nc187, nc65, nc7, nc292, nc129, nc275, 
        nc8, nc223, nc13, nc305, nc180, nc26, nc291, nc177, nc139, 
        nc310, nc259, nc245, nc233, nc163, nc318, nc268, nc112, 
        nc68, nc49, nc314, nc217, nc170, nc91, nc225, nc5, nc20, 
        nc198, nc147, nc316, nc67, nc289, nc294, nc152, nc127, 
        nc103, nc235, nc76, nc208, nc140, nc257, nc86, nc95, 
        nc120, nc165, nc279, nc137, nc64, nc19, nc312, nc70, 
        nc182, nc62, nc199, nc80, nc130, nc287, nc98, nc293, 
        nc249, nc114, nc56, nc105, nc63, nc313, nc309, nc172, 
        nc229, nc277, nc97, nc161, nc31, nc295, nc154, nc50, 
        nc260, nc239, nc142, nc320, nc315, nc247, nc94, nc197, 
        nc122, nc266, nc35, nc4, nc227, nc92, nc101, nc184, nc200, 
        nc190, nc166, nc132, nc21, nc237, nc93, nc262, nc69, 
        nc206, nc174, nc38, nc113, nc218, nc106, nc261, nc25, nc1, 
        nc299, nc37, nc202, nc144, nc153, nc46, nc258, nc71, 
        nc124, nc81, nc201, nc168, nc34, nc28, nc115, nc264, 
        nc192, nc319, nc134, nc32, nc40, nc297, nc99, nc75, nc183, 
        nc288, nc85, nc27, nc108, nc16, nc155, nc51, nc301, nc33, 
        nc204, nc173, nc278, nc169, nc78, nc263, nc24, nc88, 
        nc111, nc55, nc10, nc22, nc210, nc185, nc143, nc248, nc77, 
        nc6, nc109, nc87, nc123 : std_logic;

begin 


    MMUART_1_TXD_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, PAD
         => MMUART_1_TXD);
    
    MSS_ADLIB_INST_RNO_20 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(21), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[21]\);
    
    MSS_ADLIB_INST_RNO_23 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(24), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[24]\);
    
    MSS_ADLIB_INST_RNO_29 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(30), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[30]\);
    
    MSS_ADLIB_INST_RNO_21 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(22), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[22]\);
    
    MSS_ADLIB_INST_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(0), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[0]\);
    
    MSS_ADLIB_INST_RNO_22 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(23), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[23]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    MSS_ADLIB_INST_RNO_27 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(28), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[28]\);
    
    MSS_ADLIB_INST_RNO_10 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(11), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[11]\);
    
    MSS_ADLIB_INST_RNO_13 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(14), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[14]\);
    
    MSS_ADLIB_INST_RNO_19 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(20), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[20]\);
    
    MSS_ADLIB_INST_RNO_11 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(12), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[12]\);
    
    SPI_0_DO_PAD : TRIBUFF
      port map(D => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        E => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, PAD => 
        SPI_0_DO);
    
    MSS_ADLIB_INST_RNO_12 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(13), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[13]\);
    
    MSS_ADLIB_INST_RNO_2 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(3), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[3]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    MSS_ADLIB_INST_RNO_4 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(5), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[5]\);
    
    SPI_0_DI_PAD : INBUF
      port map(PAD => SPI_0_DI, Y => SPI_0_DI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_17 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(18), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[18]\);
    
    MSS_ADLIB_INST_RNO_7 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(8), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[8]\);
    
    MSS_ADLIB_INST : MSS_075

              generic map(INIT => "00" & x"0000000000000000000000000000036100080000000000000000000000000000000000000000000000000000000000001203610000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C35C00000000609300000003FFFFE4000000000000100000000F0E11C00000182DF34010842108421000001FE34001FF8000000400000000000451007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem", RTC_MAIN_XTL_FREQ => 0.0,
         DDR_CLK_FREQ => 50.0)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => OPEN, CAN_TX_EBL_MGPIO4A_H2F_A
         => OPEN, CAN_TX_EBL_MGPIO4A_H2F_B => OPEN, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => OPEN, CLK_CONFIG_APB => OPEN, COMMS_INT => OPEN, 
        CONFIG_PRESET_N => 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        EDAC_ERROR(7) => nc228, EDAC_ERROR(6) => nc203, 
        EDAC_ERROR(5) => nc265, EDAC_ERROR(4) => nc216, 
        EDAC_ERROR(3) => nc194, EDAC_ERROR(2) => nc151, 
        EDAC_ERROR(1) => nc23, EDAC_ERROR(0) => nc175, 
        F_FM0_RDATA(31) => nc250, F_FM0_RDATA(30) => nc58, 
        F_FM0_RDATA(29) => nc116, F_FM0_RDATA(28) => nc74, 
        F_FM0_RDATA(27) => nc133, F_FM0_RDATA(26) => nc238, 
        F_FM0_RDATA(25) => nc167, F_FM0_RDATA(24) => nc84, 
        F_FM0_RDATA(23) => nc39, F_FM0_RDATA(22) => nc72, 
        F_FM0_RDATA(21) => nc256, F_FM0_RDATA(20) => nc212, 
        F_FM0_RDATA(19) => nc205, F_FM0_RDATA(18) => nc82, 
        F_FM0_RDATA(17) => nc145, F_FM0_RDATA(16) => nc181, 
        F_FM0_RDATA(15) => nc160, F_FM0_RDATA(14) => nc57, 
        F_FM0_RDATA(13) => nc156, F_FM0_RDATA(12) => nc280, 
        F_FM0_RDATA(11) => nc125, F_FM0_RDATA(10) => nc211, 
        F_FM0_RDATA(9) => nc73, F_FM0_RDATA(8) => nc107, 
        F_FM0_RDATA(7) => nc66, F_FM0_RDATA(6) => nc83, 
        F_FM0_RDATA(5) => nc9, F_FM0_RDATA(4) => nc252, 
        F_FM0_RDATA(3) => nc171, F_FM0_RDATA(2) => nc54, 
        F_FM0_RDATA(1) => nc286, F_FM0_RDATA(0) => nc307, 
        F_FM0_READYOUT => OPEN, F_FM0_RESP => OPEN, 
        F_HM0_ADDR(31) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        F_HM0_ADDR(30) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        F_HM0_ADDR(29) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        F_HM0_ADDR(28) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        F_HM0_ADDR(27) => nc135, F_HM0_ADDR(26) => nc41, 
        F_HM0_ADDR(25) => nc100, F_HM0_ADDR(24) => nc270, 
        F_HM0_ADDR(23) => nc52, F_HM0_ADDR(22) => nc251, 
        F_HM0_ADDR(21) => nc186, F_HM0_ADDR(20) => nc29, 
        F_HM0_ADDR(19) => nc269, F_HM0_ADDR(18) => nc118, 
        F_HM0_ADDR(17) => nc60, F_HM0_ADDR(16) => nc141, 
        F_HM0_ADDR(15) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15, 
        F_HM0_ADDR(14) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14, 
        F_HM0_ADDR(13) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13, 
        F_HM0_ADDR(12) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12, 
        F_HM0_ADDR(11) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11, 
        F_HM0_ADDR(10) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10, 
        F_HM0_ADDR(9) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9, 
        F_HM0_ADDR(8) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        F_HM0_ADDR(7) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7, 
        F_HM0_ADDR(6) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        F_HM0_ADDR(5) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        F_HM0_ADDR(4) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        F_HM0_ADDR(3) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        F_HM0_ADDR(2) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        F_HM0_ADDR(1) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        F_HM0_ADDR(0) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        F_HM0_ENABLE => OPEN, F_HM0_SEL => OPEN, F_HM0_SIZE(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1), 
        F_HM0_SIZE(0) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0), 
        F_HM0_TRANS1 => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        F_HM0_WDATA(31) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        F_HM0_WDATA(30) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        F_HM0_WDATA(29) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        F_HM0_WDATA(28) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        F_HM0_WDATA(27) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        F_HM0_WDATA(26) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        F_HM0_WDATA(25) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        F_HM0_WDATA(24) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        F_HM0_WDATA(23) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        F_HM0_WDATA(22) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        F_HM0_WDATA(21) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        F_HM0_WDATA(20) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        F_HM0_WDATA(19) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        F_HM0_WDATA(18) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        F_HM0_WDATA(17) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        F_HM0_WDATA(16) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        F_HM0_WDATA(15) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        F_HM0_WDATA(14) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        F_HM0_WDATA(13) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        F_HM0_WDATA(12) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        F_HM0_WDATA(11) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        F_HM0_WDATA(10) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        F_HM0_WDATA(9) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        F_HM0_WDATA(8) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        F_HM0_WDATA(7) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        F_HM0_WDATA(6) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        F_HM0_WDATA(5) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        F_HM0_WDATA(4) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        F_HM0_WDATA(3) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        F_HM0_WDATA(2) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        F_HM0_WDATA(1) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        F_HM0_WDATA(0) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        F_HM0_WRITE => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        FAB_CHRGVBUS => OPEN, FAB_DISCHRGVBUS => OPEN, 
        FAB_DMPULLDOWN => OPEN, FAB_DPPULLDOWN => OPEN, 
        FAB_DRVVBUS => OPEN, FAB_IDPULLUP => OPEN, FAB_OPMODE(1)
         => nc311, FAB_OPMODE(0) => nc276, FAB_SUSPENDM => OPEN, 
        FAB_TERMSEL => OPEN, FAB_TXVALID => OPEN, FAB_VCONTROL(3)
         => nc193, FAB_VCONTROL(2) => nc214, FAB_VCONTROL(1) => 
        nc298, FAB_VCONTROL(0) => nc282, FAB_VCONTROLLOADM => 
        OPEN, FAB_XCVRSEL(1) => nc240, FAB_XCVRSEL(0) => nc45, 
        FAB_XDATAOUT(7) => nc53, FAB_XDATAOUT(6) => nc121, 
        FAB_XDATAOUT(5) => nc176, FAB_XDATAOUT(4) => nc220, 
        FAB_XDATAOUT(3) => nc158, FAB_XDATAOUT(2) => nc281, 
        FAB_XDATAOUT(1) => nc209, FAB_XDATAOUT(0) => nc246, 
        FACC_GLMUX_SEL => OPEN, FIC32_0_MASTER(1) => nc162, 
        FIC32_0_MASTER(0) => nc11, FIC32_1_MASTER(1) => nc272, 
        FIC32_1_MASTER(0) => nc131, FPGA_RESET_N => 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, GTX_CLK
         => OPEN, H2F_INTERRUPT(15) => nc254, H2F_INTERRUPT(14)
         => nc267, H2F_INTERRUPT(13) => nc96, H2F_INTERRUPT(12)
         => nc79, H2F_INTERRUPT(11) => nc226, H2F_INTERRUPT(10)
         => nc146, H2F_INTERRUPT(9) => nc230, H2F_INTERRUPT(8)
         => nc89, H2F_INTERRUPT(7) => nc119, H2F_INTERRUPT(6) => 
        nc48, H2F_INTERRUPT(5) => nc271, H2F_INTERRUPT(4) => 
        nc213, H2F_INTERRUPT(3) => nc300, H2F_INTERRUPT(2) => 
        nc126, H2F_INTERRUPT(1) => nc195, H2F_INTERRUPT(0) => 
        nc188, H2F_NMI => OPEN, H2FCALIB => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_A => OPEN, I2C0_SCL_MGPIO31B_H2F_B
         => OPEN, I2C0_SDA_MGPIO30B_H2F_A => OPEN, 
        I2C0_SDA_MGPIO30B_H2F_B => OPEN, I2C1_SCL_MGPIO1A_H2F_A
         => OPEN, I2C1_SCL_MGPIO1A_H2F_B => OPEN, 
        I2C1_SDA_MGPIO0A_H2F_A => OPEN, I2C1_SDA_MGPIO0A_H2F_B
         => GPIO_0_M2F_c, MDCF => OPEN, MDOENF => OPEN, MDOF => 
        OPEN, MMUART0_CTS_MGPIO19B_H2F_A => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => OPEN, MPLL_LOCK => OPEN, 
        PER2_FABRIC_PADDR(15) => nc242, PER2_FABRIC_PADDR(14) => 
        nc15, PER2_FABRIC_PADDR(13) => nc308, 
        PER2_FABRIC_PADDR(12) => nc236, PER2_FABRIC_PADDR(11) => 
        nc102, PER2_FABRIC_PADDR(10) => nc304, 
        PER2_FABRIC_PADDR(9) => nc3, PER2_FABRIC_PADDR(8) => 
        nc207, PER2_FABRIC_PADDR(7) => nc47, PER2_FABRIC_PADDR(6)
         => nc90, PER2_FABRIC_PADDR(5) => nc284, 
        PER2_FABRIC_PADDR(4) => nc222, PER2_FABRIC_PADDR(3) => 
        nc159, PER2_FABRIC_PADDR(2) => nc136, PER2_FABRIC_PENABLE
         => OPEN, PER2_FABRIC_PSEL => OPEN, 
        PER2_FABRIC_PWDATA(31) => nc241, PER2_FABRIC_PWDATA(30)
         => nc253, PER2_FABRIC_PWDATA(29) => nc178, 
        PER2_FABRIC_PWDATA(28) => nc306, PER2_FABRIC_PWDATA(27)
         => nc215, PER2_FABRIC_PWDATA(26) => nc59, 
        PER2_FABRIC_PWDATA(25) => nc221, PER2_FABRIC_PWDATA(24)
         => nc232, PER2_FABRIC_PWDATA(23) => nc274, 
        PER2_FABRIC_PWDATA(22) => nc18, PER2_FABRIC_PWDATA(21)
         => nc44, PER2_FABRIC_PWDATA(20) => nc117, 
        PER2_FABRIC_PWDATA(19) => nc189, PER2_FABRIC_PWDATA(18)
         => nc164, PER2_FABRIC_PWDATA(17) => nc148, 
        PER2_FABRIC_PWDATA(16) => nc42, PER2_FABRIC_PWDATA(15)
         => nc231, PER2_FABRIC_PWDATA(14) => nc191, 
        PER2_FABRIC_PWDATA(13) => nc255, PER2_FABRIC_PWDATA(12)
         => nc283, PER2_FABRIC_PWDATA(11) => nc317, 
        PER2_FABRIC_PWDATA(10) => nc290, PER2_FABRIC_PWDATA(9)
         => nc17, PER2_FABRIC_PWDATA(8) => nc2, 
        PER2_FABRIC_PWDATA(7) => nc302, PER2_FABRIC_PWDATA(6) => 
        nc110, PER2_FABRIC_PWDATA(5) => nc128, 
        PER2_FABRIC_PWDATA(4) => nc244, PER2_FABRIC_PWDATA(3) => 
        nc321, PER2_FABRIC_PWDATA(2) => nc43, 
        PER2_FABRIC_PWDATA(1) => nc179, PER2_FABRIC_PWDATA(0) => 
        nc157, PER2_FABRIC_PWRITE => OPEN, RTC_MATCH => OPEN, 
        SLEEPDEEP => OPEN, SLEEPHOLDACK => OPEN, SLEEPING => OPEN, 
        SMBALERT_NO0 => OPEN, SMBALERT_NO1 => OPEN, SMBSUS_NO0
         => OPEN, SMBSUS_NO1 => OPEN, SPI0_CLK_OUT => OPEN, 
        SPI0_SDI_MGPIO5A_H2F_A => OPEN, SPI0_SDI_MGPIO5A_H2F_B
         => OPEN, SPI0_SDO_MGPIO6A_H2F_A => OPEN, 
        SPI0_SDO_MGPIO6A_H2F_B => OPEN, SPI0_SS0_MGPIO7A_H2F_A
         => OPEN, SPI0_SS0_MGPIO7A_H2F_B => OPEN, 
        SPI0_SS1_MGPIO8A_H2F_A => OPEN, SPI0_SS1_MGPIO8A_H2F_B
         => OPEN, SPI0_SS2_MGPIO9A_H2F_A => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_B => OPEN, SPI0_SS3_MGPIO10A_H2F_A
         => OPEN, SPI0_SS3_MGPIO10A_H2F_B => OPEN, 
        SPI0_SS4_MGPIO19A_H2F_A => OPEN, SPI0_SS5_MGPIO20A_H2F_A
         => OPEN, SPI0_SS6_MGPIO21A_H2F_A => OPEN, 
        SPI0_SS7_MGPIO22A_H2F_A => OPEN, SPI1_CLK_OUT => OPEN, 
        SPI1_SDI_MGPIO11A_H2F_A => OPEN, SPI1_SDI_MGPIO11A_H2F_B
         => OPEN, SPI1_SDO_MGPIO12A_H2F_A => OPEN, 
        SPI1_SDO_MGPIO12A_H2F_B => OPEN, SPI1_SS0_MGPIO13A_H2F_A
         => OPEN, SPI1_SS0_MGPIO13A_H2F_B => OPEN, 
        SPI1_SS1_MGPIO14A_H2F_A => OPEN, SPI1_SS1_MGPIO14A_H2F_B
         => OPEN, SPI1_SS2_MGPIO15A_H2F_A => OPEN, 
        SPI1_SS2_MGPIO15A_H2F_B => OPEN, SPI1_SS3_MGPIO16A_H2F_A
         => OPEN, SPI1_SS3_MGPIO16A_H2F_B => OPEN, 
        SPI1_SS4_MGPIO17A_H2F_A => OPEN, SPI1_SS5_MGPIO18A_H2F_A
         => OPEN, SPI1_SS6_MGPIO23A_H2F_A => OPEN, 
        SPI1_SS7_MGPIO24A_H2F_A => OPEN, TCGF(9) => nc36, TCGF(8)
         => nc224, TCGF(7) => nc296, TCGF(6) => nc273, TCGF(5)
         => nc61, TCGF(4) => nc104, TCGF(3) => nc138, TCGF(2) => 
        nc14, TCGF(1) => nc285, TCGF(0) => nc303, TRACECLK => 
        OPEN, TRACEDATA(3) => nc150, TRACEDATA(2) => nc196, 
        TRACEDATA(1) => nc234, TRACEDATA(0) => nc149, TX_CLK => 
        OPEN, TX_ENF => OPEN, TX_ERRF => OPEN, TXCTL_EN_RIF => 
        OPEN, TXD_RIF(3) => nc12, TXD_RIF(2) => nc219, TXD_RIF(1)
         => nc30, TXD_RIF(0) => nc243, TXDF(7) => nc187, TXDF(6)
         => nc65, TXDF(5) => nc7, TXDF(4) => nc292, TXDF(3) => 
        nc129, TXDF(2) => nc275, TXDF(1) => nc8, TXDF(0) => nc223, 
        TXEV => OPEN, WDOGTIMEOUT => OPEN, F_ARREADY_HREADYOUT1
         => OPEN, F_AWREADY_HREADYOUT0 => OPEN, F_BID(3) => nc13, 
        F_BID(2) => nc305, F_BID(1) => nc180, F_BID(0) => nc26, 
        F_BRESP_HRESP0(1) => nc291, F_BRESP_HRESP0(0) => nc177, 
        F_BVALID => OPEN, F_RDATA_HRDATA01(63) => nc139, 
        F_RDATA_HRDATA01(62) => nc310, F_RDATA_HRDATA01(61) => 
        nc259, F_RDATA_HRDATA01(60) => nc245, 
        F_RDATA_HRDATA01(59) => nc233, F_RDATA_HRDATA01(58) => 
        nc163, F_RDATA_HRDATA01(57) => nc318, 
        F_RDATA_HRDATA01(56) => nc268, F_RDATA_HRDATA01(55) => 
        nc112, F_RDATA_HRDATA01(54) => nc68, F_RDATA_HRDATA01(53)
         => nc49, F_RDATA_HRDATA01(52) => nc314, 
        F_RDATA_HRDATA01(51) => nc217, F_RDATA_HRDATA01(50) => 
        nc170, F_RDATA_HRDATA01(49) => nc91, F_RDATA_HRDATA01(48)
         => nc225, F_RDATA_HRDATA01(47) => nc5, 
        F_RDATA_HRDATA01(46) => nc20, F_RDATA_HRDATA01(45) => 
        nc198, F_RDATA_HRDATA01(44) => nc147, 
        F_RDATA_HRDATA01(43) => nc316, F_RDATA_HRDATA01(42) => 
        nc67, F_RDATA_HRDATA01(41) => nc289, F_RDATA_HRDATA01(40)
         => nc294, F_RDATA_HRDATA01(39) => nc152, 
        F_RDATA_HRDATA01(38) => nc127, F_RDATA_HRDATA01(37) => 
        nc103, F_RDATA_HRDATA01(36) => nc235, 
        F_RDATA_HRDATA01(35) => nc76, F_RDATA_HRDATA01(34) => 
        nc208, F_RDATA_HRDATA01(33) => nc140, 
        F_RDATA_HRDATA01(32) => nc257, F_RDATA_HRDATA01(31) => 
        nc86, F_RDATA_HRDATA01(30) => nc95, F_RDATA_HRDATA01(29)
         => nc120, F_RDATA_HRDATA01(28) => nc165, 
        F_RDATA_HRDATA01(27) => nc279, F_RDATA_HRDATA01(26) => 
        nc137, F_RDATA_HRDATA01(25) => nc64, F_RDATA_HRDATA01(24)
         => nc19, F_RDATA_HRDATA01(23) => nc312, 
        F_RDATA_HRDATA01(22) => nc70, F_RDATA_HRDATA01(21) => 
        nc182, F_RDATA_HRDATA01(20) => nc62, F_RDATA_HRDATA01(19)
         => nc199, F_RDATA_HRDATA01(18) => nc80, 
        F_RDATA_HRDATA01(17) => nc130, F_RDATA_HRDATA01(16) => 
        nc287, F_RDATA_HRDATA01(15) => nc98, F_RDATA_HRDATA01(14)
         => nc293, F_RDATA_HRDATA01(13) => nc249, 
        F_RDATA_HRDATA01(12) => nc114, F_RDATA_HRDATA01(11) => 
        nc56, F_RDATA_HRDATA01(10) => nc105, F_RDATA_HRDATA01(9)
         => nc63, F_RDATA_HRDATA01(8) => nc313, 
        F_RDATA_HRDATA01(7) => nc309, F_RDATA_HRDATA01(6) => 
        nc172, F_RDATA_HRDATA01(5) => nc229, F_RDATA_HRDATA01(4)
         => nc277, F_RDATA_HRDATA01(3) => nc97, 
        F_RDATA_HRDATA01(2) => nc161, F_RDATA_HRDATA01(1) => nc31, 
        F_RDATA_HRDATA01(0) => nc295, F_RID(3) => nc154, F_RID(2)
         => nc50, F_RID(1) => nc260, F_RID(0) => nc239, F_RLAST
         => OPEN, F_RRESP_HRESP1(1) => nc142, F_RRESP_HRESP1(0)
         => nc320, F_RVALID => OPEN, F_WREADY => OPEN, 
        MDDR_FABRIC_PRDATA(15) => nc315, MDDR_FABRIC_PRDATA(14)
         => nc247, MDDR_FABRIC_PRDATA(13) => nc94, 
        MDDR_FABRIC_PRDATA(12) => nc197, MDDR_FABRIC_PRDATA(11)
         => nc122, MDDR_FABRIC_PRDATA(10) => nc266, 
        MDDR_FABRIC_PRDATA(9) => nc35, MDDR_FABRIC_PRDATA(8) => 
        nc4, MDDR_FABRIC_PRDATA(7) => nc227, 
        MDDR_FABRIC_PRDATA(6) => nc92, MDDR_FABRIC_PRDATA(5) => 
        nc101, MDDR_FABRIC_PRDATA(4) => nc184, 
        MDDR_FABRIC_PRDATA(3) => nc200, MDDR_FABRIC_PRDATA(2) => 
        nc190, MDDR_FABRIC_PRDATA(1) => nc166, 
        MDDR_FABRIC_PRDATA(0) => nc132, MDDR_FABRIC_PREADY => 
        OPEN, MDDR_FABRIC_PSLVERR => OPEN, CAN_RXBUS_F2H_SCP => 
        VCC_net_1, CAN_TX_EBL_F2H_SCP => VCC_net_1, 
        CAN_TXBUS_F2H_SCP => VCC_net_1, COLF => VCC_net_1, CRSF
         => VCC_net_1, F2_DMAREADY(1) => VCC_net_1, 
        F2_DMAREADY(0) => VCC_net_1, F2H_INTERRUPT(15) => 
        GND_net_1, F2H_INTERRUPT(14) => GND_net_1, 
        F2H_INTERRUPT(13) => GND_net_1, F2H_INTERRUPT(12) => 
        GND_net_1, F2H_INTERRUPT(11) => GND_net_1, 
        F2H_INTERRUPT(10) => GND_net_1, F2H_INTERRUPT(9) => 
        GND_net_1, F2H_INTERRUPT(8) => GND_net_1, 
        F2H_INTERRUPT(7) => GND_net_1, F2H_INTERRUPT(6) => 
        GND_net_1, F2H_INTERRUPT(5) => GND_net_1, 
        F2H_INTERRUPT(4) => GND_net_1, F2H_INTERRUPT(3) => 
        GND_net_1, F2H_INTERRUPT(2) => GND_net_1, 
        F2H_INTERRUPT(1) => GND_net_1, F2H_INTERRUPT(0) => 
        GND_net_1, F2HCALIB => VCC_net_1, F_DMAREADY(1) => 
        VCC_net_1, F_DMAREADY(0) => VCC_net_1, F_FM0_ADDR(31) => 
        GND_net_1, F_FM0_ADDR(30) => GND_net_1, F_FM0_ADDR(29)
         => GND_net_1, F_FM0_ADDR(28) => GND_net_1, 
        F_FM0_ADDR(27) => GND_net_1, F_FM0_ADDR(26) => GND_net_1, 
        F_FM0_ADDR(25) => GND_net_1, F_FM0_ADDR(24) => GND_net_1, 
        F_FM0_ADDR(23) => GND_net_1, F_FM0_ADDR(22) => GND_net_1, 
        F_FM0_ADDR(21) => GND_net_1, F_FM0_ADDR(20) => GND_net_1, 
        F_FM0_ADDR(19) => GND_net_1, F_FM0_ADDR(18) => GND_net_1, 
        F_FM0_ADDR(17) => GND_net_1, F_FM0_ADDR(16) => GND_net_1, 
        F_FM0_ADDR(15) => GND_net_1, F_FM0_ADDR(14) => GND_net_1, 
        F_FM0_ADDR(13) => GND_net_1, F_FM0_ADDR(12) => GND_net_1, 
        F_FM0_ADDR(11) => GND_net_1, F_FM0_ADDR(10) => GND_net_1, 
        F_FM0_ADDR(9) => GND_net_1, F_FM0_ADDR(8) => GND_net_1, 
        F_FM0_ADDR(7) => GND_net_1, F_FM0_ADDR(6) => GND_net_1, 
        F_FM0_ADDR(5) => GND_net_1, F_FM0_ADDR(4) => GND_net_1, 
        F_FM0_ADDR(3) => GND_net_1, F_FM0_ADDR(2) => GND_net_1, 
        F_FM0_ADDR(1) => GND_net_1, F_FM0_ADDR(0) => GND_net_1, 
        F_FM0_ENABLE => GND_net_1, F_FM0_MASTLOCK => GND_net_1, 
        F_FM0_READY => VCC_net_1, F_FM0_SEL => GND_net_1, 
        F_FM0_SIZE(1) => GND_net_1, F_FM0_SIZE(0) => GND_net_1, 
        F_FM0_TRANS1 => GND_net_1, F_FM0_WDATA(31) => GND_net_1, 
        F_FM0_WDATA(30) => GND_net_1, F_FM0_WDATA(29) => 
        GND_net_1, F_FM0_WDATA(28) => GND_net_1, F_FM0_WDATA(27)
         => GND_net_1, F_FM0_WDATA(26) => GND_net_1, 
        F_FM0_WDATA(25) => GND_net_1, F_FM0_WDATA(24) => 
        GND_net_1, F_FM0_WDATA(23) => GND_net_1, F_FM0_WDATA(22)
         => GND_net_1, F_FM0_WDATA(21) => GND_net_1, 
        F_FM0_WDATA(20) => GND_net_1, F_FM0_WDATA(19) => 
        GND_net_1, F_FM0_WDATA(18) => GND_net_1, F_FM0_WDATA(17)
         => GND_net_1, F_FM0_WDATA(16) => GND_net_1, 
        F_FM0_WDATA(15) => GND_net_1, F_FM0_WDATA(14) => 
        GND_net_1, F_FM0_WDATA(13) => GND_net_1, F_FM0_WDATA(12)
         => GND_net_1, F_FM0_WDATA(11) => GND_net_1, 
        F_FM0_WDATA(10) => GND_net_1, F_FM0_WDATA(9) => GND_net_1, 
        F_FM0_WDATA(8) => GND_net_1, F_FM0_WDATA(7) => GND_net_1, 
        F_FM0_WDATA(6) => GND_net_1, F_FM0_WDATA(5) => GND_net_1, 
        F_FM0_WDATA(4) => GND_net_1, F_FM0_WDATA(3) => GND_net_1, 
        F_FM0_WDATA(2) => GND_net_1, F_FM0_WDATA(1) => GND_net_1, 
        F_FM0_WDATA(0) => GND_net_1, F_FM0_WRITE => GND_net_1, 
        F_HM0_RDATA(31) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[31]\, F_HM0_RDATA(30)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[30]\, 
        F_HM0_RDATA(29) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[29]\, F_HM0_RDATA(28)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[28]\, 
        F_HM0_RDATA(27) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[27]\, F_HM0_RDATA(26)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[26]\, 
        F_HM0_RDATA(25) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[25]\, F_HM0_RDATA(24)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[24]\, 
        F_HM0_RDATA(23) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[23]\, F_HM0_RDATA(22)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[22]\, 
        F_HM0_RDATA(21) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[21]\, F_HM0_RDATA(20)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[20]\, 
        F_HM0_RDATA(19) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[19]\, F_HM0_RDATA(18)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[18]\, 
        F_HM0_RDATA(17) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[17]\, F_HM0_RDATA(16)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[16]\, 
        F_HM0_RDATA(15) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[15]\, F_HM0_RDATA(14)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[14]\, 
        F_HM0_RDATA(13) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[13]\, F_HM0_RDATA(12)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[12]\, 
        F_HM0_RDATA(11) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[11]\, F_HM0_RDATA(10)
         => \CoreAHBLite_0_AHBmslave3_HRDATA_m[10]\, 
        F_HM0_RDATA(9) => \CoreAHBLite_0_AHBmslave3_HRDATA_m[9]\, 
        F_HM0_RDATA(8) => \CoreAHBLite_0_AHBmslave3_HRDATA_m[8]\, 
        F_HM0_RDATA(7) => \CoreAHBLite_0_AHBmslave3_HRDATA_m[7]\, 
        F_HM0_RDATA(6) => \CoreAHBLite_0_AHBmslave3_HRDATA_m[6]\, 
        F_HM0_RDATA(5) => \CoreAHBLite_0_AHBmslave3_HRDATA_m[5]\, 
        F_HM0_RDATA(4) => \CoreAHBLite_0_AHBmslave3_HRDATA_m[4]\, 
        F_HM0_RDATA(3) => \CoreAHBLite_0_AHBmslave3_HRDATA_m[3]\, 
        F_HM0_RDATA(2) => \CoreAHBLite_0_AHBmslave3_HRDATA_m[2]\, 
        F_HM0_RDATA(1) => \CoreAHBLite_0_AHBmslave3_HRDATA_m[1]\, 
        F_HM0_RDATA(0) => \CoreAHBLite_0_AHBmslave3_HRDATA_m[0]\, 
        F_HM0_READY => HREADY_M_iv_i_0, F_HM0_RESP => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        FAB_AVALID => VCC_net_1, FAB_HOSTDISCON => VCC_net_1, 
        FAB_IDDIG => VCC_net_1, FAB_LINESTATE(1) => VCC_net_1, 
        FAB_LINESTATE(0) => VCC_net_1, FAB_M3_RESET_N => 
        VCC_net_1, FAB_PLL_LOCK => FAB_CCC_LOCK, FAB_RXACTIVE => 
        VCC_net_1, FAB_RXERROR => VCC_net_1, FAB_RXVALID => 
        VCC_net_1, FAB_RXVALIDH => GND_net_1, FAB_SESSEND => 
        VCC_net_1, FAB_TXREADY => VCC_net_1, FAB_VBUSVALID => 
        VCC_net_1, FAB_VSTATUS(7) => VCC_net_1, FAB_VSTATUS(6)
         => VCC_net_1, FAB_VSTATUS(5) => VCC_net_1, 
        FAB_VSTATUS(4) => VCC_net_1, FAB_VSTATUS(3) => VCC_net_1, 
        FAB_VSTATUS(2) => VCC_net_1, FAB_VSTATUS(1) => VCC_net_1, 
        FAB_VSTATUS(0) => VCC_net_1, FAB_XDATAIN(7) => VCC_net_1, 
        FAB_XDATAIN(6) => VCC_net_1, FAB_XDATAIN(5) => VCC_net_1, 
        FAB_XDATAIN(4) => VCC_net_1, FAB_XDATAIN(3) => VCC_net_1, 
        FAB_XDATAIN(2) => VCC_net_1, FAB_XDATAIN(1) => VCC_net_1, 
        FAB_XDATAIN(0) => VCC_net_1, GTX_CLKPF => VCC_net_1, 
        I2C0_BCLK => VCC_net_1, I2C0_SCL_F2H_SCP => VCC_net_1, 
        I2C0_SDA_F2H_SCP => VCC_net_1, I2C1_BCLK => VCC_net_1, 
        I2C1_SCL_F2H_SCP => VCC_net_1, I2C1_SDA_F2H_SCP => 
        VCC_net_1, MDIF => VCC_net_1, MGPIO0A_F2H_GPIN => 
        VCC_net_1, MGPIO10A_F2H_GPIN => VCC_net_1, 
        MGPIO11A_F2H_GPIN => VCC_net_1, MGPIO11B_F2H_GPIN => 
        VCC_net_1, MGPIO12A_F2H_GPIN => VCC_net_1, 
        MGPIO13A_F2H_GPIN => VCC_net_1, MGPIO14A_F2H_GPIN => 
        VCC_net_1, MGPIO15A_F2H_GPIN => VCC_net_1, 
        MGPIO16A_F2H_GPIN => VCC_net_1, MGPIO17B_F2H_GPIN => 
        VCC_net_1, MGPIO18B_F2H_GPIN => VCC_net_1, 
        MGPIO19B_F2H_GPIN => VCC_net_1, MGPIO1A_F2H_GPIN => 
        VCC_net_1, MGPIO20B_F2H_GPIN => VCC_net_1, 
        MGPIO21B_F2H_GPIN => VCC_net_1, MGPIO22B_F2H_GPIN => 
        VCC_net_1, MGPIO24B_F2H_GPIN => VCC_net_1, 
        MGPIO25B_F2H_GPIN => VCC_net_1, MGPIO26B_F2H_GPIN => 
        VCC_net_1, MGPIO27B_F2H_GPIN => VCC_net_1, 
        MGPIO28B_F2H_GPIN => VCC_net_1, MGPIO29B_F2H_GPIN => 
        VCC_net_1, MGPIO2A_F2H_GPIN => VCC_net_1, 
        MGPIO30B_F2H_GPIN => VCC_net_1, MGPIO31B_F2H_GPIN => 
        VCC_net_1, MGPIO3A_F2H_GPIN => VCC_net_1, 
        MGPIO4A_F2H_GPIN => VCC_net_1, MGPIO5A_F2H_GPIN => 
        VCC_net_1, MGPIO6A_F2H_GPIN => VCC_net_1, 
        MGPIO7A_F2H_GPIN => VCC_net_1, MGPIO8A_F2H_GPIN => 
        VCC_net_1, MGPIO9A_F2H_GPIN => VCC_net_1, 
        MMUART0_CTS_F2H_SCP => VCC_net_1, MMUART0_DCD_F2H_SCP => 
        VCC_net_1, MMUART0_DSR_F2H_SCP => VCC_net_1, 
        MMUART0_DTR_F2H_SCP => VCC_net_1, MMUART0_RI_F2H_SCP => 
        VCC_net_1, MMUART0_RTS_F2H_SCP => VCC_net_1, 
        MMUART0_RXD_F2H_SCP => VCC_net_1, MMUART0_SCK_F2H_SCP => 
        VCC_net_1, MMUART0_TXD_F2H_SCP => VCC_net_1, 
        MMUART1_CTS_F2H_SCP => VCC_net_1, MMUART1_DCD_F2H_SCP => 
        VCC_net_1, MMUART1_DSR_F2H_SCP => VCC_net_1, 
        MMUART1_RI_F2H_SCP => VCC_net_1, MMUART1_RTS_F2H_SCP => 
        VCC_net_1, MMUART1_RXD_F2H_SCP => VCC_net_1, 
        MMUART1_SCK_F2H_SCP => VCC_net_1, MMUART1_TXD_F2H_SCP => 
        VCC_net_1, PER2_FABRIC_PRDATA(31) => GND_net_1, 
        PER2_FABRIC_PRDATA(30) => GND_net_1, 
        PER2_FABRIC_PRDATA(29) => GND_net_1, 
        PER2_FABRIC_PRDATA(28) => GND_net_1, 
        PER2_FABRIC_PRDATA(27) => GND_net_1, 
        PER2_FABRIC_PRDATA(26) => GND_net_1, 
        PER2_FABRIC_PRDATA(25) => GND_net_1, 
        PER2_FABRIC_PRDATA(24) => GND_net_1, 
        PER2_FABRIC_PRDATA(23) => GND_net_1, 
        PER2_FABRIC_PRDATA(22) => GND_net_1, 
        PER2_FABRIC_PRDATA(21) => GND_net_1, 
        PER2_FABRIC_PRDATA(20) => GND_net_1, 
        PER2_FABRIC_PRDATA(19) => GND_net_1, 
        PER2_FABRIC_PRDATA(18) => GND_net_1, 
        PER2_FABRIC_PRDATA(17) => GND_net_1, 
        PER2_FABRIC_PRDATA(16) => GND_net_1, 
        PER2_FABRIC_PRDATA(15) => GND_net_1, 
        PER2_FABRIC_PRDATA(14) => GND_net_1, 
        PER2_FABRIC_PRDATA(13) => GND_net_1, 
        PER2_FABRIC_PRDATA(12) => GND_net_1, 
        PER2_FABRIC_PRDATA(11) => GND_net_1, 
        PER2_FABRIC_PRDATA(10) => GND_net_1, 
        PER2_FABRIC_PRDATA(9) => GND_net_1, PER2_FABRIC_PRDATA(8)
         => GND_net_1, PER2_FABRIC_PRDATA(7) => GND_net_1, 
        PER2_FABRIC_PRDATA(6) => GND_net_1, PER2_FABRIC_PRDATA(5)
         => GND_net_1, PER2_FABRIC_PRDATA(4) => GND_net_1, 
        PER2_FABRIC_PRDATA(3) => GND_net_1, PER2_FABRIC_PRDATA(2)
         => GND_net_1, PER2_FABRIC_PRDATA(1) => GND_net_1, 
        PER2_FABRIC_PRDATA(0) => GND_net_1, PER2_FABRIC_PREADY
         => VCC_net_1, PER2_FABRIC_PSLVERR => GND_net_1, RCGF(9)
         => VCC_net_1, RCGF(8) => VCC_net_1, RCGF(7) => VCC_net_1, 
        RCGF(6) => VCC_net_1, RCGF(5) => VCC_net_1, RCGF(4) => 
        VCC_net_1, RCGF(3) => VCC_net_1, RCGF(2) => VCC_net_1, 
        RCGF(1) => VCC_net_1, RCGF(0) => VCC_net_1, RX_CLKPF => 
        VCC_net_1, RX_DVF => VCC_net_1, RX_ERRF => VCC_net_1, 
        RX_EV => VCC_net_1, RXDF(7) => VCC_net_1, RXDF(6) => 
        VCC_net_1, RXDF(5) => VCC_net_1, RXDF(4) => VCC_net_1, 
        RXDF(3) => VCC_net_1, RXDF(2) => VCC_net_1, RXDF(1) => 
        VCC_net_1, RXDF(0) => VCC_net_1, SLEEPHOLDREQ => 
        GND_net_1, SMBALERT_NI0 => VCC_net_1, SMBALERT_NI1 => 
        VCC_net_1, SMBSUS_NI0 => VCC_net_1, SMBSUS_NI1 => 
        VCC_net_1, SPI0_CLK_IN => VCC_net_1, SPI0_SDI_F2H_SCP => 
        VCC_net_1, SPI0_SDO_F2H_SCP => VCC_net_1, 
        SPI0_SS0_F2H_SCP => VCC_net_1, SPI0_SS1_F2H_SCP => 
        VCC_net_1, SPI0_SS2_F2H_SCP => VCC_net_1, 
        SPI0_SS3_F2H_SCP => VCC_net_1, SPI1_CLK_IN => VCC_net_1, 
        SPI1_SDI_F2H_SCP => VCC_net_1, SPI1_SDO_F2H_SCP => 
        VCC_net_1, SPI1_SS0_F2H_SCP => VCC_net_1, 
        SPI1_SS1_F2H_SCP => VCC_net_1, SPI1_SS2_F2H_SCP => 
        VCC_net_1, SPI1_SS3_F2H_SCP => VCC_net_1, TX_CLKPF => 
        VCC_net_1, USER_MSS_GPIO_RESET_N => VCC_net_1, 
        USER_MSS_RESET_N => VCC_net_1, XCLK_FAB => VCC_net_1, 
        CLK_BASE => FAB_CCC_GL0, CLK_MDDR_APB => VCC_net_1, 
        F_ARADDR_HADDR1(31) => VCC_net_1, F_ARADDR_HADDR1(30) => 
        VCC_net_1, F_ARADDR_HADDR1(29) => VCC_net_1, 
        F_ARADDR_HADDR1(28) => VCC_net_1, F_ARADDR_HADDR1(27) => 
        VCC_net_1, F_ARADDR_HADDR1(26) => VCC_net_1, 
        F_ARADDR_HADDR1(25) => VCC_net_1, F_ARADDR_HADDR1(24) => 
        VCC_net_1, F_ARADDR_HADDR1(23) => VCC_net_1, 
        F_ARADDR_HADDR1(22) => VCC_net_1, F_ARADDR_HADDR1(21) => 
        VCC_net_1, F_ARADDR_HADDR1(20) => VCC_net_1, 
        F_ARADDR_HADDR1(19) => VCC_net_1, F_ARADDR_HADDR1(18) => 
        VCC_net_1, F_ARADDR_HADDR1(17) => VCC_net_1, 
        F_ARADDR_HADDR1(16) => VCC_net_1, F_ARADDR_HADDR1(15) => 
        VCC_net_1, F_ARADDR_HADDR1(14) => VCC_net_1, 
        F_ARADDR_HADDR1(13) => VCC_net_1, F_ARADDR_HADDR1(12) => 
        VCC_net_1, F_ARADDR_HADDR1(11) => VCC_net_1, 
        F_ARADDR_HADDR1(10) => VCC_net_1, F_ARADDR_HADDR1(9) => 
        VCC_net_1, F_ARADDR_HADDR1(8) => VCC_net_1, 
        F_ARADDR_HADDR1(7) => VCC_net_1, F_ARADDR_HADDR1(6) => 
        VCC_net_1, F_ARADDR_HADDR1(5) => VCC_net_1, 
        F_ARADDR_HADDR1(4) => VCC_net_1, F_ARADDR_HADDR1(3) => 
        VCC_net_1, F_ARADDR_HADDR1(2) => VCC_net_1, 
        F_ARADDR_HADDR1(1) => VCC_net_1, F_ARADDR_HADDR1(0) => 
        VCC_net_1, F_ARBURST_HTRANS1(1) => GND_net_1, 
        F_ARBURST_HTRANS1(0) => GND_net_1, F_ARID_HSEL1(3) => 
        GND_net_1, F_ARID_HSEL1(2) => GND_net_1, F_ARID_HSEL1(1)
         => GND_net_1, F_ARID_HSEL1(0) => GND_net_1, 
        F_ARLEN_HBURST1(3) => GND_net_1, F_ARLEN_HBURST1(2) => 
        GND_net_1, F_ARLEN_HBURST1(1) => GND_net_1, 
        F_ARLEN_HBURST1(0) => GND_net_1, F_ARLOCK_HMASTLOCK1(1)
         => GND_net_1, F_ARLOCK_HMASTLOCK1(0) => GND_net_1, 
        F_ARSIZE_HSIZE1(1) => GND_net_1, F_ARSIZE_HSIZE1(0) => 
        GND_net_1, F_ARVALID_HWRITE1 => GND_net_1, 
        F_AWADDR_HADDR0(31) => VCC_net_1, F_AWADDR_HADDR0(30) => 
        VCC_net_1, F_AWADDR_HADDR0(29) => VCC_net_1, 
        F_AWADDR_HADDR0(28) => VCC_net_1, F_AWADDR_HADDR0(27) => 
        VCC_net_1, F_AWADDR_HADDR0(26) => VCC_net_1, 
        F_AWADDR_HADDR0(25) => VCC_net_1, F_AWADDR_HADDR0(24) => 
        VCC_net_1, F_AWADDR_HADDR0(23) => VCC_net_1, 
        F_AWADDR_HADDR0(22) => VCC_net_1, F_AWADDR_HADDR0(21) => 
        VCC_net_1, F_AWADDR_HADDR0(20) => VCC_net_1, 
        F_AWADDR_HADDR0(19) => VCC_net_1, F_AWADDR_HADDR0(18) => 
        VCC_net_1, F_AWADDR_HADDR0(17) => VCC_net_1, 
        F_AWADDR_HADDR0(16) => VCC_net_1, F_AWADDR_HADDR0(15) => 
        VCC_net_1, F_AWADDR_HADDR0(14) => VCC_net_1, 
        F_AWADDR_HADDR0(13) => VCC_net_1, F_AWADDR_HADDR0(12) => 
        VCC_net_1, F_AWADDR_HADDR0(11) => VCC_net_1, 
        F_AWADDR_HADDR0(10) => VCC_net_1, F_AWADDR_HADDR0(9) => 
        VCC_net_1, F_AWADDR_HADDR0(8) => VCC_net_1, 
        F_AWADDR_HADDR0(7) => VCC_net_1, F_AWADDR_HADDR0(6) => 
        VCC_net_1, F_AWADDR_HADDR0(5) => VCC_net_1, 
        F_AWADDR_HADDR0(4) => VCC_net_1, F_AWADDR_HADDR0(3) => 
        VCC_net_1, F_AWADDR_HADDR0(2) => VCC_net_1, 
        F_AWADDR_HADDR0(1) => VCC_net_1, F_AWADDR_HADDR0(0) => 
        VCC_net_1, F_AWBURST_HTRANS0(1) => GND_net_1, 
        F_AWBURST_HTRANS0(0) => GND_net_1, F_AWID_HSEL0(3) => 
        GND_net_1, F_AWID_HSEL0(2) => GND_net_1, F_AWID_HSEL0(1)
         => GND_net_1, F_AWID_HSEL0(0) => GND_net_1, 
        F_AWLEN_HBURST0(3) => GND_net_1, F_AWLEN_HBURST0(2) => 
        GND_net_1, F_AWLEN_HBURST0(1) => GND_net_1, 
        F_AWLEN_HBURST0(0) => GND_net_1, F_AWLOCK_HMASTLOCK0(1)
         => GND_net_1, F_AWLOCK_HMASTLOCK0(0) => GND_net_1, 
        F_AWSIZE_HSIZE0(1) => GND_net_1, F_AWSIZE_HSIZE0(0) => 
        GND_net_1, F_AWVALID_HWRITE0 => GND_net_1, F_BREADY => 
        GND_net_1, F_RMW_AXI => GND_net_1, F_RREADY => GND_net_1, 
        F_WDATA_HWDATA01(63) => VCC_net_1, F_WDATA_HWDATA01(62)
         => VCC_net_1, F_WDATA_HWDATA01(61) => VCC_net_1, 
        F_WDATA_HWDATA01(60) => VCC_net_1, F_WDATA_HWDATA01(59)
         => VCC_net_1, F_WDATA_HWDATA01(58) => VCC_net_1, 
        F_WDATA_HWDATA01(57) => VCC_net_1, F_WDATA_HWDATA01(56)
         => VCC_net_1, F_WDATA_HWDATA01(55) => VCC_net_1, 
        F_WDATA_HWDATA01(54) => VCC_net_1, F_WDATA_HWDATA01(53)
         => VCC_net_1, F_WDATA_HWDATA01(52) => VCC_net_1, 
        F_WDATA_HWDATA01(51) => VCC_net_1, F_WDATA_HWDATA01(50)
         => VCC_net_1, F_WDATA_HWDATA01(49) => VCC_net_1, 
        F_WDATA_HWDATA01(48) => VCC_net_1, F_WDATA_HWDATA01(47)
         => VCC_net_1, F_WDATA_HWDATA01(46) => VCC_net_1, 
        F_WDATA_HWDATA01(45) => VCC_net_1, F_WDATA_HWDATA01(44)
         => VCC_net_1, F_WDATA_HWDATA01(43) => VCC_net_1, 
        F_WDATA_HWDATA01(42) => VCC_net_1, F_WDATA_HWDATA01(41)
         => VCC_net_1, F_WDATA_HWDATA01(40) => VCC_net_1, 
        F_WDATA_HWDATA01(39) => VCC_net_1, F_WDATA_HWDATA01(38)
         => VCC_net_1, F_WDATA_HWDATA01(37) => VCC_net_1, 
        F_WDATA_HWDATA01(36) => VCC_net_1, F_WDATA_HWDATA01(35)
         => VCC_net_1, F_WDATA_HWDATA01(34) => VCC_net_1, 
        F_WDATA_HWDATA01(33) => VCC_net_1, F_WDATA_HWDATA01(32)
         => VCC_net_1, F_WDATA_HWDATA01(31) => VCC_net_1, 
        F_WDATA_HWDATA01(30) => VCC_net_1, F_WDATA_HWDATA01(29)
         => VCC_net_1, F_WDATA_HWDATA01(28) => VCC_net_1, 
        F_WDATA_HWDATA01(27) => VCC_net_1, F_WDATA_HWDATA01(26)
         => VCC_net_1, F_WDATA_HWDATA01(25) => VCC_net_1, 
        F_WDATA_HWDATA01(24) => VCC_net_1, F_WDATA_HWDATA01(23)
         => VCC_net_1, F_WDATA_HWDATA01(22) => VCC_net_1, 
        F_WDATA_HWDATA01(21) => VCC_net_1, F_WDATA_HWDATA01(20)
         => VCC_net_1, F_WDATA_HWDATA01(19) => VCC_net_1, 
        F_WDATA_HWDATA01(18) => VCC_net_1, F_WDATA_HWDATA01(17)
         => VCC_net_1, F_WDATA_HWDATA01(16) => VCC_net_1, 
        F_WDATA_HWDATA01(15) => VCC_net_1, F_WDATA_HWDATA01(14)
         => VCC_net_1, F_WDATA_HWDATA01(13) => VCC_net_1, 
        F_WDATA_HWDATA01(12) => VCC_net_1, F_WDATA_HWDATA01(11)
         => VCC_net_1, F_WDATA_HWDATA01(10) => VCC_net_1, 
        F_WDATA_HWDATA01(9) => VCC_net_1, F_WDATA_HWDATA01(8) => 
        VCC_net_1, F_WDATA_HWDATA01(7) => VCC_net_1, 
        F_WDATA_HWDATA01(6) => VCC_net_1, F_WDATA_HWDATA01(5) => 
        VCC_net_1, F_WDATA_HWDATA01(4) => VCC_net_1, 
        F_WDATA_HWDATA01(3) => VCC_net_1, F_WDATA_HWDATA01(2) => 
        VCC_net_1, F_WDATA_HWDATA01(1) => VCC_net_1, 
        F_WDATA_HWDATA01(0) => VCC_net_1, F_WID_HREADY01(3) => 
        GND_net_1, F_WID_HREADY01(2) => GND_net_1, 
        F_WID_HREADY01(1) => GND_net_1, F_WID_HREADY01(0) => 
        GND_net_1, F_WLAST => GND_net_1, F_WSTRB(7) => GND_net_1, 
        F_WSTRB(6) => GND_net_1, F_WSTRB(5) => GND_net_1, 
        F_WSTRB(4) => GND_net_1, F_WSTRB(3) => GND_net_1, 
        F_WSTRB(2) => GND_net_1, F_WSTRB(1) => GND_net_1, 
        F_WSTRB(0) => GND_net_1, F_WVALID => GND_net_1, 
        FPGA_MDDR_ARESET_N => VCC_net_1, MDDR_FABRIC_PADDR(10)
         => VCC_net_1, MDDR_FABRIC_PADDR(9) => VCC_net_1, 
        MDDR_FABRIC_PADDR(8) => VCC_net_1, MDDR_FABRIC_PADDR(7)
         => VCC_net_1, MDDR_FABRIC_PADDR(6) => VCC_net_1, 
        MDDR_FABRIC_PADDR(5) => VCC_net_1, MDDR_FABRIC_PADDR(4)
         => VCC_net_1, MDDR_FABRIC_PADDR(3) => VCC_net_1, 
        MDDR_FABRIC_PADDR(2) => VCC_net_1, MDDR_FABRIC_PENABLE
         => VCC_net_1, MDDR_FABRIC_PSEL => VCC_net_1, 
        MDDR_FABRIC_PWDATA(15) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(14) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(13) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(12) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(11) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(10) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(9) => VCC_net_1, MDDR_FABRIC_PWDATA(8)
         => VCC_net_1, MDDR_FABRIC_PWDATA(7) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(6) => VCC_net_1, MDDR_FABRIC_PWDATA(5)
         => VCC_net_1, MDDR_FABRIC_PWDATA(4) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(3) => VCC_net_1, MDDR_FABRIC_PWDATA(2)
         => VCC_net_1, MDDR_FABRIC_PWDATA(1) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(0) => VCC_net_1, MDDR_FABRIC_PWRITE
         => VCC_net_1, PRESET_N => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => GND_net_1, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => GND_net_1, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => GND_net_1, DM_IN(2)
         => GND_net_1, DM_IN(1) => GND_net_1, DM_IN(0) => 
        GND_net_1, DRAM_DQ_IN(17) => GND_net_1, DRAM_DQ_IN(16)
         => GND_net_1, DRAM_DQ_IN(15) => GND_net_1, 
        DRAM_DQ_IN(14) => GND_net_1, DRAM_DQ_IN(13) => GND_net_1, 
        DRAM_DQ_IN(12) => GND_net_1, DRAM_DQ_IN(11) => GND_net_1, 
        DRAM_DQ_IN(10) => GND_net_1, DRAM_DQ_IN(9) => GND_net_1, 
        DRAM_DQ_IN(8) => GND_net_1, DRAM_DQ_IN(7) => GND_net_1, 
        DRAM_DQ_IN(6) => GND_net_1, DRAM_DQ_IN(5) => GND_net_1, 
        DRAM_DQ_IN(4) => GND_net_1, DRAM_DQ_IN(3) => GND_net_1, 
        DRAM_DQ_IN(2) => GND_net_1, DRAM_DQ_IN(1) => GND_net_1, 
        DRAM_DQ_IN(0) => GND_net_1, DRAM_DQS_IN(2) => GND_net_1, 
        DRAM_DQS_IN(1) => GND_net_1, DRAM_DQS_IN(0) => GND_net_1, 
        DRAM_FIFO_WE_IN(1) => GND_net_1, DRAM_FIFO_WE_IN(0) => 
        GND_net_1, I2C0_SCL_USBC_DATA1_MGPIO31B_IN => GND_net_1, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => GND_net_1, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => GND_net_1, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => GND_net_1, MGPIO0B_IN
         => GND_net_1, MGPIO10B_IN => GND_net_1, MGPIO1B_IN => 
        GND_net_1, MGPIO25A_IN => GND_net_1, MGPIO26A_IN => 
        GND_net_1, MGPIO27A_IN => GND_net_1, MGPIO28A_IN => 
        GND_net_1, MGPIO29A_IN => GND_net_1, MGPIO2B_IN => 
        GND_net_1, MGPIO30A_IN => GND_net_1, MGPIO31A_IN => 
        GND_net_1, MGPIO3B_IN => GND_net_1, MGPIO4B_IN => 
        GND_net_1, MGPIO5B_IN => GND_net_1, MGPIO6B_IN => 
        GND_net_1, MGPIO7B_IN => GND_net_1, MGPIO8B_IN => 
        GND_net_1, MGPIO9B_IN => GND_net_1, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => GND_net_1, 
        MMUART0_DCD_MGPIO22B_IN => GND_net_1, 
        MMUART0_DSR_MGPIO20B_IN => GND_net_1, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => GND_net_1, 
        MMUART0_RI_MGPIO21B_IN => GND_net_1, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => GND_net_1, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => GND_net_1, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => GND_net_1, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => GND_net_1, 
        MMUART1_CTS_MGPIO13B_IN => GND_net_1, 
        MMUART1_DCD_MGPIO16B_IN => GND_net_1, 
        MMUART1_DSR_MGPIO14B_IN => GND_net_1, 
        MMUART1_DTR_MGPIO12B_IN => GND_net_1, 
        MMUART1_RI_MGPIO15B_IN => GND_net_1, 
        MMUART1_RTS_MGPIO11B_IN => GND_net_1, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => MMUART_1_RXD_PAD_Y, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => GND_net_1, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => GND_net_1, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => GND_net_1, 
        RGMII_MDC_RMII_MDC_IN => GND_net_1, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => GND_net_1, 
        RGMII_RX_CLK_IN => GND_net_1, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => GND_net_1, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => GND_net_1, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => GND_net_1, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => GND_net_1, 
        RGMII_RXD3_USBB_DATA4_IN => GND_net_1, RGMII_TX_CLK_IN
         => GND_net_1, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => 
        GND_net_1, RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => GND_net_1, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => GND_net_1, 
        RGMII_TXD2_USBB_DATA5_IN => GND_net_1, 
        RGMII_TXD3_USBB_DATA6_IN => GND_net_1, 
        SPI0_SCK_USBA_XCLK_IN => SPI_0_CLK_PAD_Y, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => SPI_0_DI_PAD_Y, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => GND_net_1, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => SPI_0_SS0_PAD_Y, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => GND_net_1, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => GND_net_1, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => GND_net_1, 
        SPI0_SS4_MGPIO19A_IN => GND_net_1, SPI0_SS5_MGPIO20A_IN
         => GND_net_1, SPI0_SS6_MGPIO21A_IN => GND_net_1, 
        SPI0_SS7_MGPIO22A_IN => GND_net_1, SPI1_SCK_IN => 
        GND_net_1, SPI1_SDI_MGPIO11A_IN => GND_net_1, 
        SPI1_SDO_MGPIO12A_IN => GND_net_1, SPI1_SS0_MGPIO13A_IN
         => GND_net_1, SPI1_SS1_MGPIO14A_IN => GND_net_1, 
        SPI1_SS2_MGPIO15A_IN => GND_net_1, SPI1_SS3_MGPIO16A_IN
         => GND_net_1, SPI1_SS4_MGPIO17A_IN => GND_net_1, 
        SPI1_SS5_MGPIO18A_IN => GND_net_1, SPI1_SS6_MGPIO23A_IN
         => GND_net_1, SPI1_SS7_MGPIO24A_IN => GND_net_1, 
        USBC_XCLK_IN => GND_net_1, USBD_DATA0_IN => GND_net_1, 
        USBD_DATA1_IN => GND_net_1, USBD_DATA2_IN => GND_net_1, 
        USBD_DATA3_IN => GND_net_1, USBD_DATA4_IN => GND_net_1, 
        USBD_DATA5_IN => GND_net_1, USBD_DATA6_IN => GND_net_1, 
        USBD_DATA7_MGPIO23B_IN => GND_net_1, USBD_DIR_IN => 
        GND_net_1, USBD_NXT_IN => GND_net_1, USBD_STP_IN => 
        GND_net_1, USBD_XCLK_IN => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => OPEN, DRAM_ADDR(15)
         => nc21, DRAM_ADDR(14) => nc237, DRAM_ADDR(13) => nc93, 
        DRAM_ADDR(12) => nc262, DRAM_ADDR(11) => nc69, 
        DRAM_ADDR(10) => nc206, DRAM_ADDR(9) => nc174, 
        DRAM_ADDR(8) => nc38, DRAM_ADDR(7) => nc113, DRAM_ADDR(6)
         => nc218, DRAM_ADDR(5) => nc106, DRAM_ADDR(4) => nc261, 
        DRAM_ADDR(3) => nc25, DRAM_ADDR(2) => nc1, DRAM_ADDR(1)
         => nc299, DRAM_ADDR(0) => nc37, DRAM_BA(2) => nc202, 
        DRAM_BA(1) => nc144, DRAM_BA(0) => nc153, DRAM_CASN => 
        OPEN, DRAM_CKE => OPEN, DRAM_CLK => OPEN, DRAM_CSN => 
        OPEN, DRAM_DM_RDQS_OUT(2) => nc46, DRAM_DM_RDQS_OUT(1)
         => nc258, DRAM_DM_RDQS_OUT(0) => nc71, DRAM_DQ_OUT(17)
         => nc124, DRAM_DQ_OUT(16) => nc81, DRAM_DQ_OUT(15) => 
        nc201, DRAM_DQ_OUT(14) => nc168, DRAM_DQ_OUT(13) => nc34, 
        DRAM_DQ_OUT(12) => nc28, DRAM_DQ_OUT(11) => nc115, 
        DRAM_DQ_OUT(10) => nc264, DRAM_DQ_OUT(9) => nc192, 
        DRAM_DQ_OUT(8) => nc319, DRAM_DQ_OUT(7) => nc134, 
        DRAM_DQ_OUT(6) => nc32, DRAM_DQ_OUT(5) => nc40, 
        DRAM_DQ_OUT(4) => nc297, DRAM_DQ_OUT(3) => nc99, 
        DRAM_DQ_OUT(2) => nc75, DRAM_DQ_OUT(1) => nc183, 
        DRAM_DQ_OUT(0) => nc288, DRAM_DQS_OUT(2) => nc85, 
        DRAM_DQS_OUT(1) => nc27, DRAM_DQS_OUT(0) => nc108, 
        DRAM_FIFO_WE_OUT(1) => nc16, DRAM_FIFO_WE_OUT(0) => nc155, 
        DRAM_ODT => OPEN, DRAM_RASN => OPEN, DRAM_RSTN => OPEN, 
        DRAM_WEN => OPEN, I2C0_SCL_USBC_DATA1_MGPIO31B_OUT => 
        OPEN, I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => OPEN, MGPIO0B_OUT => 
        OPEN, MGPIO10B_OUT => OPEN, MGPIO1B_OUT => OPEN, 
        MGPIO25A_OUT => OPEN, MGPIO26A_OUT => OPEN, MGPIO27A_OUT
         => OPEN, MGPIO28A_OUT => OPEN, MGPIO29A_OUT => OPEN, 
        MGPIO2B_OUT => OPEN, MGPIO30A_OUT => OPEN, MGPIO31A_OUT
         => OPEN, MGPIO3B_OUT => OPEN, MGPIO4B_OUT => OPEN, 
        MGPIO5B_OUT => OPEN, MGPIO6B_OUT => OPEN, MGPIO7B_OUT => 
        OPEN, MGPIO8B_OUT => OPEN, MGPIO9B_OUT => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT => OPEN, 
        MMUART0_DCD_MGPIO22B_OUT => OPEN, 
        MMUART0_DSR_MGPIO20B_OUT => OPEN, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => OPEN, 
        MMUART1_CTS_MGPIO13B_OUT => OPEN, 
        MMUART1_DCD_MGPIO16B_OUT => OPEN, 
        MMUART1_DSR_MGPIO14B_OUT => OPEN, 
        MMUART1_DTR_MGPIO12B_OUT => OPEN, MMUART1_RI_MGPIO15B_OUT
         => OPEN, MMUART1_RTS_MGPIO11B_OUT => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => OPEN, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => OPEN, 
        RGMII_RXD3_USBB_DATA4_OUT => OPEN, RGMII_TX_CLK_OUT => 
        OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => OPEN, 
        RGMII_TXD2_USBB_DATA5_OUT => OPEN, 
        RGMII_TXD3_USBB_DATA6_OUT => OPEN, SPI0_SCK_USBA_XCLK_OUT
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => OPEN, 
        SPI0_SS4_MGPIO19A_OUT => OPEN, SPI0_SS5_MGPIO20A_OUT => 
        OPEN, SPI0_SS6_MGPIO21A_OUT => OPEN, 
        SPI0_SS7_MGPIO22A_OUT => OPEN, SPI1_SCK_OUT => OPEN, 
        SPI1_SDI_MGPIO11A_OUT => OPEN, SPI1_SDO_MGPIO12A_OUT => 
        OPEN, SPI1_SS0_MGPIO13A_OUT => OPEN, 
        SPI1_SS1_MGPIO14A_OUT => OPEN, SPI1_SS2_MGPIO15A_OUT => 
        OPEN, SPI1_SS3_MGPIO16A_OUT => OPEN, 
        SPI1_SS4_MGPIO17A_OUT => OPEN, SPI1_SS5_MGPIO18A_OUT => 
        OPEN, SPI1_SS6_MGPIO23A_OUT => OPEN, 
        SPI1_SS7_MGPIO24A_OUT => OPEN, USBC_XCLK_OUT => OPEN, 
        USBD_DATA0_OUT => OPEN, USBD_DATA1_OUT => OPEN, 
        USBD_DATA2_OUT => OPEN, USBD_DATA3_OUT => OPEN, 
        USBD_DATA4_OUT => OPEN, USBD_DATA5_OUT => OPEN, 
        USBD_DATA6_OUT => OPEN, USBD_DATA7_MGPIO23B_OUT => OPEN, 
        USBD_DIR_OUT => OPEN, USBD_NXT_OUT => OPEN, USBD_STP_OUT
         => OPEN, USBD_XCLK_OUT => OPEN, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => OPEN, DM_OE(2) => nc51, 
        DM_OE(1) => nc301, DM_OE(0) => nc33, DRAM_DQ_OE(17) => 
        nc204, DRAM_DQ_OE(16) => nc173, DRAM_DQ_OE(15) => nc278, 
        DRAM_DQ_OE(14) => nc169, DRAM_DQ_OE(13) => nc78, 
        DRAM_DQ_OE(12) => nc263, DRAM_DQ_OE(11) => nc24, 
        DRAM_DQ_OE(10) => nc88, DRAM_DQ_OE(9) => nc111, 
        DRAM_DQ_OE(8) => nc55, DRAM_DQ_OE(7) => nc10, 
        DRAM_DQ_OE(6) => nc22, DRAM_DQ_OE(5) => nc210, 
        DRAM_DQ_OE(4) => nc185, DRAM_DQ_OE(3) => nc143, 
        DRAM_DQ_OE(2) => nc248, DRAM_DQ_OE(1) => nc77, 
        DRAM_DQ_OE(0) => nc6, DRAM_DQS_OE(2) => nc109, 
        DRAM_DQS_OE(1) => nc87, DRAM_DQS_OE(0) => nc123, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => OPEN, MGPIO0B_OE => 
        OPEN, MGPIO10B_OE => OPEN, MGPIO1B_OE => OPEN, 
        MGPIO25A_OE => OPEN, MGPIO26A_OE => OPEN, MGPIO27A_OE => 
        OPEN, MGPIO28A_OE => OPEN, MGPIO29A_OE => OPEN, 
        MGPIO2B_OE => OPEN, MGPIO30A_OE => OPEN, MGPIO31A_OE => 
        OPEN, MGPIO3B_OE => OPEN, MGPIO4B_OE => OPEN, MGPIO5B_OE
         => OPEN, MGPIO6B_OE => OPEN, MGPIO7B_OE => OPEN, 
        MGPIO8B_OE => OPEN, MGPIO9B_OE => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => OPEN, 
        MMUART0_DCD_MGPIO22B_OE => OPEN, MMUART0_DSR_MGPIO20B_OE
         => OPEN, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => OPEN, 
        MMUART1_CTS_MGPIO13B_OE => OPEN, MMUART1_DCD_MGPIO16B_OE
         => OPEN, MMUART1_DSR_MGPIO14B_OE => OPEN, 
        MMUART1_DTR_MGPIO12B_OE => OPEN, MMUART1_RI_MGPIO15B_OE
         => OPEN, MMUART1_RTS_MGPIO11B_OE => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => OPEN, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => OPEN, 
        RGMII_RXD3_USBB_DATA4_OE => OPEN, RGMII_TX_CLK_OE => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => OPEN, 
        RGMII_TXD2_USBB_DATA5_OE => OPEN, 
        RGMII_TXD3_USBB_DATA6_OE => OPEN, SPI0_SCK_USBA_XCLK_OE
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => OPEN, 
        SPI0_SS4_MGPIO19A_OE => OPEN, SPI0_SS5_MGPIO20A_OE => 
        OPEN, SPI0_SS6_MGPIO21A_OE => OPEN, SPI0_SS7_MGPIO22A_OE
         => OPEN, SPI1_SCK_OE => OPEN, SPI1_SDI_MGPIO11A_OE => 
        OPEN, SPI1_SDO_MGPIO12A_OE => OPEN, SPI1_SS0_MGPIO13A_OE
         => OPEN, SPI1_SS1_MGPIO14A_OE => OPEN, 
        SPI1_SS2_MGPIO15A_OE => OPEN, SPI1_SS3_MGPIO16A_OE => 
        OPEN, SPI1_SS4_MGPIO17A_OE => OPEN, SPI1_SS5_MGPIO18A_OE
         => OPEN, SPI1_SS6_MGPIO23A_OE => OPEN, 
        SPI1_SS7_MGPIO24A_OE => OPEN, USBC_XCLK_OE => OPEN, 
        USBD_DATA0_OE => OPEN, USBD_DATA1_OE => OPEN, 
        USBD_DATA2_OE => OPEN, USBD_DATA3_OE => OPEN, 
        USBD_DATA4_OE => OPEN, USBD_DATA5_OE => OPEN, 
        USBD_DATA6_OE => OPEN, USBD_DATA7_MGPIO23B_OE => OPEN, 
        USBD_DIR_OE => OPEN, USBD_NXT_OE => OPEN, USBD_STP_OE => 
        OPEN, USBD_XCLK_OE => OPEN);
    
    MSS_ADLIB_INST_RNO_5 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(6), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[6]\);
    
    SPI_0_CLK_PAD : BIBUF
      port map(PAD => SPI_0_CLK, D => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, E => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, Y => 
        SPI_0_CLK_PAD_Y);
    
    MSS_ADLIB_INST_RNO_25 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(26), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[26]\);
    
    MSS_ADLIB_INST_RNO_24 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(25), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[25]\);
    
    MSS_ADLIB_INST_RNO_1 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(2), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[2]\);
    
    MSS_ADLIB_INST_RNO_30 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(31), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[31]\);
    
    MSS_ADLIB_INST_RNO_26 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(27), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[27]\);
    
    SPI_0_SS0_PAD : BIBUF
      port map(PAD => SPI_0_SS0, D => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, Y => 
        SPI_0_SS0_PAD_Y);
    
    MSS_ADLIB_INST_RNO_8 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(9), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[9]\);
    
    MSS_ADLIB_INST_RNO_6 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(7), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[7]\);
    
    MSS_ADLIB_INST_RNO_28 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(29), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[29]\);
    
    MSS_ADLIB_INST_RNO_9 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(10), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[10]\);
    
    MSS_ADLIB_INST_RNO_15 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(16), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[16]\);
    
    MSS_ADLIB_INST_RNO_0 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(1), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[1]\);
    
    MSS_ADLIB_INST_RNO_14 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(15), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[15]\);
    
    MMUART_1_RXD_PAD : INBUF
      port map(PAD => MMUART_1_RXD, Y => MMUART_1_RXD_PAD_Y);
    
    MSS_ADLIB_INST_RNO_16 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(17), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[17]\);
    
    MSS_ADLIB_INST_RNO_18 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(19), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[19]\);
    
    MSS_ADLIB_INST_RNO_3 : CFG2
      generic map(INIT => x"8")

      port map(A => xhdl1250_i_m_1(0), B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(4), Y => 
        \CoreAHBLite_0_AHBmslave3_HRDATA_m[4]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_CCC_0_FCCC is

    port( FAB_CCC_GL0                                        : out   std_logic;
          FAB_CCC_LOCK                                       : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic
        );

end CertificationSystem_sb_CCC_0_FCCC;

architecture DEF_ARCH of CertificationSystem_sb_CCC_0_FCCC is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => FAB_CCC_GL0);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007FB8000045174000318C6318C1F18C61EC0404040400101",
         VCOFREQUENCY => 800.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => FAB_CCC_LOCK, 
        BUSY => OPEN, CLK0 => VCC_net_1, CLK1 => VCC_net_1, CLK2
         => VCC_net_1, CLK3 => VCC_net_1, NGMUX0_SEL => GND_net_1, 
        NGMUX1_SEL => GND_net_1, NGMUX2_SEL => GND_net_1, 
        NGMUX3_SEL => GND_net_1, NGMUX0_HOLD_N => VCC_net_1, 
        NGMUX1_HOLD_N => VCC_net_1, NGMUX2_HOLD_N => VCC_net_1, 
        NGMUX3_HOLD_N => VCC_net_1, NGMUX0_ARST_N => VCC_net_1, 
        NGMUX1_ARST_N => VCC_net_1, NGMUX2_ARST_N => VCC_net_1, 
        NGMUX3_ARST_N => VCC_net_1, PLL_BYPASS_N => VCC_net_1, 
        PLL_ARST_N => VCC_net_1, PLL_POWERDOWN_N => VCC_net_1, 
        GPD0_ARST_N => VCC_net_1, GPD1_ARST_N => VCC_net_1, 
        GPD2_ARST_N => VCC_net_1, GPD3_ARST_N => VCC_net_1, 
        PRESET_N => GND_net_1, PCLK => VCC_net_1, PSEL => 
        VCC_net_1, PENABLE => VCC_net_1, PWRITE => VCC_net_1, 
        PADDR(7) => VCC_net_1, PADDR(6) => VCC_net_1, PADDR(5)
         => VCC_net_1, PADDR(4) => VCC_net_1, PADDR(3) => 
        VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7) => VCC_net_1, 
        PWDATA(6) => VCC_net_1, PWDATA(5) => VCC_net_1, PWDATA(4)
         => VCC_net_1, PWDATA(3) => VCC_net_1, PWDATA(2) => 
        VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0) => VCC_net_1, 
        CLK0_PAD => GND_net_1, CLK1_PAD => GND_net_1, CLK2_PAD
         => GND_net_1, CLK3_PAD => GND_net_1, GL0 => GL0_net, GL1
         => OPEN, GL2 => OPEN, GL3 => OPEN, RCOSC_25_50MHZ => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        RCOSC_1MHZ => GND_net_1, XTLOSC => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity 
        CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8 is

    port( ram_rdata                       : out   std_logic_vector(31 downto 0);
          sram_wen_mem                    : in    std_logic_vector(3 downto 0);
          ahbsram_addr                    : in    std_logic_vector(15 downto 2);
          CoreAHBLite_0_AHBmslave3_HWDATA : in    std_logic_vector(31 downto 0);
          FAB_CCC_GL0                     : in    std_logic;
          MSS_READY                       : in    std_logic;
          N_21_i_0                        : in    std_logic
        );

end CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8;

architecture DEF_ARCH of 
        CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal readdata_xhdl1419_0_a2_0, \wen_b1_1[1]\, 
        \wen_b1_1[0]\, \readData_31_am_RNO[0]_net_1\, 
        \readData_31_am_1_1[0]_net_1\, 
        \readData_31_am_RNO_0[0]_net_1\, 
        \readData_31_am[0]_net_1\, 
        \readData_31_am_1_1_RNO[0]_net_1\, 
        \readData_31_am_1_1_RNO_0[0]_net_1\, 
        \readData_31_bm_RNO[0]_net_1\, 
        \readData_31_bm_1_1[0]_net_1\, 
        \readData_31_bm_RNO_0[0]_net_1\, 
        \readData_31_bm[0]_net_1\, 
        \readData_31_bm_1_1_RNO[0]_net_1\, 
        \readData_31_bm_1_1_RNO_0[0]_net_1\, 
        \readData_31_am_RNO[1]_net_1\, 
        \readData_31_am_1_1[1]_net_1\, 
        \readData_31_am_RNO_0[1]_net_1\, 
        \readData_31_am[1]_net_1\, 
        \readData_31_am_1_1_RNO[1]_net_1\, 
        \readData_31_am_1_1_RNO_0[1]_net_1\, 
        \readData_31_bm_RNO[1]_net_1\, 
        \readData_31_bm_1_1[1]_net_1\, 
        \readData_31_bm_RNO_0[1]_net_1\, 
        \readData_31_bm[1]_net_1\, 
        \readData_31_bm_1_1_RNO[1]_net_1\, 
        \readData_31_bm_1_1_RNO_0[1]_net_1\, 
        \readData_31_am_RNO[2]_net_1\, 
        \readData_31_am_1_1[2]_net_1\, 
        \readData_31_am_RNO_0[2]_net_1\, 
        \readData_31_am[2]_net_1\, 
        \readData_31_am_1_1_RNO[2]_net_1\, 
        \readData_31_am_1_1_RNO_0[2]_net_1\, 
        \readData_31_bm_RNO[2]_net_1\, 
        \readData_31_bm_1_1[2]_net_1\, 
        \readData_31_bm_RNO_0[2]_net_1\, 
        \readData_31_bm[2]_net_1\, 
        \readData_31_bm_1_1_RNO[2]_net_1\, 
        \readData_31_bm_1_1_RNO_0[2]_net_1\, 
        \readData_31_am_RNO[3]_net_1\, 
        \readData_31_am_1_1[3]_net_1\, 
        \readData_31_am_RNO_0[3]_net_1\, 
        \readData_31_am[3]_net_1\, 
        \readData_31_am_1_1_RNO[3]_net_1\, 
        \readData_31_am_1_1_RNO_0[3]_net_1\, 
        \readData_31_bm_RNO[3]_net_1\, 
        \readData_31_bm_1_1[3]_net_1\, 
        \readData_31_bm_RNO_0[3]_net_1\, 
        \readData_31_bm[3]_net_1\, 
        \readData_31_bm_1_1_RNO[3]_net_1\, 
        \readData_31_bm_1_1_RNO_0[3]_net_1\, 
        \readData_31_am_RNO[4]_net_1\, 
        \readData_31_am_1_1[4]_net_1\, 
        \readData_31_am_RNO_0[4]_net_1\, 
        \readData_31_am[4]_net_1\, 
        \readData_31_am_1_1_RNO[4]_net_1\, 
        \readData_31_am_1_1_RNO_0[4]_net_1\, 
        \readData_31_bm_RNO[4]_net_1\, 
        \readData_31_bm_1_1[4]_net_1\, 
        \readData_31_bm_RNO_0[4]_net_1\, 
        \readData_31_bm[4]_net_1\, 
        \readData_31_bm_1_1_RNO[4]_net_1\, 
        \readData_31_bm_1_1_RNO_0[4]_net_1\, 
        \readData_31_am_RNO[5]_net_1\, 
        \readData_31_am_1_1[5]_net_1\, 
        \readData_31_am_RNO_0[5]_net_1\, 
        \readData_31_am[5]_net_1\, 
        \readData_31_am_1_1_RNO[5]_net_1\, 
        \readData_31_am_1_1_RNO_0[5]_net_1\, 
        \readData_31_bm_RNO[5]_net_1\, 
        \readData_31_bm_1_1[5]_net_1\, 
        \readData_31_bm_RNO_0[5]_net_1\, 
        \readData_31_bm[5]_net_1\, 
        \readData_31_bm_1_1_RNO[5]_net_1\, 
        \readData_31_bm_1_1_RNO_0[5]_net_1\, 
        \readData_31_am_RNO[6]_net_1\, 
        \readData_31_am_1_1[6]_net_1\, 
        \readData_31_am_RNO_0[6]_net_1\, 
        \readData_31_am[6]_net_1\, 
        \readData_31_am_1_1_RNO[6]_net_1\, 
        \readData_31_am_1_1_RNO_0[6]_net_1\, 
        \readData_31_bm_RNO[6]_net_1\, 
        \readData_31_bm_1_1[6]_net_1\, 
        \readData_31_bm_RNO_0[6]_net_1\, 
        \readData_31_bm[6]_net_1\, 
        \readData_31_bm_1_1_RNO[6]_net_1\, 
        \readData_31_bm_1_1_RNO_0[6]_net_1\, 
        \readData_31_am_RNO[7]_net_1\, 
        \readData_31_am_1_1[7]_net_1\, 
        \readData_31_am_RNO_0[7]_net_1\, 
        \readData_31_am[7]_net_1\, 
        \readData_31_am_1_1_RNO[7]_net_1\, 
        \readData_31_am_1_1_RNO_0[7]_net_1\, 
        \readData_31_bm_RNO[7]_net_1\, 
        \readData_31_bm_1_1[7]_net_1\, 
        \readData_31_bm_RNO_0[7]_net_1\, 
        \readData_31_bm[7]_net_1\, 
        \readData_31_bm_1_1_RNO[7]_net_1\, 
        \readData_31_bm_1_1_RNO_0[7]_net_1\, 
        \readData_31_am_RNO[8]_net_1\, 
        \readData_31_am_1_1[8]_net_1\, 
        \readData_31_am_RNO_0[8]_net_1\, 
        \readData_31_am[8]_net_1\, 
        \readData_31_am_1_1_RNO[8]_net_1\, 
        \readData_31_am_1_1_RNO_0[8]_net_1\, 
        \readData_31_bm_RNO[8]_net_1\, 
        \readData_31_bm_1_1[8]_net_1\, 
        \readData_31_bm_RNO_0[8]_net_1\, 
        \readData_31_bm[8]_net_1\, 
        \readData_31_bm_1_1_RNO[8]_net_1\, 
        \readData_31_bm_1_1_RNO_0[8]_net_1\, 
        \readData_31_am_RNO[9]_net_1\, 
        \readData_31_am_1_1[9]_net_1\, 
        \readData_31_am_RNO_0[9]_net_1\, 
        \readData_31_am[9]_net_1\, 
        \readData_31_am_1_1_RNO[9]_net_1\, 
        \readData_31_am_1_1_RNO_0[9]_net_1\, 
        \readData_31_bm_RNO[9]_net_1\, 
        \readData_31_bm_1_1[9]_net_1\, 
        \readData_31_bm_RNO_0[9]_net_1\, 
        \readData_31_bm[9]_net_1\, 
        \readData_31_bm_1_1_RNO[9]_net_1\, 
        \readData_31_bm_1_1_RNO_0[9]_net_1\, 
        \readData_31_am_RNO[10]_net_1\, 
        \readData_31_am_1_1[10]_net_1\, 
        \readData_31_am_RNO_0[10]_net_1\, 
        \readData_31_am[10]_net_1\, 
        \readData_31_am_1_1_RNO[10]_net_1\, 
        \readData_31_am_1_1_RNO_0[10]_net_1\, 
        \readData_31_bm_RNO[10]_net_1\, 
        \readData_31_bm_1_1[10]_net_1\, 
        \readData_31_bm_RNO_0[10]_net_1\, 
        \readData_31_bm[10]_net_1\, 
        \readData_31_bm_1_1_RNO[10]_net_1\, 
        \readData_31_bm_1_1_RNO_0[10]_net_1\, 
        \readData_31_am_RNO[11]_net_1\, 
        \readData_31_am_1_1[11]_net_1\, 
        \readData_31_am_RNO_0[11]_net_1\, 
        \readData_31_am[11]_net_1\, 
        \readData_31_am_1_1_RNO[11]_net_1\, 
        \readData_31_am_1_1_RNO_0[11]_net_1\, 
        \readData_31_bm_RNO[11]_net_1\, 
        \readData_31_bm_1_1[11]_net_1\, 
        \readData_31_bm_RNO_0[11]_net_1\, 
        \readData_31_bm[11]_net_1\, 
        \readData_31_bm_1_1_RNO[11]_net_1\, 
        \readData_31_bm_1_1_RNO_0[11]_net_1\, 
        \readData_31_am_RNO[12]_net_1\, 
        \readData_31_am_1_1[12]_net_1\, 
        \readData_31_am_RNO_0[12]_net_1\, 
        \readData_31_am[12]_net_1\, 
        \readData_31_am_1_1_RNO[12]_net_1\, 
        \readData_31_am_1_1_RNO_0[12]_net_1\, 
        \readData_31_bm_RNO[12]_net_1\, 
        \readData_31_bm_1_1[12]_net_1\, 
        \readData_31_bm_RNO_0[12]_net_1\, 
        \readData_31_bm[12]_net_1\, 
        \readData_31_bm_1_1_RNO[12]_net_1\, 
        \readData_31_bm_1_1_RNO_0[12]_net_1\, 
        \readData_31_am_RNO[13]_net_1\, 
        \readData_31_am_1_1[13]_net_1\, 
        \readData_31_am_RNO_0[13]_net_1\, 
        \readData_31_am[13]_net_1\, 
        \readData_31_am_1_1_RNO[13]_net_1\, 
        \readData_31_am_1_1_RNO_0[13]_net_1\, 
        \readData_31_bm_RNO[13]_net_1\, 
        \readData_31_bm_1_1[13]_net_1\, 
        \readData_31_bm_RNO_0[13]_net_1\, 
        \readData_31_bm[13]_net_1\, 
        \readData_31_bm_1_1_RNO[13]_net_1\, 
        \readData_31_bm_1_1_RNO_0[13]_net_1\, 
        \readData_31_am_RNO[14]_net_1\, 
        \readData_31_am_1_1[14]_net_1\, 
        \readData_31_am_RNO_0[14]_net_1\, 
        \readData_31_am[14]_net_1\, 
        \readData_31_am_1_1_RNO[14]_net_1\, 
        \readData_31_am_1_1_RNO_0[14]_net_1\, 
        \readData_31_bm_RNO[14]_net_1\, 
        \readData_31_bm_1_1[14]_net_1\, 
        \readData_31_bm_RNO_0[14]_net_1\, 
        \readData_31_bm[14]_net_1\, 
        \readData_31_bm_1_1_RNO[14]_net_1\, 
        \readData_31_bm_1_1_RNO_0[14]_net_1\, 
        \readData_31_am_RNO[15]_net_1\, 
        \readData_31_am_1_1[15]_net_1\, 
        \readData_31_am_RNO_0[15]_net_1\, 
        \readData_31_am[15]_net_1\, 
        \readData_31_am_1_1_RNO[15]_net_1\, 
        \readData_31_am_1_1_RNO_0[15]_net_1\, 
        \readData_31_bm_RNO[15]_net_1\, 
        \readData_31_bm_1_1[15]_net_1\, 
        \readData_31_bm_RNO_0[15]_net_1\, 
        \readData_31_bm[15]_net_1\, 
        \readData_31_bm_1_1_RNO[15]_net_1\, 
        \readData_31_bm_1_1_RNO_0[15]_net_1\, 
        \readData_31_am_RNO[16]_net_1\, 
        \readData_31_am_1_1[16]_net_1\, 
        \readData_31_am_RNO_0[16]_net_1\, 
        \readData_31_am[16]_net_1\, 
        \readData_31_am_1_1_RNO[16]_net_1\, 
        \readData_31_am_1_1_RNO_0[16]_net_1\, 
        \readData_31_bm_RNO[16]_net_1\, 
        \readData_31_bm_1_1[16]_net_1\, 
        \readData_31_bm_RNO_0[16]_net_1\, 
        \readData_31_bm[16]_net_1\, 
        \readData_31_bm_1_1_RNO[16]_net_1\, 
        \readData_31_bm_1_1_RNO_0[16]_net_1\, 
        \readData_31_am_RNO[17]_net_1\, 
        \readData_31_am_1_1[17]_net_1\, 
        \readData_31_am_RNO_0[17]_net_1\, 
        \readData_31_am[17]_net_1\, 
        \readData_31_am_1_1_RNO[17]_net_1\, 
        \readData_31_am_1_1_RNO_0[17]_net_1\, 
        \readData_31_bm_RNO[17]_net_1\, 
        \readData_31_bm_1_1[17]_net_1\, 
        \readData_31_bm_RNO_0[17]_net_1\, 
        \readData_31_bm[17]_net_1\, 
        \readData_31_bm_1_1_RNO[17]_net_1\, 
        \readData_31_bm_1_1_RNO_0[17]_net_1\, 
        \readData_31_am_RNO[18]_net_1\, 
        \readData_31_am_1_1[18]_net_1\, 
        \readData_31_am_RNO_0[18]_net_1\, 
        \readData_31_am[18]_net_1\, 
        \readData_31_am_1_1_RNO[18]_net_1\, 
        \readData_31_am_1_1_RNO_0[18]_net_1\, 
        \readData_31_bm_RNO[18]_net_1\, 
        \readData_31_bm_1_1[18]_net_1\, 
        \readData_31_bm_RNO_0[18]_net_1\, 
        \readData_31_bm[18]_net_1\, 
        \readData_31_bm_1_1_RNO[18]_net_1\, 
        \readData_31_bm_1_1_RNO_0[18]_net_1\, 
        \readData_31_am_RNO[19]_net_1\, 
        \readData_31_am_1_1[19]_net_1\, 
        \readData_31_am_RNO_0[19]_net_1\, 
        \readData_31_am[19]_net_1\, 
        \readData_31_am_1_1_RNO[19]_net_1\, 
        \readData_31_am_1_1_RNO_0[19]_net_1\, 
        \readData_31_bm_RNO[19]_net_1\, 
        \readData_31_bm_1_1[19]_net_1\, 
        \readData_31_bm_RNO_0[19]_net_1\, 
        \readData_31_bm[19]_net_1\, 
        \readData_31_bm_1_1_RNO[19]_net_1\, 
        \readData_31_bm_1_1_RNO_0[19]_net_1\, 
        \readData_31_am_RNO[20]_net_1\, 
        \readData_31_am_1_1[20]_net_1\, 
        \readData_31_am_RNO_0[20]_net_1\, 
        \readData_31_am[20]_net_1\, 
        \readData_31_am_1_1_RNO[20]_net_1\, 
        \readData_31_am_1_1_RNO_0[20]_net_1\, 
        \readData_31_bm_RNO[20]_net_1\, 
        \readData_31_bm_1_1[20]_net_1\, 
        \readData_31_bm_RNO_0[20]_net_1\, 
        \readData_31_bm[20]_net_1\, 
        \readData_31_bm_1_1_RNO[20]_net_1\, 
        \readData_31_bm_1_1_RNO_0[20]_net_1\, 
        \readData_31_am_RNO[21]_net_1\, 
        \readData_31_am_1_1[21]_net_1\, 
        \readData_31_am_RNO_0[21]_net_1\, 
        \readData_31_am[21]_net_1\, 
        \readData_31_am_1_1_RNO[21]_net_1\, 
        \readData_31_am_1_1_RNO_0[21]_net_1\, 
        \readData_31_bm_RNO[21]_net_1\, 
        \readData_31_bm_1_1[21]_net_1\, 
        \readData_31_bm_RNO_0[21]_net_1\, 
        \readData_31_bm[21]_net_1\, 
        \readData_31_bm_1_1_RNO[21]_net_1\, 
        \readData_31_bm_1_1_RNO_0[21]_net_1\, 
        \readData_31_am_RNO[22]_net_1\, 
        \readData_31_am_1_1[22]_net_1\, 
        \readData_31_am_RNO_0[22]_net_1\, 
        \readData_31_am[22]_net_1\, 
        \readData_31_am_1_1_RNO[22]_net_1\, 
        \readData_31_am_1_1_RNO_0[22]_net_1\, 
        \readData_31_bm_RNO[22]_net_1\, 
        \readData_31_bm_1_1[22]_net_1\, 
        \readData_31_bm_RNO_0[22]_net_1\, 
        \readData_31_bm[22]_net_1\, 
        \readData_31_bm_1_1_RNO[22]_net_1\, 
        \readData_31_bm_1_1_RNO_0[22]_net_1\, 
        \readData_31_am_RNO[23]_net_1\, 
        \readData_31_am_1_1[23]_net_1\, 
        \readData_31_am_RNO_0[23]_net_1\, 
        \readData_31_am[23]_net_1\, 
        \readData_31_am_1_1_RNO[23]_net_1\, 
        \readData_31_am_1_1_RNO_0[23]_net_1\, 
        \readData_31_bm_RNO[23]_net_1\, 
        \readData_31_bm_1_1[23]_net_1\, 
        \readData_31_bm_RNO_0[23]_net_1\, 
        \readData_31_bm[23]_net_1\, 
        \readData_31_bm_1_1_RNO[23]_net_1\, 
        \readData_31_bm_1_1_RNO_0[23]_net_1\, 
        \readData_31_am_RNO[24]_net_1\, 
        \readData_31_am_1_1[24]_net_1\, 
        \readData_31_am_RNO_0[24]_net_1\, 
        \readData_31_am[24]_net_1\, 
        \readData_31_am_1_1_RNO[24]_net_1\, 
        \readData_31_am_1_1_RNO_0[24]_net_1\, 
        \readData_31_bm_RNO[24]_net_1\, 
        \readData_31_bm_1_1[24]_net_1\, 
        \readData_31_bm_RNO_0[24]_net_1\, 
        \readData_31_bm[24]_net_1\, 
        \readData_31_bm_1_1_RNO[24]_net_1\, 
        \readData_31_bm_1_1_RNO_0[24]_net_1\, 
        \readData_31_am_RNO[25]_net_1\, 
        \readData_31_am_1_1[25]_net_1\, 
        \readData_31_am_RNO_0[25]_net_1\, 
        \readData_31_am[25]_net_1\, 
        \readData_31_am_1_1_RNO[25]_net_1\, 
        \readData_31_am_1_1_RNO_0[25]_net_1\, 
        \readData_31_bm_RNO[25]_net_1\, 
        \readData_31_bm_1_1[25]_net_1\, 
        \readData_31_bm_RNO_0[25]_net_1\, 
        \readData_31_bm[25]_net_1\, 
        \readData_31_bm_1_1_RNO[25]_net_1\, 
        \readData_31_bm_1_1_RNO_0[25]_net_1\, 
        \readData_31_am_RNO[26]_net_1\, 
        \readData_31_am_1_1[26]_net_1\, 
        \readData_31_am_RNO_0[26]_net_1\, 
        \readData_31_am[26]_net_1\, 
        \readData_31_am_1_1_RNO[26]_net_1\, 
        \readData_31_am_1_1_RNO_0[26]_net_1\, 
        \readData_31_bm_RNO[26]_net_1\, 
        \readData_31_bm_1_1[26]_net_1\, 
        \readData_31_bm_RNO_0[26]_net_1\, 
        \readData_31_bm[26]_net_1\, 
        \readData_31_bm_1_1_RNO[26]_net_1\, 
        \readData_31_bm_1_1_RNO_0[26]_net_1\, 
        \readData_31_am_RNO[27]_net_1\, 
        \readData_31_am_1_1[27]_net_1\, 
        \readData_31_am_RNO_0[27]_net_1\, 
        \readData_31_am[27]_net_1\, 
        \readData_31_am_1_1_RNO[27]_net_1\, 
        \readData_31_am_1_1_RNO_0[27]_net_1\, 
        \readData_31_bm_RNO[27]_net_1\, 
        \readData_31_bm_1_1[27]_net_1\, 
        \readData_31_bm_RNO_0[27]_net_1\, 
        \readData_31_bm[27]_net_1\, 
        \readData_31_bm_1_1_RNO[27]_net_1\, 
        \readData_31_bm_1_1_RNO_0[27]_net_1\, 
        \readData_31_am_RNO[28]_net_1\, 
        \readData_31_am_1_1[28]_net_1\, 
        \readData_31_am_RNO_0[28]_net_1\, 
        \readData_31_am[28]_net_1\, 
        \readData_31_am_1_1_RNO[28]_net_1\, 
        \readData_31_am_1_1_RNO_0[28]_net_1\, 
        \readData_31_bm_RNO[28]_net_1\, 
        \readData_31_bm_1_1[28]_net_1\, 
        \readData_31_bm_RNO_0[28]_net_1\, 
        \readData_31_bm[28]_net_1\, 
        \readData_31_bm_1_1_RNO[28]_net_1\, 
        \readData_31_bm_1_1_RNO_0[28]_net_1\, 
        \readData_31_am_RNO[29]_net_1\, 
        \readData_31_am_1_1[29]_net_1\, 
        \readData_31_am_RNO_0[29]_net_1\, 
        \readData_31_am[29]_net_1\, 
        \readData_31_am_1_1_RNO[29]_net_1\, 
        \readData_31_am_1_1_RNO_0[29]_net_1\, 
        \readData_31_bm_RNO[29]_net_1\, 
        \readData_31_bm_1_1[29]_net_1\, 
        \readData_31_bm_RNO_0[29]_net_1\, 
        \readData_31_bm[29]_net_1\, 
        \readData_31_bm_1_1_RNO[29]_net_1\, 
        \readData_31_bm_1_1_RNO_0[29]_net_1\, 
        \readData_31_am_RNO[30]_net_1\, 
        \readData_31_am_1_1[30]_net_1\, 
        \readData_31_am_RNO_0[30]_net_1\, 
        \readData_31_am[30]_net_1\, 
        \readData_31_am_1_1_RNO[30]_net_1\, 
        \readData_31_am_1_1_RNO_0[30]_net_1\, 
        \readData_31_bm_RNO[30]_net_1\, 
        \readData_31_bm_1_1[30]_net_1\, 
        \readData_31_bm_RNO_0[30]_net_1\, 
        \readData_31_bm[30]_net_1\, 
        \readData_31_bm_1_1_RNO[30]_net_1\, 
        \readData_31_bm_1_1_RNO_0[30]_net_1\, 
        \readData_31_am_RNO[31]_net_1\, 
        \readData_31_am_1_1[31]_net_1\, 
        \readData_31_am_RNO_0[31]_net_1\, 
        \readData_31_am[31]_net_1\, 
        \readData_31_am_1_1_RNO[31]_net_1\, 
        \readData_31_am_1_1_RNO_0[31]_net_1\, 
        \readData_31_bm_RNO[31]_net_1\, 
        \readData_31_bm_1_1[31]_net_1\, 
        \readData_31_bm_RNO_0[31]_net_1\, 
        \readData_31_bm[31]_net_1\, 
        \readData_31_bm_1_1_RNO[31]_net_1\, 
        \readData_31_bm_1_1_RNO_0[31]_net_1\, \readData30[7]\, 
        \readData_13_1_1[7]\, \readData14[7]\, \readData22[7]\, 
        \readData6[7]\, \readData30[6]\, \readData_13_1_1[6]\, 
        \readData14[6]\, \readData22[6]\, \readData6[6]\, 
        \readData31[7]\, \readData_28_1_1[7]\, \readData15[7]\, 
        \readData23[7]\, \readData7[7]\, \readData28[2]\, 
        \readData_6_1_1[2]\, \readData12[2]\, \readData20[2]\, 
        \readData4[2]\, \readData30[5]\, \readData_13_1_1[5]\, 
        \readData14[5]\, \readData22[5]\, \readData6[5]\, 
        \readData28[4]\, \readData_6_1_1[4]\, \readData12[4]\, 
        \readData20[4]\, \readData4[4]\, \readData31[9]\, 
        \readData_28_1_1[8]\, \readData15[9]\, \readData23[9]\, 
        \readData7[9]\, \readData31[10]\, \readData_28_1_1[9]\, 
        \readData15[10]\, \readData23[10]\, \readData7[10]\, 
        \readData30[4]\, \readData_13_1_1[4]\, \readData14[4]\, 
        \readData22[4]\, \readData6[4]\, \readData28[9]\, 
        \readData_6_1_1[8]\, \readData12[9]\, \readData20[9]\, 
        \readData4[9]\, \readData28[5]\, \readData_6_1_1[5]\, 
        \readData12[5]\, \readData20[5]\, \readData4[5]\, 
        \readData28[6]\, \readData_6_1_1[6]\, \readData12[6]\, 
        \readData20[6]\, \readData4[6]\, \readData28[3]\, 
        \readData_6_1_1[3]\, \readData12[3]\, \readData20[3]\, 
        \readData4[3]\, \readData30[3]\, \readData_13_1_1[3]\, 
        \readData14[3]\, \readData22[3]\, \readData6[3]\, 
        \readData30[19]\, \readData_13_1_1[17]\, \readData14[19]\, 
        \readData22[19]\, \readData6[19]\, \readData28[0]\, 
        \readData_6_1_1[0]\, \readData12[0]\, \readData20[0]\, 
        \readData4[0]\, \readData28[7]\, \readData_6_1_1[7]\, 
        \readData12[7]\, \readData20[7]\, \readData4[7]\, 
        \readData31[11]\, \readData_28_1_1[10]\, \readData15[11]\, 
        \readData23[11]\, \readData7[11]\, \readData30[9]\, 
        \readData_13_1_1[8]\, \readData14[9]\, \readData22[9]\, 
        \readData6[9]\, \readData30[10]\, \readData_13_1_1[9]\, 
        \readData14[10]\, \readData22[10]\, \readData6[10]\, 
        \readData28[1]\, \readData_6_1_1[1]\, \readData12[1]\, 
        \readData20[1]\, \readData4[1]\, \readData30[12]\, 
        \readData_13_1_1[11]\, \readData14[12]\, \readData22[12]\, 
        \readData6[12]\, \readData30[13]\, \readData_13_1_1[12]\, 
        \readData14[13]\, \readData22[13]\, \readData6[13]\, 
        \readData28[10]\, \readData_6_1_1[9]\, \readData12[10]\, 
        \readData20[10]\, \readData4[10]\, \readData30[11]\, 
        \readData_13_1_1[10]\, \readData14[11]\, \readData22[11]\, 
        \readData6[11]\, \readData26[2]\, \readData_10_1_1[2]\, 
        \readData10[2]\, \readData18[2]\, \readData2[2]\, 
        \readData28[11]\, \readData_6_1_1[10]\, \readData12[11]\, 
        \readData20[11]\, \readData4[11]\, \readData28[12]\, 
        \readData_6_1_1[11]\, \readData12[12]\, \readData20[12]\, 
        \readData4[12]\, \readData28[13]\, \readData_6_1_1[12]\, 
        \readData12[13]\, \readData20[13]\, \readData4[13]\, 
        \readData28[14]\, \readData_6_1_1[13]\, \readData12[14]\, 
        \readData20[14]\, \readData4[14]\, \readData30[21]\, 
        \readData_13_1_1[19]\, \readData14[21]\, \readData22[21]\, 
        \readData6[21]\, \readData30[22]\, \readData_13_1_1[20]\, 
        \readData14[22]\, \readData22[22]\, \readData6[22]\, 
        \readData30[23]\, \readData_13_1_1[21]\, \readData14[23]\, 
        \readData22[23]\, \readData6[23]\, \readData30[24]\, 
        \readData_13_1_1[22]\, \readData14[24]\, \readData22[24]\, 
        \readData6[24]\, \readData30[25]\, \readData_13_1_1[23]\, 
        \readData14[25]\, \readData22[25]\, \readData6[25]\, 
        \readData30[27]\, \readData_13_1_1[24]\, \readData14[27]\, 
        \readData22[27]\, \readData6[27]\, \readData26[0]\, 
        \readData_10_1_1[0]\, \readData10[0]\, \readData18[0]\, 
        \readData2[0]\, \readData26[1]\, \readData_10_1_1[1]\, 
        \readData10[1]\, \readData18[1]\, \readData2[1]\, 
        \readData30[0]\, \readData_13_1_1[0]\, \readData14[0]\, 
        \readData22[0]\, \readData6[0]\, \readData30[1]\, 
        \readData_13_1_1[1]\, \readData14[1]\, \readData22[1]\, 
        \readData6[1]\, \readData30[2]\, \readData_13_1_1[2]\, 
        \readData14[2]\, \readData22[2]\, \readData6[2]\, 
        \readData31[6]\, \readData_28_1_1[6]\, \readData15[6]\, 
        \readData23[6]\, \readData7[6]\, \readData24[0]\, 
        \readData_3_1_1[0]\, \readData8[0]\, \readData16[0]\, 
        \readData0[0]\, \readData24[1]\, \readData_3_1_1[1]\, 
        \readData8[1]\, \readData16[1]\, \readData0[1]\, 
        \readData24[2]\, \readData_3_1_1[2]\, \readData8[2]\, 
        \readData16[2]\, \readData0[2]\, \readData31[12]\, 
        \readData_28_1_1[11]\, \readData15[12]\, \readData23[12]\, 
        \readData7[12]\, \readData31[13]\, \readData_28_1_1[12]\, 
        \readData15[13]\, \readData23[13]\, \readData7[13]\, 
        \readData31[14]\, \readData_28_1_1[13]\, \readData15[14]\, 
        \readData23[14]\, \readData7[14]\, \readData31[15]\, 
        \readData_28_1_1[14]\, \readData15[15]\, \readData23[15]\, 
        \readData7[15]\, \readData31[16]\, \readData_28_1_1[15]\, 
        \readData15[16]\, \readData23[16]\, \readData7[16]\, 
        \readData30[14]\, \readData_13_1_1[13]\, \readData14[14]\, 
        \readData22[14]\, \readData6[14]\, \readData30[15]\, 
        \readData_13_1_1[14]\, \readData14[15]\, \readData22[15]\, 
        \readData6[15]\, \readData30[16]\, \readData_13_1_1[15]\, 
        \readData14[16]\, \readData22[16]\, \readData6[16]\, 
        \readData30[18]\, \readData_13_1_1[16]\, \readData14[18]\, 
        \readData22[18]\, \readData6[18]\, \readData29[2]\, 
        \readData_21_1_1[2]\, \readData13[2]\, \readData21[2]\, 
        \readData5[2]\, \readData29[3]\, \readData_21_1_1[3]\, 
        \readData13[3]\, \readData21[3]\, \readData5[3]\, 
        \readData30[20]\, \readData_13_1_1[18]\, \readData14[20]\, 
        \readData22[20]\, \readData6[20]\, \readData29[4]\, 
        \readData_21_1_1[4]\, \readData13[4]\, \readData21[4]\, 
        \readData5[4]\, \readData29[5]\, \readData_21_1_1[5]\, 
        \readData13[5]\, \readData21[5]\, \readData5[5]\, 
        \readData29[6]\, \readData_21_1_1[6]\, \readData13[6]\, 
        \readData21[6]\, \readData5[6]\, \readData29[7]\, 
        \readData_21_1_1[7]\, \readData13[7]\, \readData21[7]\, 
        \readData5[7]\, \readData29[9]\, \readData_21_1_1[8]\, 
        \readData13[9]\, \readData21[9]\, \readData5[9]\, 
        \readData29[10]\, \readData_21_1_1[9]\, \readData13[10]\, 
        \readData21[10]\, \readData5[10]\, \readData29[11]\, 
        \readData_21_1_1[10]\, \readData13[11]\, \readData21[11]\, 
        \readData5[11]\, \readData30[28]\, \readData_13_1_1[25]\, 
        \readData14[28]\, \readData22[28]\, \readData6[28]\, 
        \readData30[29]\, \readData_13_1_1[26]\, \readData14[29]\, 
        \readData22[29]\, \readData6[29]\, \readData30[30]\, 
        \readData_13_1_1[27]\, \readData14[30]\, \readData22[30]\, 
        \readData6[30]\, \readData26[3]\, \readData_10_1_1[3]\, 
        \readData10[3]\, \readData18[3]\, \readData2[3]\, 
        \readData26[4]\, \readData_10_1_1[4]\, \readData10[4]\, 
        \readData18[4]\, \readData2[4]\, \readData26[5]\, 
        \readData_10_1_1[5]\, \readData10[5]\, \readData18[5]\, 
        \readData2[5]\, \readData26[6]\, \readData_10_1_1[6]\, 
        \readData10[6]\, \readData18[6]\, \readData2[6]\, 
        \readData28[15]\, \readData_6_1_1[14]\, \readData12[15]\, 
        \readData20[15]\, \readData4[15]\, \readData28[16]\, 
        \readData_6_1_1[15]\, \readData12[16]\, \readData20[16]\, 
        \readData4[16]\, \readData28[18]\, \readData_6_1_1[16]\, 
        \readData12[18]\, \readData20[18]\, \readData4[18]\, 
        \readData31[0]\, \readData_28_1_1[0]\, \readData15[0]\, 
        \readData23[0]\, \readData7[0]\, \readData31[1]\, 
        \readData_28_1_1[1]\, \readData15[1]\, \readData23[1]\, 
        \readData7[1]\, \readData31[2]\, \readData_28_1_1[2]\, 
        \readData15[2]\, \readData23[2]\, \readData7[2]\, 
        \readData31[3]\, \readData_28_1_1[3]\, \readData15[3]\, 
        \readData23[3]\, \readData7[3]\, \readData28[23]\, 
        \readData_6_1_1[21]\, \readData12[23]\, \readData20[23]\, 
        \readData4[23]\, \readData31[4]\, \readData_28_1_1[4]\, 
        \readData15[4]\, \readData23[4]\, \readData7[4]\, 
        \readData31[5]\, \readData_28_1_1[5]\, \readData15[5]\, 
        \readData23[5]\, \readData7[5]\, \readData28[27]\, 
        \readData_6_1_1[24]\, \readData12[27]\, \readData20[27]\, 
        \readData4[27]\, \readData26[19]\, \readData_10_1_1[17]\, 
        \readData10[19]\, \readData18[19]\, \readData2[19]\, 
        \readData28[28]\, \readData_6_1_1[25]\, \readData12[28]\, 
        \readData20[28]\, \readData4[28]\, \readData28[29]\, 
        \readData_6_1_1[26]\, \readData12[29]\, \readData20[29]\, 
        \readData4[29]\, \readData28[30]\, \readData_6_1_1[27]\, 
        \readData12[30]\, \readData20[30]\, \readData4[30]\, 
        \readData24[3]\, \readData_3_1_1[3]\, \readData8[3]\, 
        \readData16[3]\, \readData0[3]\, \readData24[4]\, 
        \readData_3_1_1[4]\, \readData8[4]\, \readData16[4]\, 
        \readData0[4]\, \readData24[5]\, \readData_3_1_1[5]\, 
        \readData8[5]\, \readData16[5]\, \readData0[5]\, 
        \readData24[6]\, \readData_3_1_1[6]\, \readData8[6]\, 
        \readData16[6]\, \readData0[6]\, \readData31[18]\, 
        \readData_28_1_1[16]\, \readData15[18]\, \readData23[18]\, 
        \readData7[18]\, \readData31[19]\, \readData_28_1_1[17]\, 
        \readData15[19]\, \readData23[19]\, \readData7[19]\, 
        \readData29[0]\, \readData_21_1_1[0]\, \readData13[0]\, 
        \readData21[0]\, \readData5[0]\, \readData29[1]\, 
        \readData_21_1_1[1]\, \readData13[1]\, \readData21[1]\, 
        \readData5[1]\, \readData31[21]\, \readData_28_1_1[19]\, 
        \readData15[21]\, \readData23[21]\, \readData7[21]\, 
        \readData31[22]\, \readData_28_1_1[20]\, \readData15[22]\, 
        \readData23[22]\, \readData7[22]\, \readData31[23]\, 
        \readData_28_1_1[21]\, \readData15[23]\, \readData23[23]\, 
        \readData7[23]\, \readData24[14]\, \readData_3_1_1[13]\, 
        \readData8[14]\, \readData16[14]\, \readData0[14]\, 
        \readData31[24]\, \readData_28_1_1[22]\, \readData15[24]\, 
        \readData23[24]\, \readData7[24]\, \readData31[25]\, 
        \readData_28_1_1[23]\, \readData15[25]\, \readData23[25]\, 
        \readData7[25]\, \readData31[27]\, \readData_28_1_1[24]\, 
        \readData15[27]\, \readData23[27]\, \readData7[27]\, 
        \readData27[0]\, \readData_25_1_1[0]\, \readData11[0]\, 
        \readData19[0]\, \readData3[0]\, \readData27[1]\, 
        \readData_25_1_1[1]\, \readData11[1]\, \readData19[1]\, 
        \readData3[1]\, \readData27[2]\, \readData_25_1_1[2]\, 
        \readData11[2]\, \readData19[2]\, \readData3[2]\, 
        \readData27[3]\, \readData_25_1_1[3]\, \readData11[3]\, 
        \readData19[3]\, \readData3[3]\, \readData29[12]\, 
        \readData_21_1_1[11]\, \readData13[12]\, \readData21[12]\, 
        \readData5[12]\, \readData29[13]\, \readData_21_1_1[12]\, 
        \readData13[13]\, \readData21[13]\, \readData5[13]\, 
        \readData29[14]\, \readData_21_1_1[13]\, \readData13[14]\, 
        \readData21[14]\, \readData5[14]\, \readData30[31]\, 
        \readData_13_1_1[28]\, \readData14[31]\, \readData22[31]\, 
        \readData6[31]\, \readData30[32]\, \readData_13_1_1[29]\, 
        \readData14[32]\, \readData22[32]\, \readData6[32]\, 
        \readData30[33]\, \readData_13_1_1[30]\, \readData14[33]\, 
        \readData22[33]\, \readData6[33]\, \readData30[34]\, 
        \readData_13_1_1[31]\, \readData14[34]\, \readData22[34]\, 
        \readData6[34]\, \readData26[7]\, \readData_10_1_1[7]\, 
        \readData10[7]\, \readData18[7]\, \readData2[7]\, 
        \readData26[9]\, \readData_10_1_1[8]\, \readData10[9]\, 
        \readData18[9]\, \readData2[9]\, \readData28[19]\, 
        \readData_6_1_1[17]\, \readData12[19]\, \readData20[19]\, 
        \readData4[19]\, \readData28[20]\, \readData_6_1_1[18]\, 
        \readData12[20]\, \readData20[20]\, \readData4[20]\, 
        \readData28[21]\, \readData_6_1_1[19]\, \readData12[21]\, 
        \readData20[21]\, \readData4[21]\, \readData28[22]\, 
        \readData_6_1_1[20]\, \readData12[22]\, \readData20[22]\, 
        \readData4[22]\, \readData26[14]\, \readData_10_1_1[13]\, 
        \readData10[14]\, \readData18[14]\, \readData2[14]\, 
        \readData28[24]\, \readData_6_1_1[22]\, \readData12[24]\, 
        \readData20[24]\, \readData4[24]\, \readData28[25]\, 
        \readData_6_1_1[23]\, \readData12[25]\, \readData20[25]\, 
        \readData4[25]\, \readData26[18]\, \readData_10_1_1[16]\, 
        \readData10[18]\, \readData18[18]\, \readData2[18]\, 
        \readData25[2]\, \readData_18_1_1[2]\, \readData9[2]\, 
        \readData17[2]\, \readData1[2]\, \readData25[3]\, 
        \readData_18_1_1[3]\, \readData9[3]\, \readData17[3]\, 
        \readData1[3]\, \readData26[20]\, \readData_10_1_1[18]\, 
        \readData10[20]\, \readData18[20]\, \readData2[20]\, 
        \readData26[21]\, \readData_10_1_1[19]\, \readData10[21]\, 
        \readData18[21]\, \readData2[21]\, \readData26[22]\, 
        \readData_10_1_1[20]\, \readData10[22]\, \readData18[22]\, 
        \readData2[22]\, \readData28[31]\, \readData_6_1_1[28]\, 
        \readData12[31]\, \readData20[31]\, \readData4[31]\, 
        \readData28[32]\, \readData_6_1_1[29]\, \readData12[32]\, 
        \readData20[32]\, \readData4[32]\, \readData28[33]\, 
        \readData_6_1_1[30]\, \readData12[33]\, \readData20[33]\, 
        \readData4[33]\, \readData28[34]\, \readData_6_1_1[31]\, 
        \readData12[34]\, \readData20[34]\, \readData4[34]\, 
        \readData24[7]\, \readData_3_1_1[7]\, \readData8[7]\, 
        \readData16[7]\, \readData0[7]\, \readData24[9]\, 
        \readData_3_1_1[8]\, \readData8[9]\, \readData16[9]\, 
        \readData0[9]\, \readData31[20]\, \readData_28_1_1[18]\, 
        \readData15[20]\, \readData23[20]\, \readData7[20]\, 
        \readData24[11]\, \readData_3_1_1[10]\, \readData8[11]\, 
        \readData16[11]\, \readData0[11]\, \readData24[12]\, 
        \readData_3_1_1[11]\, \readData8[12]\, \readData16[12]\, 
        \readData0[12]\, \readData24[13]\, \readData_3_1_1[12]\, 
        \readData8[13]\, \readData16[13]\, \readData0[13]\, 
        \readData26[33]\, \readData_10_1_1[30]\, \readData10[33]\, 
        \readData18[33]\, \readData2[33]\, \readData24[15]\, 
        \readData_3_1_1[14]\, \readData8[15]\, \readData16[15]\, 
        \readData0[15]\, \readData24[16]\, \readData_3_1_1[15]\, 
        \readData8[16]\, \readData16[16]\, \readData0[16]\, 
        \readData24[18]\, \readData_3_1_1[16]\, \readData8[18]\, 
        \readData16[18]\, \readData0[18]\, \readData24[19]\, 
        \readData_3_1_1[17]\, \readData8[19]\, \readData16[19]\, 
        \readData0[19]\, \readData31[28]\, \readData_28_1_1[25]\, 
        \readData15[28]\, \readData23[28]\, \readData7[28]\, 
        \readData31[29]\, \readData_28_1_1[26]\, \readData15[29]\, 
        \readData23[29]\, \readData7[29]\, \readData31[30]\, 
        \readData_28_1_1[27]\, \readData15[30]\, \readData23[30]\, 
        \readData7[30]\, \readData31[31]\, \readData_28_1_1[28]\, 
        \readData15[31]\, \readData23[31]\, \readData7[31]\, 
        \readData27[4]\, \readData_25_1_1[4]\, \readData11[4]\, 
        \readData19[4]\, \readData3[4]\, \readData27[5]\, 
        \readData_25_1_1[5]\, \readData11[5]\, \readData19[5]\, 
        \readData3[5]\, \readData27[6]\, \readData_25_1_1[6]\, 
        \readData11[6]\, \readData19[6]\, \readData3[6]\, 
        \readData29[15]\, \readData_21_1_1[14]\, \readData13[15]\, 
        \readData21[15]\, \readData5[15]\, \readData29[16]\, 
        \readData_21_1_1[15]\, \readData13[16]\, \readData21[16]\, 
        \readData5[16]\, \readData29[18]\, \readData_21_1_1[16]\, 
        \readData13[18]\, \readData21[18]\, \readData5[18]\, 
        \readData29[19]\, \readData_21_1_1[17]\, \readData13[19]\, 
        \readData21[19]\, \readData5[19]\, \readData29[20]\, 
        \readData_21_1_1[18]\, \readData13[20]\, \readData21[20]\, 
        \readData5[20]\, \readData26[10]\, \readData_10_1_1[9]\, 
        \readData10[10]\, \readData18[10]\, \readData2[10]\, 
        \readData26[11]\, \readData_10_1_1[10]\, \readData10[11]\, 
        \readData18[11]\, \readData2[11]\, \readData26[12]\, 
        \readData_10_1_1[11]\, \readData10[12]\, \readData18[12]\, 
        \readData2[12]\, \readData26[13]\, \readData_10_1_1[12]\, 
        \readData10[13]\, \readData18[13]\, \readData2[13]\, 
        \readData29[25]\, \readData_21_1_1[23]\, \readData13[25]\, 
        \readData21[25]\, \readData5[25]\, \readData26[15]\, 
        \readData_10_1_1[14]\, \readData10[15]\, \readData18[15]\, 
        \readData2[15]\, \readData26[16]\, \readData_10_1_1[15]\, 
        \readData10[16]\, \readData18[16]\, \readData2[16]\, 
        \readData25[1]\, \readData_18_1_1[1]\, \readData9[1]\, 
        \readData17[1]\, \readData1[1]\, \readData29[29]\, 
        \readData_21_1_1[26]\, \readData13[29]\, \readData21[29]\, 
        \readData5[29]\, \readData29[30]\, \readData_21_1_1[27]\, 
        \readData13[30]\, \readData21[30]\, \readData5[30]\, 
        \readData29[31]\, \readData_21_1_1[28]\, \readData13[31]\, 
        \readData21[31]\, \readData5[31]\, \readData25[4]\, 
        \readData_18_1_1[4]\, \readData9[4]\, \readData17[4]\, 
        \readData1[4]\, \readData25[5]\, \readData_18_1_1[5]\, 
        \readData9[5]\, \readData17[5]\, \readData1[5]\, 
        \readData25[6]\, \readData_18_1_1[6]\, \readData9[6]\, 
        \readData17[6]\, \readData1[6]\, \readData26[23]\, 
        \readData_10_1_1[21]\, \readData10[23]\, \readData18[23]\, 
        \readData2[23]\, \readData26[24]\, \readData_10_1_1[22]\, 
        \readData10[24]\, \readData18[24]\, \readData2[24]\, 
        \readData26[25]\, \readData_10_1_1[23]\, \readData10[25]\, 
        \readData18[25]\, \readData2[25]\, \readData26[27]\, 
        \readData_10_1_1[24]\, \readData10[27]\, \readData18[27]\, 
        \readData2[27]\, \readData26[28]\, \readData_10_1_1[25]\, 
        \readData10[28]\, \readData18[28]\, \readData2[28]\, 
        \readData24[10]\, \readData_3_1_1[9]\, \readData8[10]\, 
        \readData16[10]\, \readData0[10]\, \readData26[30]\, 
        \readData_10_1_1[27]\, \readData10[30]\, \readData18[30]\, 
        \readData2[30]\, \readData26[31]\, \readData_10_1_1[28]\, 
        \readData10[31]\, \readData18[31]\, \readData2[31]\, 
        \readData26[32]\, \readData_10_1_1[29]\, \readData10[32]\, 
        \readData18[32]\, \readData2[32]\, \readData25[16]\, 
        \readData_18_1_1[15]\, \readData9[16]\, \readData17[16]\, 
        \readData1[16]\, \readData26[34]\, \readData_10_1_1[31]\, 
        \readData10[34]\, \readData18[34]\, \readData2[34]\, 
        \readData25[20]\, \readData_18_1_1[18]\, \readData9[20]\, 
        \readData17[20]\, \readData1[20]\, \readData25[21]\, 
        \readData_18_1_1[19]\, \readData9[21]\, \readData17[21]\, 
        \readData1[21]\, \readData25[22]\, \readData_18_1_1[20]\, 
        \readData9[22]\, \readData17[22]\, \readData1[22]\, 
        \readData24[20]\, \readData_3_1_1[18]\, \readData8[20]\, 
        \readData16[20]\, \readData0[20]\, \readData24[21]\, 
        \readData_3_1_1[19]\, \readData8[21]\, \readData16[21]\, 
        \readData0[21]\, \readData24[22]\, \readData_3_1_1[20]\, 
        \readData8[22]\, \readData16[22]\, \readData0[22]\, 
        \readData24[23]\, \readData_3_1_1[21]\, \readData8[23]\, 
        \readData16[23]\, \readData0[23]\, \readData24[24]\, 
        \readData_3_1_1[22]\, \readData8[24]\, \readData16[24]\, 
        \readData0[24]\, \readData24[25]\, \readData_3_1_1[23]\, 
        \readData8[25]\, \readData16[25]\, \readData0[25]\, 
        \readData24[27]\, \readData_3_1_1[24]\, \readData8[27]\, 
        \readData16[27]\, \readData0[27]\, \readData24[28]\, 
        \readData_3_1_1[25]\, \readData8[28]\, \readData16[28]\, 
        \readData0[28]\, \readData24[29]\, \readData_3_1_1[26]\, 
        \readData8[29]\, \readData16[29]\, \readData0[29]\, 
        \readData24[30]\, \readData_3_1_1[27]\, \readData8[30]\, 
        \readData16[30]\, \readData0[30]\, \readData24[31]\, 
        \readData_3_1_1[28]\, \readData8[31]\, \readData16[31]\, 
        \readData0[31]\, \readData24[32]\, \readData_3_1_1[29]\, 
        \readData8[32]\, \readData16[32]\, \readData0[32]\, 
        \readData29[21]\, \readData_21_1_1[19]\, \readData13[21]\, 
        \readData21[21]\, \readData5[21]\, \readData29[22]\, 
        \readData_21_1_1[20]\, \readData13[22]\, \readData21[22]\, 
        \readData5[22]\, \readData29[23]\, \readData_21_1_1[21]\, 
        \readData13[23]\, \readData21[23]\, \readData5[23]\, 
        \readData29[24]\, \readData_21_1_1[22]\, \readData13[24]\, 
        \readData21[24]\, \readData5[24]\, \readData27[16]\, 
        \readData_25_1_1[15]\, \readData11[16]\, \readData19[16]\, 
        \readData3[16]\, \readData29[27]\, \readData_21_1_1[24]\, 
        \readData13[27]\, \readData21[27]\, \readData5[27]\, 
        \readData25[0]\, \readData_18_1_1[0]\, \readData9[0]\, 
        \readData17[0]\, \readData1[0]\, \readData29[28]\, 
        \readData_21_1_1[25]\, \readData13[28]\, \readData21[28]\, 
        \readData5[28]\, \readData27[20]\, \readData_25_1_1[18]\, 
        \readData11[20]\, \readData19[20]\, \readData3[20]\, 
        \readData27[21]\, \readData_25_1_1[19]\, \readData11[21]\, 
        \readData19[21]\, \readData3[21]\, \readData27[22]\, 
        \readData_25_1_1[20]\, \readData11[22]\, \readData19[22]\, 
        \readData3[22]\, \readData27[23]\, \readData_25_1_1[21]\, 
        \readData11[23]\, \readData19[23]\, \readData3[23]\, 
        \readData29[32]\, \readData_21_1_1[29]\, \readData13[32]\, 
        \readData21[32]\, \readData5[32]\, \readData29[33]\, 
        \readData_21_1_1[30]\, \readData13[33]\, \readData21[33]\, 
        \readData5[33]\, \readData29[34]\, \readData_21_1_1[31]\, 
        \readData13[34]\, \readData21[34]\, \readData5[34]\, 
        \readData25[7]\, \readData_18_1_1[7]\, \readData9[7]\, 
        \readData17[7]\, \readData1[7]\, \readData25[9]\, 
        \readData_18_1_1[8]\, \readData9[9]\, \readData17[9]\, 
        \readData1[9]\, \readData25[10]\, \readData_18_1_1[9]\, 
        \readData9[10]\, \readData17[10]\, \readData1[10]\, 
        \readData25[11]\, \readData_18_1_1[10]\, \readData9[11]\, 
        \readData17[11]\, \readData1[11]\, \readData26[29]\, 
        \readData_10_1_1[26]\, \readData10[29]\, \readData18[29]\, 
        \readData2[29]\, \readData25[13]\, \readData_18_1_1[12]\, 
        \readData9[13]\, \readData17[13]\, \readData1[13]\, 
        \readData25[14]\, \readData_18_1_1[13]\, \readData9[14]\, 
        \readData17[14]\, \readData1[14]\, \readData25[15]\, 
        \readData_18_1_1[14]\, \readData9[15]\, \readData17[15]\, 
        \readData1[15]\, \readData27[7]\, \readData_25_1_1[7]\, 
        \readData11[7]\, \readData19[7]\, \readData3[7]\, 
        \readData25[18]\, \readData_18_1_1[16]\, \readData9[18]\, 
        \readData17[18]\, \readData1[18]\, \readData25[19]\, 
        \readData_18_1_1[17]\, \readData9[19]\, \readData17[19]\, 
        \readData1[19]\, \readData27[11]\, \readData_25_1_1[10]\, 
        \readData11[11]\, \readData19[11]\, \readData3[11]\, 
        \readData24[33]\, \readData_3_1_1[30]\, \readData8[33]\, 
        \readData16[33]\, \readData0[33]\, \readData25[23]\, 
        \readData_18_1_1[21]\, \readData9[23]\, \readData17[23]\, 
        \readData1[23]\, \readData25[24]\, \readData_18_1_1[22]\, 
        \readData9[24]\, \readData17[24]\, \readData1[24]\, 
        \readData25[25]\, \readData_18_1_1[23]\, \readData9[25]\, 
        \readData17[25]\, \readData1[25]\, \readData25[27]\, 
        \readData_18_1_1[24]\, \readData9[27]\, \readData17[27]\, 
        \readData1[27]\, \readData25[28]\, \readData_18_1_1[25]\, 
        \readData9[28]\, \readData17[28]\, \readData1[28]\, 
        \readData31[32]\, \readData_28_1_1[29]\, \readData15[32]\, 
        \readData23[32]\, \readData7[32]\, \readData31[33]\, 
        \readData_28_1_1[30]\, \readData15[33]\, \readData23[33]\, 
        \readData7[33]\, \readData31[34]\, \readData_28_1_1[31]\, 
        \readData15[34]\, \readData23[34]\, \readData7[34]\, 
        \readData27[34]\, \readData_25_1_1[31]\, \readData11[34]\, 
        \readData19[34]\, \readData3[34]\, \readData27[9]\, 
        \readData_25_1_1[8]\, \readData11[9]\, \readData19[9]\, 
        \readData3[9]\, \readData27[10]\, \readData_25_1_1[9]\, 
        \readData11[10]\, \readData19[10]\, \readData3[10]\, 
        \readData25[34]\, \readData_18_1_1[31]\, \readData9[34]\, 
        \readData17[34]\, \readData1[34]\, \readData27[24]\, 
        \readData_25_1_1[22]\, \readData11[24]\, \readData19[24]\, 
        \readData3[24]\, \readData24[34]\, \readData_3_1_1[31]\, 
        \readData8[34]\, \readData16[34]\, \readData0[34]\, 
        \readData27[14]\, \readData_25_1_1[13]\, \readData11[14]\, 
        \readData19[14]\, \readData3[14]\, \readData27[15]\, 
        \readData_25_1_1[14]\, \readData11[15]\, \readData19[15]\, 
        \readData3[15]\, \readData27[29]\, \readData_25_1_1[26]\, 
        \readData11[29]\, \readData19[29]\, \readData3[29]\, 
        \readData27[18]\, \readData_25_1_1[16]\, \readData11[18]\, 
        \readData19[18]\, \readData3[18]\, \readData27[19]\, 
        \readData_25_1_1[17]\, \readData11[19]\, \readData19[19]\, 
        \readData3[19]\, \readData27[32]\, \readData_25_1_1[29]\, 
        \readData11[32]\, \readData19[32]\, \readData3[32]\, 
        \readData27[33]\, \readData_25_1_1[30]\, \readData11[33]\, 
        \readData19[33]\, \readData3[33]\, \readData25[31]\, 
        \readData_18_1_1[28]\, \readData9[31]\, \readData17[31]\, 
        \readData1[31]\, \readData25[32]\, \readData_18_1_1[29]\, 
        \readData9[32]\, \readData17[32]\, \readData1[32]\, 
        \readData25[33]\, \readData_18_1_1[30]\, \readData9[33]\, 
        \readData17[33]\, \readData1[33]\, \readData27[28]\, 
        \readData_25_1_1[25]\, \readData11[28]\, \readData19[28]\, 
        \readData3[28]\, \readData25[30]\, \readData_18_1_1[27]\, 
        \readData9[30]\, \readData17[30]\, \readData1[30]\, 
        \readData27[25]\, \readData_25_1_1[23]\, \readData11[25]\, 
        \readData19[25]\, \readData3[25]\, \readData27[27]\, 
        \readData_25_1_1[24]\, \readData11[27]\, \readData19[27]\, 
        \readData3[27]\, \readData25[29]\, \readData_18_1_1[26]\, 
        \readData9[29]\, \readData17[29]\, \readData1[29]\, 
        \readData27[31]\, \readData_25_1_1[28]\, \readData11[31]\, 
        \readData19[31]\, \readData3[31]\, \readData27[30]\, 
        \readData_25_1_1[27]\, \readData11[30]\, \readData19[30]\, 
        \readData3[30]\, \readData25[12]\, \readData_18_1_1[11]\, 
        \readData9[12]\, \readData17[12]\, \readData1[12]\, 
        \readData27[13]\, \readData_25_1_1[12]\, \readData11[13]\, 
        \readData19[13]\, \readData3[13]\, \readData27[12]\, 
        \readData_25_1_1[11]\, \readData11[12]\, \readData19[12]\, 
        \readData3[12]\, readdata_xhdl1401_1, readdata_xhdl1414_1, 
        readdata_xhdl1403_0, N_1143, N_1147, N_1149, N_1150, 
        N_1144, N_1148, N_1168, wen_a3133, \wen_a5_1[1]\, 
        \wen_a5_1[0]\, \wen_a18_1[1]\, \wen_a18_1[0]\, 
        \wen_a13_1[1]\, \wen_a13_1[0]\, \wen_b5_1[1]\, 
        \wen_b5_1[0]\, \wen_b18_1[1]\, \wen_b18_1[0]\, 
        \wen_b13_1[1]\, \wen_b13_1[0]\, \wen_a4_1[1]\, 
        \wen_a4_1[0]\, \wen_a3_1[1]\, \wen_a3_1[0]\, 
        \wen_a2_1[1]\, \wen_a2_1[0]\, \wen_a1_1[1]\, 
        \wen_a1_1[0]\, \wen_a0_1[1]\, \wen_a0_1[0]\, 
        \wen_b31_1[1]\, \wen_b31_1[0]\, \wen_a31_1[1]\, 
        \wen_a31_1[0]\, \wen_a20_1[1]\, \wen_a20_1[0]\, 
        \wen_a19_1[1]\, \wen_a19_1[0]\, \wen_a17_1[1]\, 
        \wen_a17_1[0]\, \wen_a16_1[1]\, \wen_a16_1[0]\, 
        \wen_a12_1[1]\, \wen_a12_1[0]\, \wen_b4_1[1]\, 
        \wen_b4_1[0]\, \wen_b3_1[1]\, \wen_b3_1[0]\, 
        \wen_b2_1[1]\, \wen_b2_1[0]\, \wen_b0_1[1]\, 
        \wen_b0_1[0]\, \wen_b20_1[1]\, \wen_b20_1[0]\, 
        \wen_b19_1[1]\, \wen_b19_1[0]\, \wen_b17_1[1]\, 
        \wen_b17_1[0]\, \wen_b16_1[1]\, \wen_b16_1[0]\, 
        \wen_b12_1[1]\, \wen_b12_1[0]\, \wen_a30_1[1]\, 
        \wen_a30_1[0]\, \wen_a28_1[1]\, \wen_a28_1[0]\, 
        \wen_a26_1[1]\, \wen_a26_1[0]\, \wen_a24_1[1]\, 
        \wen_a24_1[0]\, \wen_a_m[1]\, \wen_a_m[0]\, 
        \wen_b30_1[1]\, \wen_b30_1[0]\, \wen_b29_1[1]\, 
        \wen_b29_1[0]\, \wen_b28_1[1]\, \wen_b28_1[0]\, 
        \wen_b27_1[1]\, \wen_b27_1[0]\, \wen_b26_1[1]\, 
        \wen_b26_1[0]\, \wen_b25_1[1]\, \wen_b25_1[0]\, 
        \wen_b24_1[1]\, \wen_b24_1[0]\, \wen_b23_1[1]\, 
        \wen_b23_1[0]\, \wen_b22_1[1]\, \wen_b22_1[0]\, 
        \wen_b_m[1]\, \wen_b_m[0]\, \wen_a6_1[1]\, \wen_a6_1[0]\, 
        \wen_a21_1[1]\, \wen_a21_1[0]\, \wen_a15_1[1]\, 
        \wen_a15_1[0]\, \wen_a14_1[1]\, \wen_a14_1[0]\, 
        \wen_a11_1[1]\, \wen_a11_1[0]\, \wen_a10_1[1]\, 
        \wen_a10_1[0]\, \wen_a9_1[1]\, \wen_a9_1[0]\, 
        \wen_a8_1[1]\, \wen_a8_1[0]\, \wen_a7_1[1]\, 
        \wen_a7_1[0]\, \wen_a29_1[1]\, \wen_a29_1[0]\, 
        \wen_a27_1[1]\, \wen_a27_1[0]\, \wen_a25_1[1]\, 
        \wen_a25_1[0]\, \wen_a23_1[1]\, \wen_a23_1[0]\, 
        \wen_b15_1[1]\, \wen_b15_1[0]\, \wen_b14_1[1]\, 
        \wen_b14_1[0]\, \wen_b11_1[1]\, \wen_b11_1[0]\, 
        \wen_b10_1[1]\, \wen_b10_1[0]\, \wen_b9_1[1]\, 
        \wen_b9_1[0]\, \wen_b8_1[1]\, \wen_b8_1[0]\, 
        \wen_b7_1[1]\, \wen_b7_1[0]\, \wen_b6_1[1]\, 
        \wen_b6_1[0]\, VCC_net_1, GND_net_1 : std_logic;
    signal nc123, nc121, nc47, nc113, nc111, nc34, nc98, nc89, 
        nc70, nc60, nc105, nc74, nc120, nc119, nc64, nc110, nc9, 
        nc92, nc91, nc13, nc23, nc55, nc80, nc33, nc84, nc16, 
        nc26, nc45, nc73, nc58, nc63, nc27, nc17, nc127, nc99, 
        nc126, nc117, nc36, nc116, nc48, nc37, nc5, nc103, nc101, 
        nc52, nc76, nc51, nc66, nc77, nc67, nc4, nc124, nc109, 
        nc42, nc114, nc100, nc83, nc41, nc90, nc94, nc122, nc112, 
        nc86, nc59, nc25, nc15, nc87, nc35, nc49, nc28, nc18, 
        nc128, nc107, nc118, nc106, nc75, nc65, nc38, nc93, nc1, 
        nc2, nc50, nc22, nc12, nc21, nc11, nc78, nc54, nc68, nc3, 
        nc32, nc104, nc40, nc31, nc96, nc44, nc7, nc97, nc85, 
        nc72, nc6, nc71, nc62, nc61, nc125, nc115, nc102, nc19, 
        nc29, nc88, nc53, nc39, nc8, nc82, nc108, nc81, nc79, 
        nc43, nc69, nc56, nc20, nc10, nc57, nc95, nc24, nc14, 
        nc46, nc30 : std_logic;

begin 


    block2_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(3), Y => \wen_b2_1[1]\);
    
    \readData_31_am_RNO_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[22]\, D => \readData6[22]\, Y => 
        \readData_13_1_1[20]\);
    
    \readData_31_am_RNO_0[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[10]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[9]\, D => \readData10[10]\, Y => 
        \readData_31_am_RNO_0[9]_net_1\);
    
    \readData_31_am_RNO_0[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[18]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[16]\, D => \readData10[18]\, Y => 
        \readData_31_am_RNO_0[16]_net_1\);
    
    \readData_31_am_1_1_RNO_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[22]\, D => \readData4[22]\, Y => 
        \readData_6_1_1[20]\);
    
    block28_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(3), Y => \wen_b28_1[1]\);
    
    \readData_31_bm[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[24]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[24]_net_1\, D
         => \readData_31_bm_RNO_0[24]_net_1\, Y => 
        \readData_31_bm[24]_net_1\);
    
    \readData_31_am_RNO_0[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[3]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[3]\, D => \readData10[3]\, Y => 
        \readData_31_am_RNO_0[3]_net_1\);
    
    \readData_31_am_1_1_RNO_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[1]\, D => \readData4[1]\, Y => 
        \readData_6_1_1[1]\);
    
    block19_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(2), Y => \wen_b19_1[0]\);
    
    \readData_31_am_RNO[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[22]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[20]\, D => \readData14[22]\, Y => 
        \readData_31_am_RNO[20]_net_1\);
    
    \readData_31_am_1_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[1]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[1]_net_1\, Y => 
        \readData_31_am_1_1[1]_net_1\);
    
    \readData_31_am_RNO[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[0]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[0]\, D => \readData14[0]\, Y => 
        \readData_31_am_RNO[0]_net_1\);
    
    \readData_31_bm_RNO_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[3]\, D => \readData7[3]\, Y => 
        \readData_28_1_1[3]\);
    
    \readData_31_am_1_1_RNO_2[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[5]\, D => \readData0[5]\, Y => 
        \readData_3_1_1[5]\);
    
    \readData_31_am[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[21]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[21]_net_1\, D
         => \readData_31_am_RNO_0[21]_net_1\, Y => 
        \readData_31_am[21]_net_1\);
    
    block28_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(0), Y => \wen_a28_1[0]\);
    
    \readData_31_am[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[23]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[23]_net_1\, D
         => \readData_31_am_RNO_0[23]_net_1\, Y => 
        \readData_31_am[23]_net_1\);
    
    block31_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(0), Y => \wen_a31_1[0]\);
    
    \readData_31_bm[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[26]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[26]_net_1\, D
         => \readData_31_bm_RNO_0[26]_net_1\, Y => 
        \readData_31_bm[26]_net_1\);
    
    \readData_31_am_1_1_RNO_2[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[27]\, D => \readData0[27]\, Y => 
        \readData_3_1_1[24]\);
    
    \readData_31_bm_RNO_2[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[0]\, D => \readData3[0]\, Y => 
        \readData_25_1_1[0]\);
    
    block7_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(2), Y => \wen_b7_1[0]\);
    
    \readData_31_am_RNO_0[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[21]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[19]\, D => \readData10[21]\, Y => 
        \readData_31_am_RNO_0[19]_net_1\);
    
    block6_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(1), Y => \wen_a6_1[1]\);
    
    \readData_31_am_1_1_RNO[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[9]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[8]\, D => \readData12[9]\, Y => 
        \readData_31_am_1_1_RNO[8]_net_1\);
    
    \readData_31_bm_RNO_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[0]\, D => \readData7[0]\, Y => 
        \readData_28_1_1[0]\);
    
    \readData_31_am_1_1_RNO_2[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[28]\, D => \readData0[28]\, Y => 
        \readData_3_1_1[25]\);
    
    \readData_31_am_RNO_2[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[29]\, D => \readData2[29]\, Y => 
        \readData_10_1_1[26]\);
    
    \readData_31_am_RNO_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[7]\, D => \readData6[7]\, Y => 
        \readData_13_1_1[7]\);
    
    \readData_31_am_RNO_0[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[15]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[14]\, D => \readData10[15]\, Y => 
        \readData_31_am_RNO_0[14]_net_1\);
    
    \readData_31_ns[22]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[22]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[22]_net_1\, Y => 
        ram_rdata(22));
    
    block2_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(0), Y => \wen_a2_1[0]\);
    
    block10_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(3), Y => \wen_b10_1[1]\);
    
    \readData_31_bm_RNO[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[19]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[17]\, D => \readData15[19]\, Y => 
        \readData_31_bm_RNO[17]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[14]\, D => \readData1[14]\, Y => 
        \readData_18_1_1[13]\);
    
    block1_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => sram_wen_mem(0), B => wen_a3133, Y => 
        \wen_a1_1[0]\);
    
    \readData_31_am_RNO[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[12]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[11]\, D => \readData14[12]\, Y => 
        \readData_31_am_RNO[11]_net_1\);
    
    block15_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(3), Y => \wen_b15_1[1]\);
    
    \readData_31_bm_1_1_RNO_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[14]\, D => \readData5[14]\, Y => 
        \readData_21_1_1[13]\);
    
    \readData_31_bm_1_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[9]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[9]_net_1\, Y => 
        \readData_31_bm_1_1[9]_net_1\);
    
    block16_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(2), Y => 
        \wen_b16_1[0]\);
    
    \readData_31_bm_RNO[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[10]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[9]\, D => \readData15[10]\, Y => 
        \readData_31_bm_RNO[9]_net_1\);
    
    \readData_31_am_RNO_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[25]\, D => \readData6[25]\, Y => 
        \readData_13_1_1[23]\);
    
    block26_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(3), Y => \wen_b26_1[1]\);
    
    block26_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(0), Y => \wen_a26_1[0]\);
    
    block23_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(3), Y => \wen_b23_1[1]\);
    
    \readData_31_bm_1_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[25]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[25]_net_1\, Y => 
        \readData_31_bm_1_1[25]_net_1\);
    
    \readData_31_bm_RNO[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[20]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[18]\, D => \readData15[20]\, Y => 
        \readData_31_bm_RNO[18]_net_1\);
    
    \readData_31_am_RNO_2[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[32]\, D => \readData2[32]\, Y => 
        \readData_10_1_1[29]\);
    
    block8_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(2), Y => \wen_b8_1[0]\);
    
    \readData_31_am[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[5]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[5]_net_1\, D
         => \readData_31_am_RNO_0[5]_net_1\, Y => 
        \readData_31_am[5]_net_1\);
    
    block11_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(0), Y => \wen_a11_1[0]\);
    
    \readData_31_am_RNO_2[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[27]\, D => \readData2[27]\, Y => 
        \readData_10_1_1[24]\);
    
    \readData_31_am_1_1_RNO_2[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[21]\, D => \readData0[21]\, Y => 
        \readData_3_1_1[19]\);
    
    block10 : RAM1K18
      port map(A_DOUT(17) => nc123, A_DOUT(16) => 
        \readData10[16]\, A_DOUT(15) => \readData10[15]\, 
        A_DOUT(14) => \readData10[14]\, A_DOUT(13) => 
        \readData10[13]\, A_DOUT(12) => \readData10[12]\, 
        A_DOUT(11) => \readData10[11]\, A_DOUT(10) => 
        \readData10[10]\, A_DOUT(9) => \readData10[9]\, A_DOUT(8)
         => nc121, A_DOUT(7) => \readData10[7]\, A_DOUT(6) => 
        \readData10[6]\, A_DOUT(5) => \readData10[5]\, A_DOUT(4)
         => \readData10[4]\, A_DOUT(3) => \readData10[3]\, 
        A_DOUT(2) => \readData10[2]\, A_DOUT(1) => 
        \readData10[1]\, A_DOUT(0) => \readData10[0]\, B_DOUT(17)
         => nc47, B_DOUT(16) => \readData10[34]\, B_DOUT(15) => 
        \readData10[33]\, B_DOUT(14) => \readData10[32]\, 
        B_DOUT(13) => \readData10[31]\, B_DOUT(12) => 
        \readData10[30]\, B_DOUT(11) => \readData10[29]\, 
        B_DOUT(10) => \readData10[28]\, B_DOUT(9) => 
        \readData10[27]\, B_DOUT(8) => nc113, B_DOUT(7) => 
        \readData10[25]\, B_DOUT(6) => \readData10[24]\, 
        B_DOUT(5) => \readData10[23]\, B_DOUT(4) => 
        \readData10[22]\, B_DOUT(3) => \readData10[21]\, 
        B_DOUT(2) => \readData10[20]\, B_DOUT(1) => 
        \readData10[19]\, B_DOUT(0) => \readData10[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a10_1[1]\, 
        A_WEN(0) => \wen_a10_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b10_1[1]\, 
        B_WEN(0) => \wen_b10_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_1_1_RNO[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[11]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[10]\, D => \readData12[11]\, Y => 
        \readData_31_am_1_1_RNO[10]_net_1\);
    
    \readData_31_am_RNO_0[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[0]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[0]\, D => \readData10[0]\, Y => 
        \readData_31_am_RNO_0[0]_net_1\);
    
    block23_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(1), Y => \wen_a23_1[1]\);
    
    \readData_31_am_RNO_0[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[28]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[25]\, D => \readData10[28]\, Y => 
        \readData_31_am_RNO_0[25]_net_1\);
    
    \readData_31_am_1_1_RNO_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[21]\, D => \readData4[21]\, Y => 
        \readData_6_1_1[19]\);
    
    \readData_31_bm_1_1_RNO_2[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[21]\, D => \readData1[21]\, Y => 
        \readData_18_1_1[19]\);
    
    \readData_31_bm_1_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[19]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[19]_net_1\, Y => 
        \readData_31_bm_1_1[19]_net_1\);
    
    \readData_31_am_1_1_RNO_0[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[19]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[17]\, D => \readData8[19]\, Y => 
        \readData_31_am_1_1_RNO_0[17]_net_1\);
    
    \readData_31_bm_RNO_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[27]\, D => \readData7[27]\, Y => 
        \readData_28_1_1[24]\);
    
    \readData_31_bm_RNO[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[9]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[8]\, D => \readData15[9]\, Y => 
        \readData_31_bm_RNO[8]_net_1\);
    
    \readData_31_bm_RNO_2[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[1]\, D => \readData3[1]\, Y => 
        \readData_25_1_1[1]\);
    
    \readData_31_bm_1_1_RNO_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[21]\, D => \readData5[21]\, Y => 
        \readData_21_1_1[19]\);
    
    \readData_31_am_1_1_RNO_0[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[3]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[3]\, D => \readData8[3]\, Y => 
        \readData_31_am_1_1_RNO_0[3]_net_1\);
    
    \readData_31_bm_RNO_0[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[18]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[16]\, D => \readData11[18]\, Y => 
        \readData_31_bm_RNO_0[16]_net_1\);
    
    \readData_31_bm_1_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[11]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[11]_net_1\, Y => 
        \readData_31_bm_1_1[11]_net_1\);
    
    block21 : RAM1K18
      port map(A_DOUT(17) => nc111, A_DOUT(16) => 
        \readData21[16]\, A_DOUT(15) => \readData21[15]\, 
        A_DOUT(14) => \readData21[14]\, A_DOUT(13) => 
        \readData21[13]\, A_DOUT(12) => \readData21[12]\, 
        A_DOUT(11) => \readData21[11]\, A_DOUT(10) => 
        \readData21[10]\, A_DOUT(9) => \readData21[9]\, A_DOUT(8)
         => nc34, A_DOUT(7) => \readData21[7]\, A_DOUT(6) => 
        \readData21[6]\, A_DOUT(5) => \readData21[5]\, A_DOUT(4)
         => \readData21[4]\, A_DOUT(3) => \readData21[3]\, 
        A_DOUT(2) => \readData21[2]\, A_DOUT(1) => 
        \readData21[1]\, A_DOUT(0) => \readData21[0]\, B_DOUT(17)
         => nc98, B_DOUT(16) => \readData21[34]\, B_DOUT(15) => 
        \readData21[33]\, B_DOUT(14) => \readData21[32]\, 
        B_DOUT(13) => \readData21[31]\, B_DOUT(12) => 
        \readData21[30]\, B_DOUT(11) => \readData21[29]\, 
        B_DOUT(10) => \readData21[28]\, B_DOUT(9) => 
        \readData21[27]\, B_DOUT(8) => nc89, B_DOUT(7) => 
        \readData21[25]\, B_DOUT(6) => \readData21[24]\, 
        B_DOUT(5) => \readData21[23]\, B_DOUT(4) => 
        \readData21[22]\, B_DOUT(3) => \readData21[21]\, 
        B_DOUT(2) => \readData21[20]\, B_DOUT(1) => 
        \readData21[19]\, B_DOUT(0) => \readData21[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a21_1[1]\, 
        A_WEN(0) => \wen_a21_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b_m[1]\, 
        B_WEN(0) => \wen_b_m[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_1_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[16]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[16]_net_1\, Y => 
        \readData_31_am_1_1[16]_net_1\);
    
    \readData_31_bm_RNO_0[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[34]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[31]\, D => \readData11[34]\, Y => 
        \readData_31_bm_RNO_0[31]_net_1\);
    
    block8 : RAM1K18
      port map(A_DOUT(17) => nc70, A_DOUT(16) => \readData8[16]\, 
        A_DOUT(15) => \readData8[15]\, A_DOUT(14) => 
        \readData8[14]\, A_DOUT(13) => \readData8[13]\, 
        A_DOUT(12) => \readData8[12]\, A_DOUT(11) => 
        \readData8[11]\, A_DOUT(10) => \readData8[10]\, A_DOUT(9)
         => \readData8[9]\, A_DOUT(8) => nc60, A_DOUT(7) => 
        \readData8[7]\, A_DOUT(6) => \readData8[6]\, A_DOUT(5)
         => \readData8[5]\, A_DOUT(4) => \readData8[4]\, 
        A_DOUT(3) => \readData8[3]\, A_DOUT(2) => \readData8[2]\, 
        A_DOUT(1) => \readData8[1]\, A_DOUT(0) => \readData8[0]\, 
        B_DOUT(17) => nc105, B_DOUT(16) => \readData8[34]\, 
        B_DOUT(15) => \readData8[33]\, B_DOUT(14) => 
        \readData8[32]\, B_DOUT(13) => \readData8[31]\, 
        B_DOUT(12) => \readData8[30]\, B_DOUT(11) => 
        \readData8[29]\, B_DOUT(10) => \readData8[28]\, B_DOUT(9)
         => \readData8[27]\, B_DOUT(8) => nc74, B_DOUT(7) => 
        \readData8[25]\, B_DOUT(6) => \readData8[24]\, B_DOUT(5)
         => \readData8[23]\, B_DOUT(4) => \readData8[22]\, 
        B_DOUT(3) => \readData8[21]\, B_DOUT(2) => 
        \readData8[20]\, B_DOUT(1) => \readData8[19]\, B_DOUT(0)
         => \readData8[18]\, BUSY => OPEN, A_CLK => FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_21_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a8_1[1]\, 
        A_WEN(0) => \wen_a8_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b8_1[1]\, 
        B_WEN(0) => \wen_b8_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block12_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(2), Y => \wen_b12_1[0]\);
    
    \readData_31_bm_RNO[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[28]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[25]\, D => \readData15[28]\, Y => 
        \readData_31_bm_RNO[25]_net_1\);
    
    \readData_31_am_RNO_0[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[34]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[31]\, D => \readData10[34]\, Y => 
        \readData_31_am_RNO_0[31]_net_1\);
    
    \readData_31_bm_RNO_0[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[30]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[27]\, D => \readData11[30]\, Y => 
        \readData_31_bm_RNO_0[27]_net_1\);
    
    \readData_31_bm[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[28]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[28]_net_1\, D
         => \readData_31_bm_RNO_0[28]_net_1\, Y => 
        \readData_31_bm[28]_net_1\);
    
    \readData_31_am_RNO_2[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[16]\, D => \readData2[16]\, Y => 
        \readData_10_1_1[15]\);
    
    \readData_31_bm_RNO_0[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[21]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[19]\, D => \readData11[21]\, Y => 
        \readData_31_bm_RNO_0[19]_net_1\);
    
    \readData_31_am_1_1_RNO_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[27]\, D => \readData4[27]\, Y => 
        \readData_6_1_1[24]\);
    
    block22 : RAM1K18
      port map(A_DOUT(17) => nc120, A_DOUT(16) => 
        \readData22[16]\, A_DOUT(15) => \readData22[15]\, 
        A_DOUT(14) => \readData22[14]\, A_DOUT(13) => 
        \readData22[13]\, A_DOUT(12) => \readData22[12]\, 
        A_DOUT(11) => \readData22[11]\, A_DOUT(10) => 
        \readData22[10]\, A_DOUT(9) => \readData22[9]\, A_DOUT(8)
         => nc119, A_DOUT(7) => \readData22[7]\, A_DOUT(6) => 
        \readData22[6]\, A_DOUT(5) => \readData22[5]\, A_DOUT(4)
         => \readData22[4]\, A_DOUT(3) => \readData22[3]\, 
        A_DOUT(2) => \readData22[2]\, A_DOUT(1) => 
        \readData22[1]\, A_DOUT(0) => \readData22[0]\, B_DOUT(17)
         => nc64, B_DOUT(16) => \readData22[34]\, B_DOUT(15) => 
        \readData22[33]\, B_DOUT(14) => \readData22[32]\, 
        B_DOUT(13) => \readData22[31]\, B_DOUT(12) => 
        \readData22[30]\, B_DOUT(11) => \readData22[29]\, 
        B_DOUT(10) => \readData22[28]\, B_DOUT(9) => 
        \readData22[27]\, B_DOUT(8) => nc110, B_DOUT(7) => 
        \readData22[25]\, B_DOUT(6) => \readData22[24]\, 
        B_DOUT(5) => \readData22[23]\, B_DOUT(4) => 
        \readData22[22]\, B_DOUT(3) => \readData22[21]\, 
        B_DOUT(2) => \readData22[20]\, B_DOUT(1) => 
        \readData22[19]\, B_DOUT(0) => \readData22[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a_m[1]\, 
        A_WEN(0) => \wen_a_m[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b22_1[1]\, 
        B_WEN(0) => \wen_b22_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_ns[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[5]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[5]_net_1\, Y => 
        ram_rdata(5));
    
    \readData_31_ns[25]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[25]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[25]_net_1\, Y => 
        ram_rdata(25));
    
    \readData_31_am_RNO_0[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[6]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[6]\, D => \readData10[6]\, Y => 
        \readData_31_am_RNO_0[6]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[20]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[18]\, D => \readData9[20]\, Y => 
        \readData_31_bm_1_1_RNO_0[18]_net_1\);
    
    \readData_31_am_RNO_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[16]\, D => \readData6[16]\, Y => 
        \readData_13_1_1[15]\);
    
    \readData_31_bm[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[13]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[13]_net_1\, D
         => \readData_31_bm_RNO_0[13]_net_1\, Y => 
        \readData_31_bm[13]_net_1\);
    
    \readData_31_am_1_1_RNO[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[22]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[20]\, D => \readData12[22]\, Y => 
        \readData_31_am_1_1_RNO[20]_net_1\);
    
    \readData_31_am_1_1_RNO_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[10]\, D => \readData4[10]\, Y => 
        \readData_6_1_1[9]\);
    
    block23 : RAM1K18
      port map(A_DOUT(17) => nc9, A_DOUT(16) => \readData23[16]\, 
        A_DOUT(15) => \readData23[15]\, A_DOUT(14) => 
        \readData23[14]\, A_DOUT(13) => \readData23[13]\, 
        A_DOUT(12) => \readData23[12]\, A_DOUT(11) => 
        \readData23[11]\, A_DOUT(10) => \readData23[10]\, 
        A_DOUT(9) => \readData23[9]\, A_DOUT(8) => nc92, 
        A_DOUT(7) => \readData23[7]\, A_DOUT(6) => 
        \readData23[6]\, A_DOUT(5) => \readData23[5]\, A_DOUT(4)
         => \readData23[4]\, A_DOUT(3) => \readData23[3]\, 
        A_DOUT(2) => \readData23[2]\, A_DOUT(1) => 
        \readData23[1]\, A_DOUT(0) => \readData23[0]\, B_DOUT(17)
         => nc91, B_DOUT(16) => \readData23[34]\, B_DOUT(15) => 
        \readData23[33]\, B_DOUT(14) => \readData23[32]\, 
        B_DOUT(13) => \readData23[31]\, B_DOUT(12) => 
        \readData23[30]\, B_DOUT(11) => \readData23[29]\, 
        B_DOUT(10) => \readData23[28]\, B_DOUT(9) => 
        \readData23[27]\, B_DOUT(8) => nc13, B_DOUT(7) => 
        \readData23[25]\, B_DOUT(6) => \readData23[24]\, 
        B_DOUT(5) => \readData23[23]\, B_DOUT(4) => 
        \readData23[22]\, B_DOUT(3) => \readData23[21]\, 
        B_DOUT(2) => \readData23[20]\, B_DOUT(1) => 
        \readData23[19]\, B_DOUT(0) => \readData23[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a23_1[1]\, 
        A_WEN(0) => \wen_a23_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b23_1[1]\, 
        B_WEN(0) => \wen_b23_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[5]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[5]\, D => \readData15[5]\, Y => 
        \readData_31_bm_RNO[5]_net_1\);
    
    \readData_31_bm_RNO_0[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[2]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[2]\, D => \readData11[2]\, Y => 
        \readData_31_bm_RNO_0[2]_net_1\);
    
    \readData_31_am_1_1_RNO[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[3]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[3]\, D => \readData12[3]\, Y => 
        \readData_31_am_1_1_RNO[3]_net_1\);
    
    \readData_31_am_1_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[12]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[12]_net_1\, Y => 
        \readData_31_am_1_1[12]_net_1\);
    
    \readData_31_am[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[27]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[27]_net_1\, D
         => \readData_31_am_RNO_0[27]_net_1\, Y => 
        \readData_31_am[27]_net_1\);
    
    \readData_31_am_1_1_RNO_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[28]\, D => \readData4[28]\, Y => 
        \readData_6_1_1[25]\);
    
    \readData_31_bm_RNO_2[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[29]\, D => \readData3[29]\, Y => 
        \readData_25_1_1[26]\);
    
    block13_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(2), Y => 
        \wen_b13_1[0]\);
    
    \readData_31_am_1_1_RNO[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[10]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[9]\, D => \readData12[10]\, Y => 
        \readData_31_am_1_1_RNO[9]_net_1\);
    
    \readData_31_am_1_1_RNO_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[0]\, D => \readData4[0]\, Y => 
        \readData_6_1_1[0]\);
    
    \readData_31_am_1_1_RNO[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[14]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[13]\, D => \readData12[14]\, Y => 
        \readData_31_am_1_1_RNO[13]_net_1\);
    
    \readData_31_bm_RNO_2[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[19]\, D => \readData3[19]\, Y => 
        \readData_25_1_1[17]\);
    
    \readData_31_bm_1_1_RNO_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[4]\, D => \readData5[4]\, Y => 
        \readData_21_1_1[4]\);
    
    \readData_31_bm_RNO_0[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[24]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[22]\, D => \readData11[24]\, Y => 
        \readData_31_bm_RNO_0[22]_net_1\);
    
    \readData_31_am_RNO[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[28]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[25]\, D => \readData14[28]\, Y => 
        \readData_31_am_RNO[25]_net_1\);
    
    \readData_31_am_1_1_RNO_0[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[31]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[28]\, D => \readData8[31]\, Y => 
        \readData_31_am_1_1_RNO_0[28]_net_1\);
    
    block28 : RAM1K18
      port map(A_DOUT(17) => nc23, A_DOUT(16) => \readData28[16]\, 
        A_DOUT(15) => \readData28[15]\, A_DOUT(14) => 
        \readData28[14]\, A_DOUT(13) => \readData28[13]\, 
        A_DOUT(12) => \readData28[12]\, A_DOUT(11) => 
        \readData28[11]\, A_DOUT(10) => \readData28[10]\, 
        A_DOUT(9) => \readData28[9]\, A_DOUT(8) => nc55, 
        A_DOUT(7) => \readData28[7]\, A_DOUT(6) => 
        \readData28[6]\, A_DOUT(5) => \readData28[5]\, A_DOUT(4)
         => \readData28[4]\, A_DOUT(3) => \readData28[3]\, 
        A_DOUT(2) => \readData28[2]\, A_DOUT(1) => 
        \readData28[1]\, A_DOUT(0) => \readData28[0]\, B_DOUT(17)
         => nc80, B_DOUT(16) => \readData28[34]\, B_DOUT(15) => 
        \readData28[33]\, B_DOUT(14) => \readData28[32]\, 
        B_DOUT(13) => \readData28[31]\, B_DOUT(12) => 
        \readData28[30]\, B_DOUT(11) => \readData28[29]\, 
        B_DOUT(10) => \readData28[28]\, B_DOUT(9) => 
        \readData28[27]\, B_DOUT(8) => nc33, B_DOUT(7) => 
        \readData28[25]\, B_DOUT(6) => \readData28[24]\, 
        B_DOUT(5) => \readData28[23]\, B_DOUT(4) => 
        \readData28[22]\, B_DOUT(3) => \readData28[21]\, 
        B_DOUT(2) => \readData28[20]\, B_DOUT(1) => 
        \readData28[19]\, B_DOUT(0) => \readData28[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a28_1[1]\, 
        A_WEN(0) => \wen_a28_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b28_1[1]\, 
        B_WEN(0) => \wen_b28_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_2[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[32]\, D => \readData3[32]\, Y => 
        \readData_25_1_1[29]\);
    
    \readData_31_am[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[14]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[14]_net_1\, D
         => \readData_31_am_RNO_0[14]_net_1\, Y => 
        \readData_31_am[14]_net_1\);
    
    \readData_31_bm_RNO_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[19]\, D => \readData7[19]\, Y => 
        \readData_28_1_1[17]\);
    
    \readData_31_am_RNO_2[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[4]\, D => \readData2[4]\, Y => 
        \readData_10_1_1[4]\);
    
    \readData_31_bm_1_1_RNO_0[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[6]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[6]\, D => \readData9[6]\, Y => 
        \readData_31_bm_1_1_RNO_0[6]_net_1\);
    
    \readData_31_bm_RNO_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[34]\, D => \readData7[34]\, Y => 
        \readData_28_1_1[31]\);
    
    \readData_31_am_RNO_0[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[24]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[22]\, D => \readData10[24]\, Y => 
        \readData_31_am_RNO_0[22]_net_1\);
    
    \readData_31_bm_RNO[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[34]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[31]\, D => \readData15[34]\, Y => 
        \readData_31_bm_RNO[31]_net_1\);
    
    \readData_31_am_RNO_2[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[6]\, D => \readData2[6]\, Y => 
        \readData_10_1_1[6]\);
    
    \readData_31_am_1_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[24]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[24]_net_1\, Y => 
        \readData_31_am_1_1[24]_net_1\);
    
    \readData_31_ns[16]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[16]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[16]_net_1\, Y => 
        ram_rdata(16));
    
    \readData_31_am_RNO_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[34]\, D => \readData6[34]\, Y => 
        \readData_13_1_1[31]\);
    
    \readData_31_bm_RNO_0[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[14]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[13]\, D => \readData11[14]\, Y => 
        \readData_31_bm_RNO_0[13]_net_1\);
    
    \readData_31_bm[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[19]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[19]_net_1\, D
         => \readData_31_bm_RNO_0[19]_net_1\, Y => 
        \readData_31_bm[19]_net_1\);
    
    \readData_31_bm_RNO_0[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[11]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[10]\, D => \readData11[11]\, Y => 
        \readData_31_bm_RNO_0[10]_net_1\);
    
    \readData_31_bm_RNO_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[9]\, D => \readData7[9]\, Y => 
        \readData_28_1_1[8]\);
    
    \readData_31_am[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[12]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[12]_net_1\, D
         => \readData_31_am_RNO_0[12]_net_1\, Y => 
        \readData_31_am[12]_net_1\);
    
    \readData_31_am_1_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[19]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[19]_net_1\, Y => 
        \readData_31_am_1_1[19]_net_1\);
    
    \readData_31_bm_RNO_2[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[13]\, D => \readData3[13]\, Y => 
        \readData_25_1_1[12]\);
    
    \readData_31_bm_1_1_RNO[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[0]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[0]\, D => \readData13[0]\, Y => 
        \readData_31_bm_1_1_RNO[0]_net_1\);
    
    \readData_31_bm_1_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[22]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[22]_net_1\, Y => 
        \readData_31_bm_1_1[22]_net_1\);
    
    block24_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(2), Y => \wen_b24_1[0]\);
    
    \readData_31_bm_RNO_2[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[9]\, D => \readData3[9]\, Y => 
        \readData_25_1_1[8]\);
    
    \readData_31_am_1_1_RNO_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[9]\, D => \readData4[9]\, Y => 
        \readData_6_1_1[8]\);
    
    \readData_31_bm_RNO[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[14]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[13]\, D => \readData15[14]\, Y => 
        \readData_31_bm_RNO[13]_net_1\);
    
    \readData_31_bm_RNO_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[13]\, D => \readData7[13]\, Y => 
        \readData_28_1_1[12]\);
    
    \readData_31_bm_RNO[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[33]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[30]\, D => \readData15[33]\, Y => 
        \readData_31_bm_RNO[30]_net_1\);
    
    \readData_31_bm[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[12]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[12]_net_1\, D
         => \readData_31_bm_RNO_0[12]_net_1\, Y => 
        \readData_31_bm[12]_net_1\);
    
    \readData_31_am_RNO_2[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[13]\, D => \readData2[13]\, Y => 
        \readData_10_1_1[12]\);
    
    \readData_31_am_1_1_RNO[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[25]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[23]\, D => \readData12[25]\, Y => 
        \readData_31_am_1_1_RNO[23]_net_1\);
    
    \readData_31_am_RNO_0[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[1]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[1]\, D => \readData10[1]\, Y => 
        \readData_31_am_RNO_0[1]_net_1\);
    
    block17 : RAM1K18
      port map(A_DOUT(17) => nc84, A_DOUT(16) => \readData17[16]\, 
        A_DOUT(15) => \readData17[15]\, A_DOUT(14) => 
        \readData17[14]\, A_DOUT(13) => \readData17[13]\, 
        A_DOUT(12) => \readData17[12]\, A_DOUT(11) => 
        \readData17[11]\, A_DOUT(10) => \readData17[10]\, 
        A_DOUT(9) => \readData17[9]\, A_DOUT(8) => nc16, 
        A_DOUT(7) => \readData17[7]\, A_DOUT(6) => 
        \readData17[6]\, A_DOUT(5) => \readData17[5]\, A_DOUT(4)
         => \readData17[4]\, A_DOUT(3) => \readData17[3]\, 
        A_DOUT(2) => \readData17[2]\, A_DOUT(1) => 
        \readData17[1]\, A_DOUT(0) => \readData17[0]\, B_DOUT(17)
         => nc26, B_DOUT(16) => \readData17[34]\, B_DOUT(15) => 
        \readData17[33]\, B_DOUT(14) => \readData17[32]\, 
        B_DOUT(13) => \readData17[31]\, B_DOUT(12) => 
        \readData17[30]\, B_DOUT(11) => \readData17[29]\, 
        B_DOUT(10) => \readData17[28]\, B_DOUT(9) => 
        \readData17[27]\, B_DOUT(8) => nc45, B_DOUT(7) => 
        \readData17[25]\, B_DOUT(6) => \readData17[24]\, 
        B_DOUT(5) => \readData17[23]\, B_DOUT(4) => 
        \readData17[22]\, B_DOUT(3) => \readData17[21]\, 
        B_DOUT(2) => \readData17[20]\, B_DOUT(1) => 
        \readData17[19]\, B_DOUT(0) => \readData17[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a17_1[1]\, 
        A_WEN(0) => \wen_a17_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b17_1[1]\, 
        B_WEN(0) => \wen_b17_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \readData_31_am_1_1_RNO_2[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[31]\, D => \readData0[31]\, Y => 
        \readData_3_1_1[28]\);
    
    \readData_31_bm_1_1_RNO_2[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[9]\, D => \readData1[9]\, Y => 
        \readData_18_1_1[8]\);
    
    \readData_31_am_RNO_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[13]\, D => \readData6[13]\, Y => 
        \readData_13_1_1[12]\);
    
    \readData_31_bm_RNO_2[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[25]\, D => \readData3[25]\, Y => 
        \readData_25_1_1[23]\);
    
    block21_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(2), Y => \wen_b_m[0]\);
    
    block30_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(1), Y => \wen_a30_1[1]\);
    
    \readData_31_ns[31]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[31]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[31]_net_1\, Y => 
        ram_rdata(31));
    
    \readData_31_am_1_1_RNO_0[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[4]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[4]\, D => \readData8[4]\, Y => 
        \readData_31_am_1_1_RNO_0[4]_net_1\);
    
    \readData_31_bm_RNO_2[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[22]\, D => \readData3[22]\, Y => 
        \readData_25_1_1[20]\);
    
    \readData_31_am_1_1_RNO_2[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[19]\, D => \readData0[19]\, Y => 
        \readData_3_1_1[17]\);
    
    block21_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(0), Y => \wen_a21_1[0]\);
    
    \readData_31_bm_1_1_RNO_0[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[16]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[15]\, D => \readData9[16]\, Y => 
        \readData_31_bm_1_1_RNO_0[15]_net_1\);
    
    \readData_31_am_1_1_RNO_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[19]\, D => \readData4[19]\, Y => 
        \readData_6_1_1[17]\);
    
    \readData_31_am_1_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[7]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[7]_net_1\, Y => 
        \readData_31_am_1_1[7]_net_1\);
    
    block7_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(1), Y => \wen_a7_1[1]\);
    
    \readData_31_bm_RNO_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[28]\, D => \readData7[28]\, Y => 
        \readData_28_1_1[25]\);
    
    block22_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(3), Y => \wen_b22_1[1]\);
    
    \readData_31_bm_1_1_RNO_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[1]\, D => \readData5[1]\, Y => 
        \readData_21_1_1[1]\);
    
    \readData_31_bm[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[5]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[5]_net_1\, D
         => \readData_31_bm_RNO_0[5]_net_1\, Y => 
        \readData_31_bm[5]_net_1\);
    
    block6_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(2), Y => \wen_b6_1[0]\);
    
    \readData_31_bm[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[27]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[27]_net_1\, D
         => \readData_31_bm_RNO_0[27]_net_1\, Y => 
        \readData_31_bm[27]_net_1\);
    
    \readData_31_am_1_1_RNO_0[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[25]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[23]\, D => \readData8[25]\, Y => 
        \readData_31_am_1_1_RNO_0[23]_net_1\);
    
    \readData_31_bm_1_1_RNO[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[14]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[13]\, D => \readData13[14]\, Y => 
        \readData_31_bm_1_1_RNO[13]_net_1\);
    
    block9_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(2), Y => \wen_b9_1[0]\);
    
    \readData_31_am_1_1_RNO_0[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[9]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[8]\, D => \readData8[9]\, Y => 
        \readData_31_am_1_1_RNO_0[8]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[5]\, D => \readData1[5]\, Y => 
        \readData_18_1_1[5]\);
    
    block24_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(3), Y => \wen_b24_1[1]\);
    
    \readData_31_bm_1_1_RNO_2[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[20]\, D => \readData1[20]\, Y => 
        \readData_18_1_1[18]\);
    
    \readData_31_bm_1_1_RNO[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[21]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[19]\, D => \readData13[21]\, Y => 
        \readData_31_bm_1_1_RNO[19]_net_1\);
    
    \readData_31_am_1_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[0]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[0]_net_1\, Y => 
        \readData_31_am_1_1[0]_net_1\);
    
    \readData_31_am_1_1_RNO[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[18]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[16]\, D => \readData12[18]\, Y => 
        \readData_31_am_1_1_RNO[16]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[20]\, D => \readData5[20]\, Y => 
        \readData_21_1_1[18]\);
    
    \readData_31_am_RNO_2[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[5]\, D => \readData2[5]\, Y => 
        \readData_10_1_1[5]\);
    
    block16_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(1), Y => 
        \wen_a16_1[1]\);
    
    \readData_31_am_RNO[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[10]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[9]\, D => \readData14[10]\, Y => 
        \readData_31_am_RNO[9]_net_1\);
    
    \readData_31_bm_1_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[28]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[28]_net_1\, Y => 
        \readData_31_bm_1_1[28]_net_1\);
    
    \readData_31_am_1_1_RNO_2[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[4]\, D => \readData0[4]\, Y => 
        \readData_3_1_1[4]\);
    
    \readData_31_am_RNO[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[13]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[12]\, D => \readData14[13]\, Y => 
        \readData_31_am_RNO[12]_net_1\);
    
    \readData_31_am_1_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[15]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[15]_net_1\, Y => 
        \readData_31_am_1_1[15]_net_1\);
    
    \readData_31_bm_RNO[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[13]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[12]\, D => \readData15[13]\, Y => 
        \readData_31_bm_RNO[12]_net_1\);
    
    \readData_31_am_RNO_0[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[4]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[4]\, D => \readData10[4]\, Y => 
        \readData_31_am_RNO_0[4]_net_1\);
    
    block31 : RAM1K18
      port map(A_DOUT(17) => nc73, A_DOUT(16) => \readData31[16]\, 
        A_DOUT(15) => \readData31[15]\, A_DOUT(14) => 
        \readData31[14]\, A_DOUT(13) => \readData31[13]\, 
        A_DOUT(12) => \readData31[12]\, A_DOUT(11) => 
        \readData31[11]\, A_DOUT(10) => \readData31[10]\, 
        A_DOUT(9) => \readData31[9]\, A_DOUT(8) => nc58, 
        A_DOUT(7) => \readData31[7]\, A_DOUT(6) => 
        \readData31[6]\, A_DOUT(5) => \readData31[5]\, A_DOUT(4)
         => \readData31[4]\, A_DOUT(3) => \readData31[3]\, 
        A_DOUT(2) => \readData31[2]\, A_DOUT(1) => 
        \readData31[1]\, A_DOUT(0) => \readData31[0]\, B_DOUT(17)
         => nc63, B_DOUT(16) => \readData31[34]\, B_DOUT(15) => 
        \readData31[33]\, B_DOUT(14) => \readData31[32]\, 
        B_DOUT(13) => \readData31[31]\, B_DOUT(12) => 
        \readData31[30]\, B_DOUT(11) => \readData31[29]\, 
        B_DOUT(10) => \readData31[28]\, B_DOUT(9) => 
        \readData31[27]\, B_DOUT(8) => nc27, B_DOUT(7) => 
        \readData31[25]\, B_DOUT(6) => \readData31[24]\, 
        B_DOUT(5) => \readData31[23]\, B_DOUT(4) => 
        \readData31[22]\, B_DOUT(3) => \readData31[21]\, 
        B_DOUT(2) => \readData31[20]\, B_DOUT(1) => 
        \readData31[19]\, B_DOUT(0) => \readData31[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a31_1[1]\, 
        A_WEN(0) => \wen_a31_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b31_1[1]\, 
        B_WEN(0) => \wen_b31_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[25]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[25]_net_1\, D
         => \readData_31_bm_RNO_0[25]_net_1\, Y => 
        \readData_31_bm[25]_net_1\);
    
    \readData_31_am_RNO_0[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[33]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[30]\, D => \readData10[33]\, Y => 
        \readData_31_am_RNO_0[30]_net_1\);
    
    block13_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(0), Y => 
        \wen_a13_1[0]\);
    
    \readData_31_am_1_1_RNO_2[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[1]\, D => \readData0[1]\, Y => 
        \readData_3_1_1[1]\);
    
    block14_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(1), Y => \wen_a14_1[1]\);
    
    \readData_31_am_1_1_RNO_0[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[10]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[9]\, D => \readData8[10]\, Y => 
        \readData_31_am_1_1_RNO_0[9]_net_1\);
    
    \readData_31_am_1_1_RNO_2[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[25]\, D => \readData0[25]\, Y => 
        \readData_3_1_1[23]\);
    
    \readData_31_ns[28]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[28]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[28]_net_1\, Y => 
        ram_rdata(28));
    
    \readData_31_bm_1_1_RNO[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[25]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[23]\, D => \readData13[25]\, Y => 
        \readData_31_bm_1_1_RNO[23]_net_1\);
    
    block26 : RAM1K18
      port map(A_DOUT(17) => nc17, A_DOUT(16) => \readData26[16]\, 
        A_DOUT(15) => \readData26[15]\, A_DOUT(14) => 
        \readData26[14]\, A_DOUT(13) => \readData26[13]\, 
        A_DOUT(12) => \readData26[12]\, A_DOUT(11) => 
        \readData26[11]\, A_DOUT(10) => \readData26[10]\, 
        A_DOUT(9) => \readData26[9]\, A_DOUT(8) => nc127, 
        A_DOUT(7) => \readData26[7]\, A_DOUT(6) => 
        \readData26[6]\, A_DOUT(5) => \readData26[5]\, A_DOUT(4)
         => \readData26[4]\, A_DOUT(3) => \readData26[3]\, 
        A_DOUT(2) => \readData26[2]\, A_DOUT(1) => 
        \readData26[1]\, A_DOUT(0) => \readData26[0]\, B_DOUT(17)
         => nc99, B_DOUT(16) => \readData26[34]\, B_DOUT(15) => 
        \readData26[33]\, B_DOUT(14) => \readData26[32]\, 
        B_DOUT(13) => \readData26[31]\, B_DOUT(12) => 
        \readData26[30]\, B_DOUT(11) => \readData26[29]\, 
        B_DOUT(10) => \readData26[28]\, B_DOUT(9) => 
        \readData26[27]\, B_DOUT(8) => nc126, B_DOUT(7) => 
        \readData26[25]\, B_DOUT(6) => \readData26[24]\, 
        B_DOUT(5) => \readData26[23]\, B_DOUT(4) => 
        \readData26[22]\, B_DOUT(3) => \readData26[21]\, 
        B_DOUT(2) => \readData26[20]\, B_DOUT(1) => 
        \readData26[19]\, B_DOUT(0) => \readData26[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a26_1[1]\, 
        A_WEN(0) => \wen_a26_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b26_1[1]\, 
        B_WEN(0) => \wen_b26_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_1_1_RNO_0[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[12]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[11]\, D => \readData8[12]\, Y => 
        \readData_31_am_1_1_RNO_0[11]_net_1\);
    
    \readData_31_ns[29]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[29]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[29]_net_1\, Y => 
        ram_rdata(29));
    
    block10_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(1), Y => \wen_a10_1[1]\);
    
    \readData_31_bm_RNO[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[1]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[1]\, D => \readData15[1]\, Y => 
        \readData_31_bm_RNO[1]_net_1\);
    
    \readData_31_bm_RNO[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[4]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[4]\, D => \readData15[4]\, Y => 
        \readData_31_bm_RNO[4]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[11]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[10]\, D => \readData9[11]\, Y => 
        \readData_31_bm_1_1_RNO_0[10]_net_1\);
    
    \readData_31_bm_1_1_RNO[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[32]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[29]\, D => \readData13[32]\, Y => 
        \readData_31_bm_1_1_RNO[29]_net_1\);
    
    \readData_31_am_RNO[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[9]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[8]\, D => \readData14[9]\, Y => 
        \readData_31_am_RNO[8]_net_1\);
    
    \readData_31_bm_RNO[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[32]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[29]\, D => \readData15[32]\, Y => 
        \readData_31_bm_RNO[29]_net_1\);
    
    \readData_31_am_1_1_RNO_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[31]\, D => \readData4[31]\, Y => 
        \readData_6_1_1[28]\);
    
    \readData_31_am_1_1_RNO_0[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[1]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[1]\, D => \readData8[1]\, Y => 
        \readData_31_am_1_1_RNO_0[1]_net_1\);
    
    \readData_31_bm_RNO_0[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[5]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[5]\, D => \readData11[5]\, Y => 
        \readData_31_bm_RNO_0[5]_net_1\);
    
    \readData_31_am_1_1_RNO[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[29]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[26]\, D => \readData12[29]\, Y => 
        \readData_31_am_1_1_RNO[26]_net_1\);
    
    \readData_31_am_1_1_RNO_0[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[33]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[30]\, D => \readData8[33]\, Y => 
        \readData_31_am_1_1_RNO_0[30]_net_1\);
    
    \readData_31_bm[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[14]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[14]_net_1\, D
         => \readData_31_bm_RNO_0[14]_net_1\, Y => 
        \readData_31_bm[14]_net_1\);
    
    \readData_31_am_1_1_RNO[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[19]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[17]\, D => \readData12[19]\, Y => 
        \readData_31_am_1_1_RNO[17]_net_1\);
    
    \readData_31_am[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[30]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[30]_net_1\, D
         => \readData_31_am_RNO_0[30]_net_1\, Y => 
        \readData_31_am[30]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[12]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[11]\, D => \readData9[12]\, Y => 
        \readData_31_bm_1_1_RNO_0[11]_net_1\);
    
    \readData_31_bm_RNO[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[3]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[3]\, D => \readData15[3]\, Y => 
        \readData_31_bm_RNO[3]_net_1\);
    
    \readData_31_am[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[11]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[11]_net_1\, D
         => \readData_31_am_RNO_0[11]_net_1\, Y => 
        \readData_31_am[11]_net_1\);
    
    block4_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(3), Y => \wen_b4_1[1]\);
    
    \readData_31_bm_1_1_RNO_0[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[19]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[17]\, D => \readData9[19]\, Y => 
        \readData_31_bm_1_1_RNO_0[17]_net_1\);
    
    \readData_31_am[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[13]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[13]_net_1\, D
         => \readData_31_am_RNO_0[13]_net_1\, Y => 
        \readData_31_am[13]_net_1\);
    
    \readData_31_bm_RNO_0[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[23]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[21]\, D => \readData11[23]\, Y => 
        \readData_31_bm_RNO_0[21]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[3]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[3]\, D => \readData9[3]\, Y => 
        \readData_31_bm_1_1_RNO_0[3]_net_1\);
    
    \readData_31_bm[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[16]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[16]_net_1\, D
         => \readData_31_bm_RNO_0[16]_net_1\, Y => 
        \readData_31_bm[16]_net_1\);
    
    \readData_31_am_RNO_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[33]\, D => \readData6[33]\, Y => 
        \readData_13_1_1[30]\);
    
    \readData_31_bm[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[31]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[31]_net_1\, D
         => \readData_31_bm_RNO_0[31]_net_1\, Y => 
        \readData_31_bm[31]_net_1\);
    
    \readData_31_am_RNO[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[5]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[5]\, D => \readData14[5]\, Y => 
        \readData_31_am_RNO[5]_net_1\);
    
    block31_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(1), Y => \wen_a31_1[1]\);
    
    \readData_31_am_RNO_0[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[23]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[21]\, D => \readData10[23]\, Y => 
        \readData_31_am_RNO_0[21]_net_1\);
    
    \readData_31_am_1_1_RNO_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[3]\, D => \readData4[3]\, Y => 
        \readData_6_1_1[3]\);
    
    readdata_xhdl1401_1_0 : CFG3
      generic map(INIT => x"40")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => ahbsram_addr(12), Y => readdata_xhdl1401_1);
    
    block6_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(3), Y => \wen_b6_1[1]\);
    
    block9_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(1), Y => \wen_a9_1[1]\);
    
    block18_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(14), C
         => readdata_xhdl1401_1, D => sram_wen_mem(1), Y => 
        \wen_a18_1[1]\);
    
    \readData_31_bm_1_1_RNO_2[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[16]\, D => \readData1[16]\, Y => 
        \readData_18_1_1[15]\);
    
    \readData_31_am[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[1]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[1]_net_1\, D
         => \readData_31_am_RNO_0[1]_net_1\, Y => 
        \readData_31_am[1]_net_1\);
    
    \readData_31_am_1_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[5]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[5]_net_1\, Y => 
        \readData_31_am_1_1[5]_net_1\);
    
    \readData_31_am[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[6]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[6]_net_1\, D
         => \readData_31_am_RNO_0[6]_net_1\, Y => 
        \readData_31_am[6]_net_1\);
    
    block8_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(1), Y => \wen_a8_1[1]\);
    
    \readData_31_ns[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[6]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[6]_net_1\, Y => 
        ram_rdata(6));
    
    \readData_31_bm_RNO_2[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[2]\, D => \readData3[2]\, Y => 
        \readData_25_1_1[2]\);
    
    \readData_31_bm_1_1_RNO_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[16]\, D => \readData5[16]\, Y => 
        \readData_21_1_1[15]\);
    
    \readData_31_bm_RNO_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[10]\, D => \readData7[10]\, Y => 
        \readData_28_1_1[9]\);
    
    \readData_31_am_1_1_RNO[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[30]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[27]\, D => \readData12[30]\, Y => 
        \readData_31_am_1_1_RNO[27]_net_1\);
    
    \readData_31_am[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[3]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[3]_net_1\, D
         => \readData_31_am_RNO_0[3]_net_1\, Y => 
        \readData_31_am[3]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[10]\, D => \readData5[10]\, Y => 
        \readData_21_1_1[9]\);
    
    \readData_31_bm_RNO_2[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[12]\, D => \readData3[12]\, Y => 
        \readData_25_1_1[11]\);
    
    \readData_31_bm_RNO_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[31]\, D => \readData7[31]\, Y => 
        \readData_28_1_1[28]\);
    
    block15_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(1), Y => \wen_a15_1[1]\);
    
    block5 : RAM1K18
      port map(A_DOUT(17) => nc117, A_DOUT(16) => \readData5[16]\, 
        A_DOUT(15) => \readData5[15]\, A_DOUT(14) => 
        \readData5[14]\, A_DOUT(13) => \readData5[13]\, 
        A_DOUT(12) => \readData5[12]\, A_DOUT(11) => 
        \readData5[11]\, A_DOUT(10) => \readData5[10]\, A_DOUT(9)
         => \readData5[9]\, A_DOUT(8) => nc36, A_DOUT(7) => 
        \readData5[7]\, A_DOUT(6) => \readData5[6]\, A_DOUT(5)
         => \readData5[5]\, A_DOUT(4) => \readData5[4]\, 
        A_DOUT(3) => \readData5[3]\, A_DOUT(2) => \readData5[2]\, 
        A_DOUT(1) => \readData5[1]\, A_DOUT(0) => \readData5[0]\, 
        B_DOUT(17) => nc116, B_DOUT(16) => \readData5[34]\, 
        B_DOUT(15) => \readData5[33]\, B_DOUT(14) => 
        \readData5[32]\, B_DOUT(13) => \readData5[31]\, 
        B_DOUT(12) => \readData5[30]\, B_DOUT(11) => 
        \readData5[29]\, B_DOUT(10) => \readData5[28]\, B_DOUT(9)
         => \readData5[27]\, B_DOUT(8) => nc48, B_DOUT(7) => 
        \readData5[25]\, B_DOUT(6) => \readData5[24]\, B_DOUT(5)
         => \readData5[23]\, B_DOUT(4) => \readData5[22]\, 
        B_DOUT(3) => \readData5[21]\, B_DOUT(2) => 
        \readData5[20]\, B_DOUT(1) => \readData5[19]\, B_DOUT(0)
         => \readData5[18]\, BUSY => OPEN, A_CLK => FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_21_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a5_1[1]\, 
        A_WEN(0) => \wen_a5_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b5_1[1]\, 
        B_WEN(0) => \wen_b5_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block31_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(3), Y => \wen_b31_1[1]\);
    
    \readData_31_am_RNO_0[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[30]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[27]\, D => \readData10[30]\, Y => 
        \readData_31_am_RNO_0[27]_net_1\);
    
    readdata_xhdl1418_0_a2_0_0 : CFG3
      generic map(INIT => x"01")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => readdata_xhdl1419_0_a2_0);
    
    \readData_31_am_RNO_2[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[12]\, D => \readData2[12]\, Y => 
        \readData_10_1_1[11]\);
    
    \readData_31_ns[12]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[12]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[12]_net_1\, Y => 
        ram_rdata(12));
    
    \readData_31_bm_RNO_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[12]\, D => \readData7[12]\, Y => 
        \readData_28_1_1[11]\);
    
    \readData_31_bm_1_1_RNO[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[18]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[16]\, D => \readData13[18]\, Y => 
        \readData_31_bm_1_1_RNO[16]_net_1\);
    
    \readData_31_am_RNO_0[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[16]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[15]\, D => \readData10[16]\, Y => 
        \readData_31_am_RNO_0[15]_net_1\);
    
    block25_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(2), Y => \wen_b25_1[0]\);
    
    \readData_31_bm_RNO_0[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[10]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[9]\, D => \readData11[10]\, Y => 
        \readData_31_bm_RNO_0[9]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[0]\, D => \readData5[0]\, Y => 
        \readData_21_1_1[0]\);
    
    \readData_31_am_RNO_0[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[31]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[28]\, D => \readData10[31]\, Y => 
        \readData_31_am_RNO_0[28]_net_1\);
    
    \readData_31_bm_1_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[29]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[29]_net_1\, Y => 
        \readData_31_bm_1_1[29]_net_1\);
    
    \readData_31_am_RNO_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[12]\, D => \readData6[12]\, Y => 
        \readData_13_1_1[11]\);
    
    \readData_31_bm_RNO_0[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[3]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[3]\, D => \readData11[3]\, Y => 
        \readData_31_bm_RNO_0[3]_net_1\);
    
    \readData_31_am_1_1_RNO_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[25]\, D => \readData4[25]\, Y => 
        \readData_6_1_1[23]\);
    
    \readData_31_am_RNO_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[1]\, D => \readData6[1]\, Y => 
        \readData_13_1_1[1]\);
    
    \readData_31_bm_1_1_RNO_0[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[25]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[23]\, D => \readData9[25]\, Y => 
        \readData_31_bm_1_1_RNO_0[23]_net_1\);
    
    \readData_31_bm_1_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[21]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[21]_net_1\, Y => 
        \readData_31_bm_1_1[21]_net_1\);
    
    \readData_31_am_1_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[26]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[26]_net_1\, Y => 
        \readData_31_am_1_1[26]_net_1\);
    
    \readData_31_ns[21]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[21]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[21]_net_1\, Y => 
        ram_rdata(21));
    
    \readData_31_am_1_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[18]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[18]_net_1\, Y => 
        \readData_31_am_1_1[18]_net_1\);
    
    block29_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(3), Y => \wen_b29_1[1]\);
    
    \readData_31_am_RNO_2[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[19]\, D => \readData2[19]\, Y => 
        \readData_10_1_1[17]\);
    
    \readData_31_bm_1_1_RNO[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[7]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[7]\, D => \readData13[7]\, Y => 
        \readData_31_bm_1_1_RNO[7]_net_1\);
    
    block1_RNO_2 : CFG4
      generic map(INIT => x"0080")

      port map(A => readdata_xhdl1419_0_a2_0, B => 
        sram_wen_mem(3), C => ahbsram_addr(11), D => 
        ahbsram_addr(15), Y => \wen_b1_1[1]\);
    
    \readData_31_am_1_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[6]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[6]_net_1\, Y => 
        \readData_31_am_1_1[6]_net_1\);
    
    \readData_31_bm_RNO_0[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[19]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[17]\, D => \readData11[19]\, Y => 
        \readData_31_bm_RNO_0[17]_net_1\);
    
    \readData_31_am_RNO[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[14]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[13]\, D => \readData14[14]\, Y => 
        \readData_31_am_RNO[13]_net_1\);
    
    \readData_31_am_RNO_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[19]\, D => \readData6[19]\, Y => 
        \readData_13_1_1[17]\);
    
    \readData_31_am_RNO_2[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[20]\, D => \readData2[20]\, Y => 
        \readData_10_1_1[18]\);
    
    \readData_31_am_1_1_RNO_2[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[12]\, D => \readData0[12]\, Y => 
        \readData_3_1_1[11]\);
    
    \readData_31_am_RNO_2[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[28]\, D => \readData2[28]\, Y => 
        \readData_10_1_1[25]\);
    
    block11_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(1), Y => \wen_a11_1[1]\);
    
    \readData_31_bm_1_1_RNO_2[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[11]\, D => \readData1[11]\, Y => 
        \readData_18_1_1[10]\);
    
    \readData_31_bm_RNO_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[7]\, D => \readData7[7]\, Y => 
        \readData_28_1_1[7]\);
    
    \readData_31_am_1_1_RNO_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[12]\, D => \readData4[12]\, Y => 
        \readData_6_1_1[11]\);
    
    \readData_31_am_1_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[22]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[22]_net_1\, Y => 
        \readData_31_am_1_1[22]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[9]\, D => \readData5[9]\, Y => 
        \readData_21_1_1[8]\);
    
    \readData_31_bm_1_1_RNO[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[29]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[26]\, D => \readData13[29]\, Y => 
        \readData_31_bm_1_1_RNO[26]_net_1\);
    
    block7_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(0), Y => \wen_a7_1[0]\);
    
    \readData_31_am_RNO_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[20]\, D => \readData6[20]\, Y => 
        \readData_13_1_1[18]\);
    
    \readData_31_am_1_1_RNO_0[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[32]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[29]\, D => \readData8[32]\, Y => 
        \readData_31_am_1_1_RNO_0[29]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[11]\, D => \readData5[11]\, Y => 
        \readData_21_1_1[10]\);
    
    \readData_31_bm[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[18]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[18]_net_1\, D
         => \readData_31_bm_RNO_0[18]_net_1\, Y => 
        \readData_31_bm[18]_net_1\);
    
    \readData_31_bm_RNO[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[27]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[24]\, D => \readData15[27]\, Y => 
        \readData_31_bm_RNO[24]_net_1\);
    
    \readData_31_am_RNO_2[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[10]\, D => \readData2[10]\, Y => 
        \readData_10_1_1[9]\);
    
    \readData_31_bm_1_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[31]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[31]_net_1\, Y => 
        \readData_31_bm_1_1[31]_net_1\);
    
    block23_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(0), Y => \wen_a23_1[0]\);
    
    \readData_31_am_1_1_RNO[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[0]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[0]\, D => \readData12[0]\, Y => 
        \readData_31_am_1_1_RNO[0]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[32]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[29]\, D => \readData9[32]\, Y => 
        \readData_31_bm_1_1_RNO_0[29]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[25]\, D => \readData1[25]\, Y => 
        \readData_18_1_1[23]\);
    
    \readData_31_am[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[17]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[17]_net_1\, D
         => \readData_31_am_RNO_0[17]_net_1\, Y => 
        \readData_31_am[17]_net_1\);
    
    \readData_31_bm_RNO_0[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[13]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[12]\, D => \readData11[13]\, Y => 
        \readData_31_bm_RNO_0[12]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[12]\, D => \readData1[12]\, Y => 
        \readData_18_1_1[11]\);
    
    \readData_31_bm_1_1_RNO_0[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[4]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[4]\, D => \readData9[4]\, Y => 
        \readData_31_bm_1_1_RNO_0[4]_net_1\);
    
    block15_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(0), Y => \wen_a15_1[0]\);
    
    block12_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(0), Y => \wen_a12_1[0]\);
    
    \readData_31_bm_RNO_2[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[30]\, D => \readData3[30]\, Y => 
        \readData_25_1_1[27]\);
    
    \readData_31_am_RNO[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[31]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[28]\, D => \readData14[31]\, Y => 
        \readData_31_am_RNO[28]_net_1\);
    
    block11_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(3), Y => \wen_b11_1[1]\);
    
    \readData_31_bm_1_1_RNO_2[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[19]\, D => \readData1[19]\, Y => 
        \readData_18_1_1[17]\);
    
    block20_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(2), Y => \wen_b20_1[0]\);
    
    \readData_31_bm_1_1_RNO_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[12]\, D => \readData5[12]\, Y => 
        \readData_21_1_1[11]\);
    
    \readData_31_am_RNO_0[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[13]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[12]\, D => \readData10[13]\, Y => 
        \readData_31_am_RNO_0[12]_net_1\);
    
    \readData_31_ns[15]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[15]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[15]_net_1\, Y => 
        ram_rdata(15));
    
    \readData_31_bm[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[20]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[20]_net_1\, D
         => \readData_31_bm_RNO_0[20]_net_1\, Y => 
        \readData_31_bm[20]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[19]\, D => \readData5[19]\, Y => 
        \readData_21_1_1[17]\);
    
    \readData_31_am_RNO[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[33]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[30]\, D => \readData14[33]\, Y => 
        \readData_31_am_RNO[30]_net_1\);
    
    \readData_31_am_RNO_2[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[3]\, D => \readData2[3]\, Y => 
        \readData_10_1_1[3]\);
    
    \readData_31_bm_RNO_0[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[0]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[0]\, D => \readData11[0]\, Y => 
        \readData_31_bm_RNO_0[0]_net_1\);
    
    \readData_31_am_RNO[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[15]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[14]\, D => \readData14[15]\, Y => 
        \readData_31_am_RNO[14]_net_1\);
    
    \readData_31_am_1_1_RNO_2[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[3]\, D => \readData0[3]\, Y => 
        \readData_3_1_1[3]\);
    
    \readData_31_am[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[4]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[4]_net_1\, D
         => \readData_31_am_RNO_0[4]_net_1\, Y => 
        \readData_31_am[4]_net_1\);
    
    block30_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(0), Y => \wen_a30_1[0]\);
    
    \readData_31_am_1_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[29]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[29]_net_1\, Y => 
        \readData_31_am_1_1[29]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[18]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[16]\, D => \readData9[18]\, Y => 
        \readData_31_bm_1_1_RNO_0[16]_net_1\);
    
    block20 : RAM1K18
      port map(A_DOUT(17) => nc37, A_DOUT(16) => \readData20[16]\, 
        A_DOUT(15) => \readData20[15]\, A_DOUT(14) => 
        \readData20[14]\, A_DOUT(13) => \readData20[13]\, 
        A_DOUT(12) => \readData20[12]\, A_DOUT(11) => 
        \readData20[11]\, A_DOUT(10) => \readData20[10]\, 
        A_DOUT(9) => \readData20[9]\, A_DOUT(8) => nc5, A_DOUT(7)
         => \readData20[7]\, A_DOUT(6) => \readData20[6]\, 
        A_DOUT(5) => \readData20[5]\, A_DOUT(4) => 
        \readData20[4]\, A_DOUT(3) => \readData20[3]\, A_DOUT(2)
         => \readData20[2]\, A_DOUT(1) => \readData20[1]\, 
        A_DOUT(0) => \readData20[0]\, B_DOUT(17) => nc103, 
        B_DOUT(16) => \readData20[34]\, B_DOUT(15) => 
        \readData20[33]\, B_DOUT(14) => \readData20[32]\, 
        B_DOUT(13) => \readData20[31]\, B_DOUT(12) => 
        \readData20[30]\, B_DOUT(11) => \readData20[29]\, 
        B_DOUT(10) => \readData20[28]\, B_DOUT(9) => 
        \readData20[27]\, B_DOUT(8) => nc101, B_DOUT(7) => 
        \readData20[25]\, B_DOUT(6) => \readData20[24]\, 
        B_DOUT(5) => \readData20[23]\, B_DOUT(4) => 
        \readData20[22]\, B_DOUT(3) => \readData20[21]\, 
        B_DOUT(2) => \readData20[20]\, B_DOUT(1) => 
        \readData20[19]\, B_DOUT(0) => \readData20[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a20_1[1]\, 
        A_WEN(0) => \wen_a20_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b20_1[1]\, 
        B_WEN(0) => \wen_b20_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_1_1_RNO_2[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[32]\, D => \readData0[32]\, Y => 
        \readData_3_1_1[29]\);
    
    \readData_31_bm_1_1_RNO_0[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[9]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[8]\, D => \readData9[9]\, Y => 
        \readData_31_bm_1_1_RNO_0[8]_net_1\);
    
    \readData_31_bm_RNO_2[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[24]\, D => \readData3[24]\, Y => 
        \readData_25_1_1[22]\);
    
    \readData_31_bm_1_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[8]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[8]_net_1\, Y => 
        \readData_31_bm_1_1[8]_net_1\);
    
    \readData_31_bm_1_1_RNO[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[16]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[15]\, D => \readData13[16]\, Y => 
        \readData_31_bm_1_1_RNO[15]_net_1\);
    
    \readData_31_bm_1_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[10]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[10]_net_1\, Y => 
        \readData_31_bm_1_1[10]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[32]\, D => \readData1[32]\, Y => 
        \readData_18_1_1[29]\);
    
    \readData_31_am_1_1_RNO_2[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[10]\, D => \readData0[10]\, Y => 
        \readData_3_1_1[9]\);
    
    \readData_31_am_RNO[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[19]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[17]\, D => \readData14[19]\, Y => 
        \readData_31_am_RNO[17]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[4]\, D => \readData1[4]\, Y => 
        \readData_18_1_1[4]\);
    
    \readData_31_am_RNO_2[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[7]\, D => \readData2[7]\, Y => 
        \readData_10_1_1[7]\);
    
    \readData_31_am_RNO_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[29]\, D => \readData6[29]\, Y => 
        \readData_13_1_1[26]\);
    
    \readData_31_am_RNO_2[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[24]\, D => \readData2[24]\, Y => 
        \readData_10_1_1[22]\);
    
    \readData_31_am_1_1_RNO_0[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[13]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[12]\, D => \readData8[13]\, Y => 
        \readData_31_am_1_1_RNO_0[12]_net_1\);
    
    \readData_31_bm_RNO[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[30]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[27]\, D => \readData15[30]\, Y => 
        \readData_31_bm_RNO[27]_net_1\);
    
    \readData_31_bm_1_1_RNO[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[12]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[11]\, D => \readData13[12]\, Y => 
        \readData_31_bm_1_1_RNO[11]_net_1\);
    
    \readData_31_am[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[9]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[9]_net_1\, D
         => \readData_31_am_RNO_0[9]_net_1\, Y => 
        \readData_31_am[9]_net_1\);
    
    \readData_31_am_RNO[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[1]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[1]\, D => \readData14[1]\, Y => 
        \readData_31_am_RNO[1]_net_1\);
    
    \readData_31_am_RNO[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[4]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[4]\, D => \readData14[4]\, Y => 
        \readData_31_am_RNO[4]_net_1\);
    
    block22_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(1), Y => \wen_a_m[1]\);
    
    \readData_31_am_RNO_0[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[22]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[20]\, D => \readData10[22]\, Y => 
        \readData_31_am_RNO_0[20]_net_1\);
    
    \readData_31_am_RNO[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[18]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[16]\, D => \readData14[18]\, Y => 
        \readData_31_am_RNO[16]_net_1\);
    
    \readData_31_ns[27]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[27]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[27]_net_1\, Y => 
        ram_rdata(27));
    
    \readData_31_am_RNO[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[23]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[21]\, D => \readData14[23]\, Y => 
        \readData_31_am_RNO[21]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[13]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[12]\, D => \readData9[13]\, Y => 
        \readData_31_bm_1_1_RNO_0[12]_net_1\);
    
    block0_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem(3), Y => 
        \wen_b0_1[1]\);
    
    \readData_31_bm_RNO_0[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[6]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[6]\, D => \readData11[6]\, Y => 
        \readData_31_bm_RNO_0[6]_net_1\);
    
    \readData_31_bm[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[1]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[1]_net_1\, D
         => \readData_31_bm_RNO_0[1]_net_1\, Y => 
        \readData_31_bm[1]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[1]\, D => \readData1[1]\, Y => 
        \readData_18_1_1[1]\);
    
    \readData_31_bm[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[6]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[6]_net_1\, D
         => \readData_31_bm_RNO_0[6]_net_1\, Y => 
        \readData_31_bm[6]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[10]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[9]\, D => \readData9[10]\, Y => 
        \readData_31_bm_1_1_RNO_0[9]_net_1\);
    
    \readData_31_bm_RNO[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[2]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[2]\, D => \readData15[2]\, Y => 
        \readData_31_bm_RNO[2]_net_1\);
    
    block5_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(3), Y => 
        \wen_b5_1[1]\);
    
    block10_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(0), Y => \wen_a10_1[0]\);
    
    \readData_31_bm_RNO[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[31]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[28]\, D => \readData15[31]\, Y => 
        \readData_31_bm_RNO[28]_net_1\);
    
    \readData_31_bm[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[3]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[3]_net_1\, D
         => \readData_31_bm_RNO_0[3]_net_1\, Y => 
        \readData_31_bm[3]_net_1\);
    
    \readData_31_am_RNO_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[32]\, D => \readData6[32]\, Y => 
        \readData_13_1_1[29]\);
    
    block18_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(14), C
         => readdata_xhdl1401_1, D => sram_wen_mem(3), Y => 
        \wen_b18_1[1]\);
    
    \readData_31_am_1_1_RNO_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[6]\, D => \readData4[6]\, Y => 
        \readData_6_1_1[6]\);
    
    \readData_31_am_RNO[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[3]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[3]\, D => \readData14[3]\, Y => 
        \readData_31_am_RNO[3]_net_1\);
    
    block14_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(0), Y => \wen_a14_1[0]\);
    
    \readData_31_am_RNO_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[27]\, D => \readData6[27]\, Y => 
        \readData_13_1_1[24]\);
    
    \readData_31_bm_1_1_RNO[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[28]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[25]\, D => \readData13[28]\, Y => 
        \readData_31_bm_1_1_RNO[25]_net_1\);
    
    \readData_31_am_RNO_2[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[11]\, D => \readData2[11]\, Y => 
        \readData_10_1_1[10]\);
    
    block0_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem(2), Y => 
        \wen_b0_1[0]\);
    
    \readData_31_bm_1_1_RNO_0[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[1]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[1]\, D => \readData9[1]\, Y => 
        \readData_31_bm_1_1_RNO_0[1]_net_1\);
    
    \readData_31_am_1_1_RNO_0[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[5]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[5]\, D => \readData8[5]\, Y => 
        \readData_31_am_1_1_RNO_0[5]_net_1\);
    
    block28_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(2), Y => \wen_b28_1[0]\);
    
    \readData_31_bm_1_1_RNO_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[25]\, D => \readData5[25]\, Y => 
        \readData_21_1_1[23]\);
    
    \readData_31_bm_RNO[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[12]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[11]\, D => \readData15[12]\, Y => 
        \readData_31_bm_RNO[11]_net_1\);
    
    \readData_31_bm_RNO_2[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[4]\, D => \readData3[4]\, Y => 
        \readData_25_1_1[4]\);
    
    \readData_31_bm[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[17]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[17]_net_1\, D
         => \readData_31_bm_RNO_0[17]_net_1\, Y => 
        \readData_31_bm[17]_net_1\);
    
    \readData_31_am_RNO_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[11]\, D => \readData6[11]\, Y => 
        \readData_13_1_1[10]\);
    
    \readData_31_bm_1_1_RNO[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[23]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[21]\, D => \readData13[23]\, Y => 
        \readData_31_bm_1_1_RNO[21]_net_1\);
    
    \readData_31_bm_1_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[2]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[2]_net_1\, Y => 
        \readData_31_bm_1_1[2]_net_1\);
    
    \readData_31_am_1_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[25]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[25]_net_1\, Y => 
        \readData_31_am_1_1[25]_net_1\);
    
    \readData_31_bm_RNO_2[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[6]\, D => \readData3[6]\, Y => 
        \readData_25_1_1[6]\);
    
    \readData_31_bm_RNO_2[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[33]\, D => \readData3[33]\, Y => 
        \readData_25_1_1[30]\);
    
    \readData_31_ns[30]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[30]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[30]_net_1\, Y => 
        ram_rdata(30));
    
    \readData_31_am_1_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[9]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[9]_net_1\, Y => 
        \readData_31_am_1_1[9]_net_1\);
    
    \readData_31_am_1_1_RNO_0[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[18]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[16]\, D => \readData8[18]\, Y => 
        \readData_31_am_1_1_RNO_0[16]_net_1\);
    
    \readData_31_am_RNO_0[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[25]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[23]\, D => \readData10[25]\, Y => 
        \readData_31_am_RNO_0[23]_net_1\);
    
    \readData_31_am_1_1_RNO_0[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[30]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[27]\, D => \readData8[30]\, Y => 
        \readData_31_am_1_1_RNO_0[27]_net_1\);
    
    \readData_31_bm_RNO[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[18]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[16]\, D => \readData15[18]\, Y => 
        \readData_31_bm_RNO[16]_net_1\);
    
    \readData_31_am_1_1_RNO_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[32]\, D => \readData4[32]\, Y => 
        \readData_6_1_1[29]\);
    
    \readData_31_bm_1_1_RNO_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[3]\, D => \readData5[3]\, Y => 
        \readData_21_1_1[3]\);
    
    \readData_31_bm_RNO[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[11]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[10]\, D => \readData15[11]\, Y => 
        \readData_31_bm_RNO[10]_net_1\);
    
    \readData_31_bm[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[15]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[15]_net_1\, D
         => \readData_31_bm_RNO_0[15]_net_1\, Y => 
        \readData_31_bm[15]_net_1\);
    
    \readData_31_am_1_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[11]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[11]_net_1\, Y => 
        \readData_31_am_1_1[11]_net_1\);
    
    block16_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(3), Y => 
        \wen_b16_1[1]\);
    
    block13_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(3), Y => 
        \wen_b13_1[1]\);
    
    \readData_31_bm_RNO_0[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[1]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[1]\, D => \readData11[1]\, Y => 
        \readData_31_bm_RNO_0[1]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[32]\, D => \readData5[32]\, Y => 
        \readData_21_1_1[29]\);
    
    \readData_31_am_RNO_0[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[9]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[8]\, D => \readData10[9]\, Y => 
        \readData_31_am_RNO_0[8]_net_1\);
    
    \readData_31_am_RNO_2[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[14]\, D => \readData2[14]\, Y => 
        \readData_10_1_1[13]\);
    
    \readData_31_bm_1_1_RNO_2[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[18]\, D => \readData1[18]\, Y => 
        \readData_18_1_1[16]\);
    
    block27 : RAM1K18
      port map(A_DOUT(17) => nc52, A_DOUT(16) => \readData27[16]\, 
        A_DOUT(15) => \readData27[15]\, A_DOUT(14) => 
        \readData27[14]\, A_DOUT(13) => \readData27[13]\, 
        A_DOUT(12) => \readData27[12]\, A_DOUT(11) => 
        \readData27[11]\, A_DOUT(10) => \readData27[10]\, 
        A_DOUT(9) => \readData27[9]\, A_DOUT(8) => nc76, 
        A_DOUT(7) => \readData27[7]\, A_DOUT(6) => 
        \readData27[6]\, A_DOUT(5) => \readData27[5]\, A_DOUT(4)
         => \readData27[4]\, A_DOUT(3) => \readData27[3]\, 
        A_DOUT(2) => \readData27[2]\, A_DOUT(1) => 
        \readData27[1]\, A_DOUT(0) => \readData27[0]\, B_DOUT(17)
         => nc51, B_DOUT(16) => \readData27[34]\, B_DOUT(15) => 
        \readData27[33]\, B_DOUT(14) => \readData27[32]\, 
        B_DOUT(13) => \readData27[31]\, B_DOUT(12) => 
        \readData27[30]\, B_DOUT(11) => \readData27[29]\, 
        B_DOUT(10) => \readData27[28]\, B_DOUT(9) => 
        \readData27[27]\, B_DOUT(8) => nc66, B_DOUT(7) => 
        \readData27[25]\, B_DOUT(6) => \readData27[24]\, 
        B_DOUT(5) => \readData27[23]\, B_DOUT(4) => 
        \readData27[22]\, B_DOUT(3) => \readData27[21]\, 
        B_DOUT(2) => \readData27[20]\, B_DOUT(1) => 
        \readData27[19]\, B_DOUT(0) => \readData27[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a27_1[1]\, 
        A_WEN(0) => \wen_a27_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b27_1[1]\, 
        B_WEN(0) => \wen_b27_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block25_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(0), Y => \wen_a25_1[0]\);
    
    block22_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(0), Y => \wen_a_m[0]\);
    
    \readData_31_bm_RNO_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[29]\, D => \readData7[29]\, Y => 
        \readData_28_1_1[26]\);
    
    \readData_31_bm_1_1_RNO_0[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[31]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[28]\, D => \readData9[31]\, Y => 
        \readData_31_bm_1_1_RNO_0[28]_net_1\);
    
    \readData_31_bm_RNO_0[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[27]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[24]\, D => \readData11[27]\, Y => 
        \readData_31_bm_RNO_0[24]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[18]\, D => \readData5[18]\, Y => 
        \readData_21_1_1[16]\);
    
    \readData_31_am_RNO_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[14]\, D => \readData6[14]\, Y => 
        \readData_13_1_1[13]\);
    
    \readData_31_am_1_1_RNO[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[33]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[30]\, D => \readData12[33]\, Y => 
        \readData_31_am_1_1_RNO[30]_net_1\);
    
    block13_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(1), Y => 
        \wen_a13_1[1]\);
    
    \readData_31_bm_RNO_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[32]\, D => \readData7[32]\, Y => 
        \readData_28_1_1[29]\);
    
    \readData_31_am_1_1_RNO_2[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[30]\, D => \readData0[30]\, Y => 
        \readData_3_1_1[27]\);
    
    block27_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(1), Y => \wen_a27_1[1]\);
    
    \readData_31_am_1_1_RNO_2[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[13]\, D => \readData0[13]\, Y => 
        \readData_3_1_1[12]\);
    
    \readData_31_ns[18]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[18]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[18]_net_1\, Y => 
        ram_rdata(18));
    
    \readData_31_bm_RNO_0[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[12]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[11]\, D => \readData11[12]\, Y => 
        \readData_31_bm_RNO_0[11]_net_1\);
    
    \readData_31_bm_RNO[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[7]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[7]\, D => \readData15[7]\, Y => 
        \readData_31_bm_RNO[7]_net_1\);
    
    \readData_31_ns[19]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[19]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[19]_net_1\, Y => 
        ram_rdata(19));
    
    \readData_31_am_1_1_RNO_2[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[2]\, D => \readData0[2]\, Y => 
        \readData_3_1_1[2]\);
    
    \readData_31_am_1_1_RNO_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[13]\, D => \readData4[13]\, Y => 
        \readData_6_1_1[12]\);
    
    \readData_31_bm_1_1_RNO_2[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[13]\, D => \readData1[13]\, Y => 
        \readData_18_1_1[12]\);
    
    \readData_31_am_RNO_0[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[12]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[11]\, D => \readData10[12]\, Y => 
        \readData_31_am_RNO_0[11]_net_1\);
    
    \readData_31_bm_RNO_2[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[15]\, D => \readData3[15]\, Y => 
        \readData_25_1_1[14]\);
    
    \readData_31_bm[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[4]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[4]_net_1\, D
         => \readData_31_bm_RNO_0[4]_net_1\, Y => 
        \readData_31_bm[4]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[13]\, D => \readData5[13]\, Y => 
        \readData_21_1_1[12]\);
    
    block30 : RAM1K18
      port map(A_DOUT(17) => nc77, A_DOUT(16) => \readData30[16]\, 
        A_DOUT(15) => \readData30[15]\, A_DOUT(14) => 
        \readData30[14]\, A_DOUT(13) => \readData30[13]\, 
        A_DOUT(12) => \readData30[12]\, A_DOUT(11) => 
        \readData30[11]\, A_DOUT(10) => \readData30[10]\, 
        A_DOUT(9) => \readData30[9]\, A_DOUT(8) => nc67, 
        A_DOUT(7) => \readData30[7]\, A_DOUT(6) => 
        \readData30[6]\, A_DOUT(5) => \readData30[5]\, A_DOUT(4)
         => \readData30[4]\, A_DOUT(3) => \readData30[3]\, 
        A_DOUT(2) => \readData30[2]\, A_DOUT(1) => 
        \readData30[1]\, A_DOUT(0) => \readData30[0]\, B_DOUT(17)
         => nc4, B_DOUT(16) => \readData30[34]\, B_DOUT(15) => 
        \readData30[33]\, B_DOUT(14) => \readData30[32]\, 
        B_DOUT(13) => \readData30[31]\, B_DOUT(12) => 
        \readData30[30]\, B_DOUT(11) => \readData30[29]\, 
        B_DOUT(10) => \readData30[28]\, B_DOUT(9) => 
        \readData30[27]\, B_DOUT(8) => nc124, B_DOUT(7) => 
        \readData30[25]\, B_DOUT(6) => \readData30[24]\, 
        B_DOUT(5) => \readData30[23]\, B_DOUT(4) => 
        \readData30[22]\, B_DOUT(3) => \readData30[21]\, 
        B_DOUT(2) => \readData30[20]\, B_DOUT(1) => 
        \readData30[19]\, B_DOUT(0) => \readData30[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a30_1[1]\, 
        A_WEN(0) => \wen_a30_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b30_1[1]\, 
        B_WEN(0) => \wen_b30_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_RNO_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[2]\, D => \readData6[2]\, Y => 
        \readData_13_1_1[2]\);
    
    \readData_31_bm_RNO_2[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[5]\, D => \readData3[5]\, Y => 
        \readData_25_1_1[5]\);
    
    block8_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(3), Y => \wen_b8_1[1]\);
    
    \readData_31_bm_RNO_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[15]\, D => \readData7[15]\, Y => 
        \readData_28_1_1[14]\);
    
    \readData_31_bm_1_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[4]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[4]_net_1\, Y => 
        \readData_31_bm_1_1[4]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[15]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[14]\, D => \readData9[15]\, Y => 
        \readData_31_bm_1_1_RNO_0[14]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[31]\, D => \readData1[31]\, Y => 
        \readData_18_1_1[28]\);
    
    \readData_31_am_1_1_RNO_2[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[6]\, D => \readData0[6]\, Y => 
        \readData_3_1_1[6]\);
    
    \readData_31_bm_RNO_0[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[4]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[4]\, D => \readData11[4]\, Y => 
        \readData_31_bm_RNO_0[4]_net_1\);
    
    \readData_31_bm_RNO[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[25]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[23]\, D => \readData15[25]\, Y => 
        \readData_31_bm_RNO[23]_net_1\);
    
    \readData_31_am_1_1_RNO[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[7]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[7]\, D => \readData12[7]\, Y => 
        \readData_31_am_1_1_RNO[7]_net_1\);
    
    \readData_31_ns[23]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[23]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[23]_net_1\, Y => 
        ram_rdata(23));
    
    \readData_31_am_1_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[13]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[13]_net_1\, Y => 
        \readData_31_am_1_1[13]_net_1\);
    
    block31_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(2), Y => \wen_b31_1[0]\);
    
    block29_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(1), Y => \wen_a29_1[1]\);
    
    \readData_31_bm[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[9]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[9]_net_1\, D
         => \readData_31_bm_RNO_0[9]_net_1\, Y => 
        \readData_31_bm[9]_net_1\);
    
    \readData_31_bm_RNO_2[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[23]\, D => \readData3[23]\, Y => 
        \readData_25_1_1[21]\);
    
    \readData_31_am_RNO_0[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[19]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[17]\, D => \readData10[19]\, Y => 
        \readData_31_am_RNO_0[17]_net_1\);
    
    \readData_31_bm_RNO_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[25]\, D => \readData7[25]\, Y => 
        \readData_28_1_1[23]\);
    
    block4 : RAM1K18
      port map(A_DOUT(17) => nc109, A_DOUT(16) => \readData4[16]\, 
        A_DOUT(15) => \readData4[15]\, A_DOUT(14) => 
        \readData4[14]\, A_DOUT(13) => \readData4[13]\, 
        A_DOUT(12) => \readData4[12]\, A_DOUT(11) => 
        \readData4[11]\, A_DOUT(10) => \readData4[10]\, A_DOUT(9)
         => \readData4[9]\, A_DOUT(8) => nc42, A_DOUT(7) => 
        \readData4[7]\, A_DOUT(6) => \readData4[6]\, A_DOUT(5)
         => \readData4[5]\, A_DOUT(4) => \readData4[4]\, 
        A_DOUT(3) => \readData4[3]\, A_DOUT(2) => \readData4[2]\, 
        A_DOUT(1) => \readData4[1]\, A_DOUT(0) => \readData4[0]\, 
        B_DOUT(17) => nc114, B_DOUT(16) => \readData4[34]\, 
        B_DOUT(15) => \readData4[33]\, B_DOUT(14) => 
        \readData4[32]\, B_DOUT(13) => \readData4[31]\, 
        B_DOUT(12) => \readData4[30]\, B_DOUT(11) => 
        \readData4[29]\, B_DOUT(10) => \readData4[28]\, B_DOUT(9)
         => \readData4[27]\, B_DOUT(8) => nc100, B_DOUT(7) => 
        \readData4[25]\, B_DOUT(6) => \readData4[24]\, B_DOUT(5)
         => \readData4[23]\, B_DOUT(4) => \readData4[22]\, 
        B_DOUT(3) => \readData4[21]\, B_DOUT(2) => 
        \readData4[20]\, B_DOUT(1) => \readData4[19]\, B_DOUT(0)
         => \readData4[18]\, BUSY => OPEN, A_CLK => FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_21_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a4_1[1]\, 
        A_WEN(0) => \wen_a4_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b4_1[1]\, 
        B_WEN(0) => \wen_b4_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block20_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(0), Y => \wen_a20_1[0]\);
    
    \readData_31_am_RNO_2[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[23]\, D => \readData2[23]\, Y => 
        \readData_10_1_1[21]\);
    
    \readData_31_bm_RNO_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[22]\, D => \readData7[22]\, Y => 
        \readData_28_1_1[20]\);
    
    \readData_31_am_1_1_RNO_2[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[7]\, D => \readData0[7]\, Y => 
        \readData_3_1_1[7]\);
    
    \readData_31_am_RNO_0[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[20]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[18]\, D => \readData10[20]\, Y => 
        \readData_31_am_RNO_0[18]_net_1\);
    
    \readData_31_am_1_1_RNO_0[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[11]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[10]\, D => \readData8[11]\, Y => 
        \readData_31_am_1_1_RNO_0[10]_net_1\);
    
    \wen_a_m_30_0_a2_0[1]\ : CFG3
      generic map(INIT => x"20")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1144);
    
    block24_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(0), Y => \wen_a24_1[0]\);
    
    \readData_31_am_1_1_RNO_2[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[18]\, D => \readData0[18]\, Y => 
        \readData_3_1_1[16]\);
    
    \readData_31_am_1_1_RNO[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[20]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[18]\, D => \readData12[20]\, Y => 
        \readData_31_am_1_1_RNO[18]_net_1\);
    
    \readData_31_bm_1_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[17]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[17]_net_1\, Y => 
        \readData_31_bm_1_1[17]_net_1\);
    
    \readData_31_am_RNO[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[21]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[19]\, D => \readData14[21]\, Y => 
        \readData_31_am_RNO[19]_net_1\);
    
    \readData_31_am_1_1_RNO_2[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[34]\, D => \readData0[34]\, Y => 
        \readData_3_1_1[31]\);
    
    \readData_31_am_1_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[28]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[28]_net_1\, Y => 
        \readData_31_am_1_1[28]_net_1\);
    
    \readData_31_am_1_1_RNO_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[18]\, D => \readData4[18]\, Y => 
        \readData_6_1_1[16]\);
    
    block27_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(3), Y => \wen_b27_1[1]\);
    
    \readData_31_am_1_1_RNO_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[34]\, D => \readData4[34]\, Y => 
        \readData_6_1_1[31]\);
    
    \readData_31_bm_1_1_RNO_2[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[33]\, D => \readData1[33]\, Y => 
        \readData_18_1_1[30]\);
    
    \readData_31_bm_1_1_RNO_0[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[28]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[25]\, D => \readData9[28]\, Y => 
        \readData_31_bm_1_1_RNO_0[25]_net_1\);
    
    block1 : RAM1K18
      port map(A_DOUT(17) => nc83, A_DOUT(16) => \readData1[16]\, 
        A_DOUT(15) => \readData1[15]\, A_DOUT(14) => 
        \readData1[14]\, A_DOUT(13) => \readData1[13]\, 
        A_DOUT(12) => \readData1[12]\, A_DOUT(11) => 
        \readData1[11]\, A_DOUT(10) => \readData1[10]\, A_DOUT(9)
         => \readData1[9]\, A_DOUT(8) => nc41, A_DOUT(7) => 
        \readData1[7]\, A_DOUT(6) => \readData1[6]\, A_DOUT(5)
         => \readData1[5]\, A_DOUT(4) => \readData1[4]\, 
        A_DOUT(3) => \readData1[3]\, A_DOUT(2) => \readData1[2]\, 
        A_DOUT(1) => \readData1[1]\, A_DOUT(0) => \readData1[0]\, 
        B_DOUT(17) => nc90, B_DOUT(16) => \readData1[34]\, 
        B_DOUT(15) => \readData1[33]\, B_DOUT(14) => 
        \readData1[32]\, B_DOUT(13) => \readData1[31]\, 
        B_DOUT(12) => \readData1[30]\, B_DOUT(11) => 
        \readData1[29]\, B_DOUT(10) => \readData1[28]\, B_DOUT(9)
         => \readData1[27]\, B_DOUT(8) => nc94, B_DOUT(7) => 
        \readData1[25]\, B_DOUT(6) => \readData1[24]\, B_DOUT(5)
         => \readData1[23]\, B_DOUT(4) => \readData1[22]\, 
        B_DOUT(3) => \readData1[21]\, B_DOUT(2) => 
        \readData1[20]\, B_DOUT(1) => \readData1[19]\, B_DOUT(0)
         => \readData1[18]\, BUSY => OPEN, A_CLK => FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_21_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a1_1[1]\, 
        A_WEN(0) => \wen_a1_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b1_1[1]\, 
        B_WEN(0) => \wen_b1_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_1_1_RNO_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[33]\, D => \readData5[33]\, Y => 
        \readData_21_1_1[30]\);
    
    block5_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(0), Y => 
        \wen_a5_1[0]\);
    
    \readData_31_bm_1_1_RNO_2[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[3]\, D => \readData1[3]\, Y => 
        \readData_18_1_1[3]\);
    
    \readData_31_am_RNO_2[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[30]\, D => \readData2[30]\, Y => 
        \readData_10_1_1[27]\);
    
    \readData_31_am_1_1_RNO[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[21]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[19]\, D => \readData12[21]\, Y => 
        \readData_31_am_1_1_RNO[19]_net_1\);
    
    block27_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(2), Y => \wen_b27_1[0]\);
    
    \readData_31_am_RNO_2[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[31]\, D => \readData2[31]\, Y => 
        \readData_10_1_1[28]\);
    
    \readData_31_am_1_1_RNO_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[30]\, D => \readData4[30]\, Y => 
        \readData_6_1_1[27]\);
    
    readdata_xhdl1400_0_a2_0 : CFG3
      generic map(INIT => x"02")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1168);
    
    \readData_31_bm_1_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[14]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[14]_net_1\, Y => 
        \readData_31_bm_1_1[14]_net_1\);
    
    \readData_31_am_RNO_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[5]\, D => \readData6[5]\, Y => 
        \readData_13_1_1[5]\);
    
    block14_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(2), Y => \wen_b14_1[0]\);
    
    \readData_31_bm_1_1_RNO_2[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[34]\, D => \readData1[34]\, Y => 
        \readData_18_1_1[31]\);
    
    \readData_31_am_1_1_RNO_0[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[0]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[0]\, D => \readData8[0]\, Y => 
        \readData_31_am_1_1_RNO_0[0]_net_1\);
    
    \readData_31_am_RNO[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[24]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[22]\, D => \readData14[24]\, Y => 
        \readData_31_am_RNO[22]_net_1\);
    
    \readData_31_bm_RNO[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[24]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[22]\, D => \readData15[24]\, Y => 
        \readData_31_bm_RNO[22]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[10]\, D => \readData1[10]\, Y => 
        \readData_18_1_1[9]\);
    
    \readData_31_bm_1_1_RNO[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[11]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[10]\, D => \readData13[11]\, Y => 
        \readData_31_bm_1_1_RNO[10]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[34]\, D => \readData5[34]\, Y => 
        \readData_21_1_1[31]\);
    
    \readData_31_am_RNO[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[2]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[2]\, D => \readData14[2]\, Y => 
        \readData_31_am_RNO[2]_net_1\);
    
    block5_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(1), Y => 
        \wen_a5_1[1]\);
    
    \readData_31_am_1_1_RNO[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[12]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[11]\, D => \readData12[12]\, Y => 
        \readData_31_am_1_1_RNO[11]_net_1\);
    
    block19 : RAM1K18
      port map(A_DOUT(17) => nc122, A_DOUT(16) => 
        \readData19[16]\, A_DOUT(15) => \readData19[15]\, 
        A_DOUT(14) => \readData19[14]\, A_DOUT(13) => 
        \readData19[13]\, A_DOUT(12) => \readData19[12]\, 
        A_DOUT(11) => \readData19[11]\, A_DOUT(10) => 
        \readData19[10]\, A_DOUT(9) => \readData19[9]\, A_DOUT(8)
         => nc112, A_DOUT(7) => \readData19[7]\, A_DOUT(6) => 
        \readData19[6]\, A_DOUT(5) => \readData19[5]\, A_DOUT(4)
         => \readData19[4]\, A_DOUT(3) => \readData19[3]\, 
        A_DOUT(2) => \readData19[2]\, A_DOUT(1) => 
        \readData19[1]\, A_DOUT(0) => \readData19[0]\, B_DOUT(17)
         => nc86, B_DOUT(16) => \readData19[34]\, B_DOUT(15) => 
        \readData19[33]\, B_DOUT(14) => \readData19[32]\, 
        B_DOUT(13) => \readData19[31]\, B_DOUT(12) => 
        \readData19[30]\, B_DOUT(11) => \readData19[29]\, 
        B_DOUT(10) => \readData19[28]\, B_DOUT(9) => 
        \readData19[27]\, B_DOUT(8) => nc59, B_DOUT(7) => 
        \readData19[25]\, B_DOUT(6) => \readData19[24]\, 
        B_DOUT(5) => \readData19[23]\, B_DOUT(4) => 
        \readData19[22]\, B_DOUT(3) => \readData19[21]\, 
        B_DOUT(2) => \readData19[20]\, B_DOUT(1) => 
        \readData19[19]\, B_DOUT(0) => \readData19[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a19_1[1]\, 
        A_WEN(0) => \wen_a19_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b19_1[1]\, 
        B_WEN(0) => \wen_b19_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    readdata_xhdl1406_1 : CFG3
      generic map(INIT => x"20")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => ahbsram_addr(13), Y => readdata_xhdl1414_1);
    
    \readData_31_am_1_1_RNO[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[31]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[28]\, D => \readData12[31]\, Y => 
        \readData_31_am_1_1_RNO[28]_net_1\);
    
    \readData_31_ns[11]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[11]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[11]_net_1\, Y => 
        ram_rdata(11));
    
    \readData_31_ns[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[1]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[1]_net_1\, Y => 
        ram_rdata(1));
    
    block0_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem(1), Y => 
        \wen_a0_1[1]\);
    
    \readData_31_bm_RNO_0[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[28]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[25]\, D => \readData11[28]\, Y => 
        \readData_31_bm_RNO_0[25]_net_1\);
    
    block11_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(2), Y => \wen_b11_1[0]\);
    
    \readData_31_ns[20]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[20]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[20]_net_1\, Y => 
        ram_rdata(20));
    
    \readData_31_bm_1_1_RNO[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[20]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[18]\, D => \readData13[20]\, Y => 
        \readData_31_bm_1_1_RNO[18]_net_1\);
    
    \readData_31_ns[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[7]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[7]_net_1\, Y => 
        ram_rdata(7));
    
    \readData_31_bm_1_1_RNO_2[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[28]\, D => \readData1[28]\, Y => 
        \readData_18_1_1[25]\);
    
    \readData_31_bm_1_1_RNO_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[31]\, D => \readData5[31]\, Y => 
        \readData_21_1_1[28]\);
    
    block2_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(2), Y => \wen_b2_1[0]\);
    
    \readData_31_am_1_1_RNO[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[32]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[29]\, D => \readData12[32]\, Y => 
        \readData_31_am_1_1_RNO[29]_net_1\);
    
    block5_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(2), Y => 
        \wen_b5_1[0]\);
    
    block14 : RAM1K18
      port map(A_DOUT(17) => nc25, A_DOUT(16) => \readData14[16]\, 
        A_DOUT(15) => \readData14[15]\, A_DOUT(14) => 
        \readData14[14]\, A_DOUT(13) => \readData14[13]\, 
        A_DOUT(12) => \readData14[12]\, A_DOUT(11) => 
        \readData14[11]\, A_DOUT(10) => \readData14[10]\, 
        A_DOUT(9) => \readData14[9]\, A_DOUT(8) => nc15, 
        A_DOUT(7) => \readData14[7]\, A_DOUT(6) => 
        \readData14[6]\, A_DOUT(5) => \readData14[5]\, A_DOUT(4)
         => \readData14[4]\, A_DOUT(3) => \readData14[3]\, 
        A_DOUT(2) => \readData14[2]\, A_DOUT(1) => 
        \readData14[1]\, A_DOUT(0) => \readData14[0]\, B_DOUT(17)
         => nc87, B_DOUT(16) => \readData14[34]\, B_DOUT(15) => 
        \readData14[33]\, B_DOUT(14) => \readData14[32]\, 
        B_DOUT(13) => \readData14[31]\, B_DOUT(12) => 
        \readData14[30]\, B_DOUT(11) => \readData14[29]\, 
        B_DOUT(10) => \readData14[28]\, B_DOUT(9) => 
        \readData14[27]\, B_DOUT(8) => nc35, B_DOUT(7) => 
        \readData14[25]\, B_DOUT(6) => \readData14[24]\, 
        B_DOUT(5) => \readData14[23]\, B_DOUT(4) => 
        \readData14[22]\, B_DOUT(3) => \readData14[21]\, 
        B_DOUT(2) => \readData14[20]\, B_DOUT(1) => 
        \readData14[19]\, B_DOUT(0) => \readData14[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a14_1[1]\, 
        A_WEN(0) => \wen_a14_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b14_1[1]\, 
        B_WEN(0) => \wen_b14_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[6]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[6]\, D => \readData15[6]\, Y => 
        \readData_31_bm_RNO[6]_net_1\);
    
    \readData_31_ns[9]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[9]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[9]_net_1\, Y => 
        ram_rdata(9));
    
    block12_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(3), Y => \wen_b12_1[1]\);
    
    \readData_31_bm_1_1_RNO_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[6]\, D => \readData5[6]\, Y => 
        \readData_21_1_1[6]\);
    
    \readData_31_am_1_1_RNO_0[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[23]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[21]\, D => \readData8[23]\, Y => 
        \readData_31_am_1_1_RNO_0[21]_net_1\);
    
    \readData_31_am[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[31]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[31]_net_1\, D
         => \readData_31_am_RNO_0[31]_net_1\, Y => 
        \readData_31_am[31]_net_1\);
    
    \readData_31_bm_1_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[3]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[3]_net_1\, Y => 
        \readData_31_bm_1_1[3]_net_1\);
    
    \readData_31_am[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[26]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[26]_net_1\, D
         => \readData_31_am_RNO_0[26]_net_1\, Y => 
        \readData_31_am[26]_net_1\);
    
    \readData_31_bm_RNO_2[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[16]\, D => \readData3[16]\, Y => 
        \readData_25_1_1[15]\);
    
    \readData_31_bm_1_1_RNO_0[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[5]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[5]\, D => \readData9[5]\, Y => 
        \readData_31_bm_1_1_RNO_0[5]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[22]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[20]\, D => \readData9[22]\, Y => 
        \readData_31_bm_1_1_RNO_0[20]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[15]\, D => \readData1[15]\, Y => 
        \readData_18_1_1[14]\);
    
    \readData_31_bm[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[10]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[10]_net_1\, D
         => \readData_31_bm_RNO_0[10]_net_1\, Y => 
        \readData_31_bm[10]_net_1\);
    
    \readData_31_am[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[29]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[29]_net_1\, D
         => \readData_31_am_RNO_0[29]_net_1\, Y => 
        \readData_31_am[29]_net_1\);
    
    block29_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(2), Y => \wen_b29_1[0]\);
    
    \readData_31_bm_RNO_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[1]\, D => \readData7[1]\, Y => 
        \readData_28_1_1[1]\);
    
    \readData_31_bm_1_1_RNO[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[22]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[20]\, D => \readData13[22]\, Y => 
        \readData_31_bm_1_1_RNO[20]_net_1\);
    
    block14_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(3), Y => \wen_b14_1[1]\);
    
    \readData_31_ns[24]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[24]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[24]_net_1\, Y => 
        ram_rdata(24));
    
    \readData_31_bm_1_1_RNO_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[15]\, D => \readData5[15]\, Y => 
        \readData_21_1_1[14]\);
    
    block15 : RAM1K18
      port map(A_DOUT(17) => nc49, A_DOUT(16) => \readData15[16]\, 
        A_DOUT(15) => \readData15[15]\, A_DOUT(14) => 
        \readData15[14]\, A_DOUT(13) => \readData15[13]\, 
        A_DOUT(12) => \readData15[12]\, A_DOUT(11) => 
        \readData15[11]\, A_DOUT(10) => \readData15[10]\, 
        A_DOUT(9) => \readData15[9]\, A_DOUT(8) => nc28, 
        A_DOUT(7) => \readData15[7]\, A_DOUT(6) => 
        \readData15[6]\, A_DOUT(5) => \readData15[5]\, A_DOUT(4)
         => \readData15[4]\, A_DOUT(3) => \readData15[3]\, 
        A_DOUT(2) => \readData15[2]\, A_DOUT(1) => 
        \readData15[1]\, A_DOUT(0) => \readData15[0]\, B_DOUT(17)
         => nc18, B_DOUT(16) => \readData15[34]\, B_DOUT(15) => 
        \readData15[33]\, B_DOUT(14) => \readData15[32]\, 
        B_DOUT(13) => \readData15[31]\, B_DOUT(12) => 
        \readData15[30]\, B_DOUT(11) => \readData15[29]\, 
        B_DOUT(10) => \readData15[28]\, B_DOUT(9) => 
        \readData15[27]\, B_DOUT(8) => nc128, B_DOUT(7) => 
        \readData15[25]\, B_DOUT(6) => \readData15[24]\, 
        B_DOUT(5) => \readData15[23]\, B_DOUT(4) => 
        \readData15[22]\, B_DOUT(3) => \readData15[21]\, 
        B_DOUT(2) => \readData15[20]\, B_DOUT(1) => 
        \readData15[19]\, B_DOUT(0) => \readData15[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a15_1[1]\, 
        A_WEN(0) => \wen_a15_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b15_1[1]\, 
        B_WEN(0) => \wen_b15_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[16]\, D => \readData7[16]\, Y => 
        \readData_28_1_1[15]\);
    
    \readData_31_bm_1_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[20]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[20]_net_1\, Y => 
        \readData_31_bm_1_1[20]_net_1\);
    
    \readData_31_am_1_1_RNO[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[23]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[21]\, D => \readData12[23]\, Y => 
        \readData_31_am_1_1_RNO[21]_net_1\);
    
    \readData_31_am_1_1_RNO_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[2]\, D => \readData4[2]\, Y => 
        \readData_6_1_1[2]\);
    
    \readData_31_bm_1_1_RNO[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[31]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[28]\, D => \readData13[31]\, Y => 
        \readData_31_bm_1_1_RNO[28]_net_1\);
    
    readdata_xhdl1388_0_a2_1 : CFG3
      generic map(INIT => x"80")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1148);
    
    \readData_31_bm_1_1_RNO_0[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[23]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[21]\, D => \readData9[23]\, Y => 
        \readData_31_bm_1_1_RNO_0[21]_net_1\);
    
    \readData_31_am_RNO_0[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[11]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[10]\, D => \readData10[11]\, Y => 
        \readData_31_am_RNO_0[10]_net_1\);
    
    \readData_31_bm_1_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[1]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[1]_net_1\, Y => 
        \readData_31_bm_1_1[1]_net_1\);
    
    \readData_31_am_1_1_RNO_0[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[15]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[14]\, D => \readData8[15]\, Y => 
        \readData_31_am_1_1_RNO_0[14]_net_1\);
    
    \readData_31_am_1_1_RNO_2[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[11]\, D => \readData0[11]\, Y => 
        \readData_3_1_1[10]\);
    
    \readData_31_bm_1_1_RNO_0[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[30]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[27]\, D => \readData9[30]\, Y => 
        \readData_31_bm_1_1_RNO_0[27]_net_1\);
    
    \readData_31_am_1_1_RNO_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[11]\, D => \readData4[11]\, Y => 
        \readData_6_1_1[10]\);
    
    block20_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(3), Y => \wen_b20_1[1]\);
    
    \readData_31_am_1_1_RNO_0[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[16]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[15]\, D => \readData8[16]\, Y => 
        \readData_31_am_1_1_RNO_0[15]_net_1\);
    
    block3_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(3), Y => \wen_b3_1[1]\);
    
    readdata_xhdl1418_0_a2 : CFG3
      generic map(INIT => x"40")

      port map(A => ahbsram_addr(15), B => 
        readdata_xhdl1419_0_a2_0, C => ahbsram_addr(11), Y => 
        wen_a3133);
    
    \readData_31_am_1_1_RNO_2[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[23]\, D => \readData0[23]\, Y => 
        \readData_3_1_1[21]\);
    
    \readData_31_bm_RNO_2[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[10]\, D => \readData3[10]\, Y => 
        \readData_25_1_1[9]\);
    
    \readData_31_am[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[25]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[25]_net_1\, D
         => \readData_31_am_RNO_0[25]_net_1\, Y => 
        \readData_31_am[25]_net_1\);
    
    readdata_xhdl1402_0 : CFG3
      generic map(INIT => x"01")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => readdata_xhdl1403_0);
    
    \readData_31_bm_1_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[30]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[30]_net_1\, Y => 
        \readData_31_bm_1_1[30]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[22]\, D => \readData1[22]\, Y => 
        \readData_18_1_1[20]\);
    
    block3_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(1), Y => \wen_a3_1[1]\);
    
    block25_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(3), Y => \wen_b25_1[1]\);
    
    block26_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(2), Y => \wen_b26_1[0]\);
    
    \readData_31_bm_1_1_RNO[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[13]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[12]\, D => \readData13[13]\, Y => 
        \readData_31_bm_1_1_RNO[12]_net_1\);
    
    \readData_31_am_1_1_RNO_0[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[2]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[2]\, D => \readData8[2]\, Y => 
        \readData_31_am_1_1_RNO_0[2]_net_1\);
    
    \readData_31_am_RNO[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[7]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[7]\, D => \readData14[7]\, Y => 
        \readData_31_am_RNO[7]_net_1\);
    
    \readData_31_am_RNO_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[4]\, D => \readData6[4]\, Y => 
        \readData_13_1_1[4]\);
    
    \readData_31_am_RNO_2[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[22]\, D => \readData2[22]\, Y => 
        \readData_10_1_1[20]\);
    
    \readData_31_ns[17]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[17]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[17]_net_1\, Y => 
        ram_rdata(17));
    
    readdata_xhdl1407_0_a2_1 : CFG3
      generic map(INIT => x"40")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1149);
    
    \readData_31_am_RNO[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[11]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[10]\, D => \readData14[11]\, Y => 
        \readData_31_am_RNO[10]_net_1\);
    
    \readData_31_am_RNO_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[6]\, D => \readData6[6]\, Y => 
        \readData_13_1_1[6]\);
    
    \readData_31_bm_1_1_RNO_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[28]\, D => \readData5[28]\, Y => 
        \readData_21_1_1[25]\);
    
    \readData_31_bm_1_1_RNO_2[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[23]\, D => \readData1[23]\, Y => 
        \readData_18_1_1[21]\);
    
    \readData_31_am[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[28]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[28]_net_1\, D
         => \readData_31_am_RNO_0[28]_net_1\, Y => 
        \readData_31_am[28]_net_1\);
    
    \readData_31_bm_RNO_2[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[3]\, D => \readData3[3]\, Y => 
        \readData_25_1_1[3]\);
    
    \readData_31_bm_1_1_RNO_2[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[30]\, D => \readData1[30]\, Y => 
        \readData_18_1_1[27]\);
    
    \readData_31_am_RNO_0[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[14]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[13]\, D => \readData10[14]\, Y => 
        \readData_31_am_RNO_0[13]_net_1\);
    
    \readData_31_am_RNO_0[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[7]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[7]\, D => \readData10[7]\, Y => 
        \readData_31_am_RNO_0[7]_net_1\);
    
    \readData_31_am_1_1_RNO_0[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[7]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[7]\, D => \readData8[7]\, Y => 
        \readData_31_am_1_1_RNO_0[7]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[2]\, D => \readData1[2]\, Y => 
        \readData_18_1_1[2]\);
    
    \readData_31_am[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[20]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[20]_net_1\, D
         => \readData_31_am_RNO_0[20]_net_1\, Y => 
        \readData_31_am[20]_net_1\);
    
    \readData_31_am_RNO[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[25]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[23]\, D => \readData14[25]\, Y => 
        \readData_31_am_RNO[23]_net_1\);
    
    block17_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(0), Y => 
        \wen_a17_1[0]\);
    
    \readData_31_am_1_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[21]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[21]_net_1\, Y => 
        \readData_31_am_1_1[21]_net_1\);
    
    \readData_31_bm_1_1_RNO[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[24]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[22]\, D => \readData13[24]\, Y => 
        \readData_31_bm_1_1_RNO[22]_net_1\);
    
    \readData_31_am_RNO_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[28]\, D => \readData6[28]\, Y => 
        \readData_13_1_1[25]\);
    
    \readData_31_bm_RNO_0[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[31]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[28]\, D => \readData11[31]\, Y => 
        \readData_31_bm_RNO_0[28]_net_1\);
    
    block22_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(2), Y => \wen_b22_1[0]\);
    
    \readData_31_bm_RNO_2[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[7]\, D => \readData3[7]\, Y => 
        \readData_25_1_1[7]\);
    
    \readData_31_bm_1_1_RNO_2[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[6]\, D => \readData1[6]\, Y => 
        \readData_18_1_1[6]\);
    
    \readData_31_bm[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[21]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[21]_net_1\, D
         => \readData_31_bm_RNO_0[21]_net_1\, Y => 
        \readData_31_bm[21]_net_1\);
    
    \readData_31_am_RNO_2[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[25]\, D => \readData2[25]\, Y => 
        \readData_10_1_1[23]\);
    
    \readData_31_am_1_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[10]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[10]_net_1\, Y => 
        \readData_31_am_1_1[10]_net_1\);
    
    \readData_31_bm_RNO_0[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[15]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[14]\, D => \readData11[15]\, Y => 
        \readData_31_bm_RNO_0[14]_net_1\);
    
    block4_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(0), Y => \wen_a4_1[0]\);
    
    block30_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(2), Y => \wen_b30_1[0]\);
    
    \readData_31_am_1_1_RNO[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[13]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[12]\, D => \readData12[13]\, Y => 
        \readData_31_am_1_1_RNO[12]_net_1\);
    
    \readData_31_bm_1_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[13]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[13]_net_1\, Y => 
        \readData_31_bm_1_1[13]_net_1\);
    
    \readData_31_bm_RNO_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[30]\, D => \readData7[30]\, Y => 
        \readData_28_1_1[27]\);
    
    \readData_31_bm_1_1_RNO_2[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[7]\, D => \readData1[7]\, Y => 
        \readData_18_1_1[7]\);
    
    block15_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(2), Y => \wen_b15_1[0]\);
    
    \readData_31_bm_RNO_2[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[20]\, D => \readData3[20]\, Y => 
        \readData_25_1_1[18]\);
    
    \readData_31_am_1_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[31]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[31]_net_1\, Y => 
        \readData_31_am_1_1[31]_net_1\);
    
    \readData_31_am_1_1_RNO_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[23]\, D => \readData4[23]\, Y => 
        \readData_6_1_1[21]\);
    
    block23_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(2), Y => \wen_b23_1[0]\);
    
    \readData_31_bm_1_1_RNO[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[5]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[5]\, D => \readData13[5]\, Y => 
        \readData_31_bm_1_1_RNO[5]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[22]\, D => \readData5[22]\, Y => 
        \readData_21_1_1[20]\);
    
    block9_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(0), Y => \wen_a9_1[0]\);
    
    \readData_31_bm_RNO_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[20]\, D => \readData7[20]\, Y => 
        \readData_28_1_1[18]\);
    
    \readData_31_am_RNO_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[3]\, D => \readData6[3]\, Y => 
        \readData_13_1_1[3]\);
    
    \readData_31_am_1_1_RNO_2[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[15]\, D => \readData0[15]\, Y => 
        \readData_3_1_1[14]\);
    
    \readData_31_am_1_1_RNO_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[5]\, D => \readData4[5]\, Y => 
        \readData_6_1_1[5]\);
    
    \readData_31_am_1_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[17]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[17]_net_1\, Y => 
        \readData_31_am_1_1[17]_net_1\);
    
    \readData_31_am_RNO[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[27]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[24]\, D => \readData14[27]\, Y => 
        \readData_31_am_RNO[24]_net_1\);
    
    \readData_31_am_1_1_RNO_2[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[0]\, D => \readData0[0]\, Y => 
        \readData_3_1_1[0]\);
    
    block19_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(3), Y => \wen_b19_1[1]\);
    
    \readData_31_am_1_1_RNO_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[15]\, D => \readData4[15]\, Y => 
        \readData_6_1_1[14]\);
    
    block6 : RAM1K18
      port map(A_DOUT(17) => nc107, A_DOUT(16) => \readData6[16]\, 
        A_DOUT(15) => \readData6[15]\, A_DOUT(14) => 
        \readData6[14]\, A_DOUT(13) => \readData6[13]\, 
        A_DOUT(12) => \readData6[12]\, A_DOUT(11) => 
        \readData6[11]\, A_DOUT(10) => \readData6[10]\, A_DOUT(9)
         => \readData6[9]\, A_DOUT(8) => nc118, A_DOUT(7) => 
        \readData6[7]\, A_DOUT(6) => \readData6[6]\, A_DOUT(5)
         => \readData6[5]\, A_DOUT(4) => \readData6[4]\, 
        A_DOUT(3) => \readData6[3]\, A_DOUT(2) => \readData6[2]\, 
        A_DOUT(1) => \readData6[1]\, A_DOUT(0) => \readData6[0]\, 
        B_DOUT(17) => nc106, B_DOUT(16) => \readData6[34]\, 
        B_DOUT(15) => \readData6[33]\, B_DOUT(14) => 
        \readData6[32]\, B_DOUT(13) => \readData6[31]\, 
        B_DOUT(12) => \readData6[30]\, B_DOUT(11) => 
        \readData6[29]\, B_DOUT(10) => \readData6[28]\, B_DOUT(9)
         => \readData6[27]\, B_DOUT(8) => nc75, B_DOUT(7) => 
        \readData6[25]\, B_DOUT(6) => \readData6[24]\, B_DOUT(5)
         => \readData6[23]\, B_DOUT(4) => \readData6[22]\, 
        B_DOUT(3) => \readData6[21]\, B_DOUT(2) => 
        \readData6[20]\, B_DOUT(1) => \readData6[19]\, B_DOUT(0)
         => \readData6[18]\, BUSY => OPEN, A_CLK => FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_21_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a6_1[1]\, 
        A_WEN(0) => \wen_a6_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b6_1[1]\, 
        B_WEN(0) => \wen_b6_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_2[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[27]\, D => \readData3[27]\, Y => 
        \readData_25_1_1[24]\);
    
    \readData_31_am_1_1_RNO_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[7]\, D => \readData4[7]\, Y => 
        \readData_6_1_1[7]\);
    
    \readData_31_am_1_1_RNO_2[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[16]\, D => \readData0[16]\, Y => 
        \readData_3_1_1[15]\);
    
    \readData_31_am_RNO_2[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[0]\, D => \readData2[0]\, Y => 
        \readData_10_1_1[0]\);
    
    \readData_31_bm_RNO_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[24]\, D => \readData7[24]\, Y => 
        \readData_28_1_1[22]\);
    
    \readData_31_am_1_1_RNO_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[16]\, D => \readData4[16]\, Y => 
        \readData_6_1_1[15]\);
    
    \readData_31_bm_1_1_RNO_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[23]\, D => \readData5[23]\, Y => 
        \readData_21_1_1[21]\);
    
    readdata_xhdl1399_0_a2_0 : CFG3
      generic map(INIT => x"10")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1150);
    
    \readData_31_bm_1_1_RNO_0[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[29]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[26]\, D => \readData9[29]\, Y => 
        \readData_31_bm_1_1_RNO_0[26]_net_1\);
    
    \readData_31_am_RNO_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[0]\, D => \readData6[0]\, Y => 
        \readData_13_1_1[0]\);
    
    \readData_31_am_1_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[23]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[23]_net_1\, Y => 
        \readData_31_am_1_1[23]_net_1\);
    
    \readData_31_bm_1_1_RNO[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[2]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[2]\, D => \readData13[2]\, Y => 
        \readData_31_bm_1_1_RNO[2]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[30]\, D => \readData5[30]\, Y => 
        \readData_21_1_1[27]\);
    
    \readData_31_am_RNO[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[30]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[27]\, D => \readData14[30]\, Y => 
        \readData_31_am_RNO[27]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[0]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[0]\, D => \readData9[0]\, Y => 
        \readData_31_bm_1_1_RNO_0[0]_net_1\);
    
    \readData_31_am_1_1_RNO[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[24]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[22]\, D => \readData12[24]\, Y => 
        \readData_31_am_1_1_RNO[22]_net_1\);
    
    \readData_31_am[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[2]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[2]_net_1\, D
         => \readData_31_am_RNO_0[2]_net_1\, Y => 
        \readData_31_am[2]_net_1\);
    
    \readData_31_bm_RNO[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[16]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[15]\, D => \readData15[16]\, Y => 
        \readData_31_bm_RNO[15]_net_1\);
    
    \readData_31_am_RNO_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[24]\, D => \readData6[24]\, Y => 
        \readData_13_1_1[22]\);
    
    \readData_31_bm_RNO_0[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[33]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[30]\, D => \readData11[33]\, Y => 
        \readData_31_bm_RNO_0[30]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    block3_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(0), Y => \wen_a3_1[0]\);
    
    \readData_31_am_RNO[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[29]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[26]\, D => \readData14[29]\, Y => 
        \readData_31_am_RNO[26]_net_1\);
    
    \readData_31_am_RNO[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[6]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[6]\, D => \readData14[6]\, Y => 
        \readData_31_am_RNO[6]_net_1\);
    
    \readData_31_am_RNO[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[34]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[31]\, D => \readData14[34]\, Y => 
        \readData_31_am_RNO[31]_net_1\);
    
    \readData_31_ns[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[4]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[4]_net_1\, Y => 
        ram_rdata(4));
    
    \wen_a_m_10_0_a2_0[1]\ : CFG3
      generic map(INIT => x"04")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1143);
    
    \readData_31_am_1_1_RNO_0[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[24]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[22]\, D => \readData8[24]\, Y => 
        \readData_31_am_1_1_RNO_0[22]_net_1\);
    
    block2_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(1), Y => \wen_a2_1[1]\);
    
    \readData_31_bm_RNO_0[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[9]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[8]\, D => \readData11[9]\, Y => 
        \readData_31_bm_RNO_0[8]_net_1\);
    
    block1_RNO_0 : CFG2
      generic map(INIT => x"8")

      port map(A => sram_wen_mem(1), B => wen_a3133, Y => 
        \wen_a1_1[1]\);
    
    \readData_31_bm_1_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[27]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[27]_net_1\, Y => 
        \readData_31_bm_1_1[27]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[24]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[22]\, D => \readData9[24]\, Y => 
        \readData_31_bm_1_1_RNO_0[22]_net_1\);
    
    \readData_31_am_1_1_RNO_0[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[20]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[18]\, D => \readData8[20]\, Y => 
        \readData_31_am_1_1_RNO_0[18]_net_1\);
    
    \readData_31_am[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[8]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[8]_net_1\, D
         => \readData_31_am_RNO_0[8]_net_1\, Y => 
        \readData_31_am[8]_net_1\);
    
    \readData_31_bm_1_1_RNO[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[4]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[4]\, D => \readData13[4]\, Y => 
        \readData_31_bm_1_1_RNO[4]_net_1\);
    
    block10_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(2), Y => \wen_b10_1[0]\);
    
    \readData_31_bm_1_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[16]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[16]_net_1\, Y => 
        \readData_31_bm_1_1[16]_net_1\);
    
    \readData_31_bm_1_1_RNO[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[15]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[14]\, D => \readData13[15]\, Y => 
        \readData_31_bm_1_1_RNO[14]_net_1\);
    
    \readData_31_am_1_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[8]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[8]_net_1\, Y => 
        \readData_31_am_1_1[8]_net_1\);
    
    \readData_31_ns[13]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[13]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[13]_net_1\, Y => 
        ram_rdata(13));
    
    \readData_31_am_RNO[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[16]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[15]\, D => \readData14[16]\, Y => 
        \readData_31_am_RNO[15]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[29]\, D => \readData1[29]\, Y => 
        \readData_18_1_1[26]\);
    
    \readData_31_bm_RNO_2[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[34]\, D => \readData3[34]\, Y => 
        \readData_25_1_1[31]\);
    
    block4_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(2), Y => \wen_b4_1[0]\);
    
    \readData_31_am_RNO_0[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[29]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[26]\, D => \readData10[29]\, Y => 
        \readData_31_am_RNO_0[26]_net_1\);
    
    \readData_31_bm_RNO[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[23]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[21]\, D => \readData15[23]\, Y => 
        \readData_31_bm_RNO[21]_net_1\);
    
    \readData_31_bm_1_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[24]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[24]_net_1\, Y => 
        \readData_31_bm_1_1[24]_net_1\);
    
    \readData_31_bm_1_1_RNO[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[6]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[6]\, D => \readData13[6]\, Y => 
        \readData_31_bm_1_1_RNO[6]_net_1\);
    
    block11 : RAM1K18
      port map(A_DOUT(17) => nc65, A_DOUT(16) => \readData11[16]\, 
        A_DOUT(15) => \readData11[15]\, A_DOUT(14) => 
        \readData11[14]\, A_DOUT(13) => \readData11[13]\, 
        A_DOUT(12) => \readData11[12]\, A_DOUT(11) => 
        \readData11[11]\, A_DOUT(10) => \readData11[10]\, 
        A_DOUT(9) => \readData11[9]\, A_DOUT(8) => nc38, 
        A_DOUT(7) => \readData11[7]\, A_DOUT(6) => 
        \readData11[6]\, A_DOUT(5) => \readData11[5]\, A_DOUT(4)
         => \readData11[4]\, A_DOUT(3) => \readData11[3]\, 
        A_DOUT(2) => \readData11[2]\, A_DOUT(1) => 
        \readData11[1]\, A_DOUT(0) => \readData11[0]\, B_DOUT(17)
         => nc93, B_DOUT(16) => \readData11[34]\, B_DOUT(15) => 
        \readData11[33]\, B_DOUT(14) => \readData11[32]\, 
        B_DOUT(13) => \readData11[31]\, B_DOUT(12) => 
        \readData11[30]\, B_DOUT(11) => \readData11[29]\, 
        B_DOUT(10) => \readData11[28]\, B_DOUT(9) => 
        \readData11[27]\, B_DOUT(8) => nc1, B_DOUT(7) => 
        \readData11[25]\, B_DOUT(6) => \readData11[24]\, 
        B_DOUT(5) => \readData11[23]\, B_DOUT(4) => 
        \readData11[22]\, B_DOUT(3) => \readData11[21]\, 
        B_DOUT(2) => \readData11[20]\, B_DOUT(1) => 
        \readData11[19]\, B_DOUT(0) => \readData11[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a11_1[1]\, 
        A_WEN(0) => \wen_a11_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b11_1[1]\, 
        B_WEN(0) => \wen_b11_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_RNO_2[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[34]\, D => \readData2[34]\, Y => 
        \readData_10_1_1[31]\);
    
    \readData_31_am_1_1_RNO[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[16]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[15]\, D => \readData12[16]\, Y => 
        \readData_31_am_1_1_RNO[15]_net_1\);
    
    \readData_31_am_RNO_2[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[1]\, D => \readData2[1]\, Y => 
        \readData_10_1_1[1]\);
    
    \readData_31_bm_RNO_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[33]\, D => \readData7[33]\, Y => 
        \readData_28_1_1[30]\);
    
    \readData_31_am_1_1_RNO_2[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[24]\, D => \readData0[24]\, Y => 
        \readData_3_1_1[22]\);
    
    block7_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(3), Y => \wen_b7_1[1]\);
    
    \readData_31_bm_1_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[7]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[7]_net_1\, Y => 
        \readData_31_bm_1_1[7]_net_1\);
    
    block27_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(0), Y => \wen_a27_1[0]\);
    
    \readData_31_bm_1_1_RNO_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[2]\, D => \readData5[2]\, Y => 
        \readData_21_1_1[2]\);
    
    block12 : RAM1K18
      port map(A_DOUT(17) => nc2, A_DOUT(16) => \readData12[16]\, 
        A_DOUT(15) => \readData12[15]\, A_DOUT(14) => 
        \readData12[14]\, A_DOUT(13) => \readData12[13]\, 
        A_DOUT(12) => \readData12[12]\, A_DOUT(11) => 
        \readData12[11]\, A_DOUT(10) => \readData12[10]\, 
        A_DOUT(9) => \readData12[9]\, A_DOUT(8) => nc50, 
        A_DOUT(7) => \readData12[7]\, A_DOUT(6) => 
        \readData12[6]\, A_DOUT(5) => \readData12[5]\, A_DOUT(4)
         => \readData12[4]\, A_DOUT(3) => \readData12[3]\, 
        A_DOUT(2) => \readData12[2]\, A_DOUT(1) => 
        \readData12[1]\, A_DOUT(0) => \readData12[0]\, B_DOUT(17)
         => nc22, B_DOUT(16) => \readData12[34]\, B_DOUT(15) => 
        \readData12[33]\, B_DOUT(14) => \readData12[32]\, 
        B_DOUT(13) => \readData12[31]\, B_DOUT(12) => 
        \readData12[30]\, B_DOUT(11) => \readData12[29]\, 
        B_DOUT(10) => \readData12[28]\, B_DOUT(9) => 
        \readData12[27]\, B_DOUT(8) => nc12, B_DOUT(7) => 
        \readData12[25]\, B_DOUT(6) => \readData12[24]\, 
        B_DOUT(5) => \readData12[23]\, B_DOUT(4) => 
        \readData12[22]\, B_DOUT(3) => \readData12[21]\, 
        B_DOUT(2) => \readData12[20]\, B_DOUT(1) => 
        \readData12[19]\, B_DOUT(0) => \readData12[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a12_1[1]\, 
        A_WEN(0) => \wen_a12_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b12_1[1]\, 
        B_WEN(0) => \wen_b12_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[2]\, D => \readData7[2]\, Y => 
        \readData_28_1_1[2]\);
    
    block26_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(1), Y => \wen_a26_1[1]\);
    
    block12_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(1), Y => \wen_a12_1[1]\);
    
    \readData_31_bm_1_1_RNO_2[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[24]\, D => \readData1[24]\, Y => 
        \readData_18_1_1[22]\);
    
    \readData_31_bm_1_1_RNO[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[34]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[31]\, D => \readData13[34]\, Y => 
        \readData_31_bm_1_1_RNO[31]_net_1\);
    
    \readData_31_bm_RNO_0[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[16]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[15]\, D => \readData11[16]\, Y => 
        \readData_31_bm_RNO_0[15]_net_1\);
    
    \readData_31_bm_RNO[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[29]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[26]\, D => \readData15[29]\, Y => 
        \readData_31_bm_RNO[26]_net_1\);
    
    block13 : RAM1K18
      port map(A_DOUT(17) => nc21, A_DOUT(16) => \readData13[16]\, 
        A_DOUT(15) => \readData13[15]\, A_DOUT(14) => 
        \readData13[14]\, A_DOUT(13) => \readData13[13]\, 
        A_DOUT(12) => \readData13[12]\, A_DOUT(11) => 
        \readData13[11]\, A_DOUT(10) => \readData13[10]\, 
        A_DOUT(9) => \readData13[9]\, A_DOUT(8) => nc11, 
        A_DOUT(7) => \readData13[7]\, A_DOUT(6) => 
        \readData13[6]\, A_DOUT(5) => \readData13[5]\, A_DOUT(4)
         => \readData13[4]\, A_DOUT(3) => \readData13[3]\, 
        A_DOUT(2) => \readData13[2]\, A_DOUT(1) => 
        \readData13[1]\, A_DOUT(0) => \readData13[0]\, B_DOUT(17)
         => nc78, B_DOUT(16) => \readData13[34]\, B_DOUT(15) => 
        \readData13[33]\, B_DOUT(14) => \readData13[32]\, 
        B_DOUT(13) => \readData13[31]\, B_DOUT(12) => 
        \readData13[30]\, B_DOUT(11) => \readData13[29]\, 
        B_DOUT(10) => \readData13[28]\, B_DOUT(9) => 
        \readData13[27]\, B_DOUT(8) => nc54, B_DOUT(7) => 
        \readData13[25]\, B_DOUT(6) => \readData13[24]\, 
        B_DOUT(5) => \readData13[23]\, B_DOUT(4) => 
        \readData13[22]\, B_DOUT(3) => \readData13[21]\, 
        B_DOUT(2) => \readData13[20]\, B_DOUT(1) => 
        \readData13[19]\, B_DOUT(0) => \readData13[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a13_1[1]\, 
        A_WEN(0) => \wen_a13_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b13_1[1]\, 
        B_WEN(0) => \wen_b13_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_RNO_0[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[32]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[29]\, D => \readData10[32]\, Y => 
        \readData_31_am_RNO_0[29]_net_1\);
    
    \readData_31_am_1_1_RNO_0[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[29]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[26]\, D => \readData8[29]\, Y => 
        \readData_31_am_1_1_RNO_0[26]_net_1\);
    
    \readData_31_bm_1_1_RNO[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[27]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[24]\, D => \readData13[27]\, Y => 
        \readData_31_bm_1_1_RNO[24]_net_1\);
    
    \readData_31_bm_RNO[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[22]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[20]\, D => \readData15[22]\, Y => 
        \readData_31_bm_RNO[20]_net_1\);
    
    \readData_31_am_RNO_2[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[18]\, D => \readData2[18]\, Y => 
        \readData_10_1_1[16]\);
    
    \readData_31_bm_1_1_RNO[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[1]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[1]\, D => \readData13[1]\, Y => 
        \readData_31_bm_1_1_RNO[1]_net_1\);
    
    \readData_31_am_RNO_0[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[27]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[24]\, D => \readData10[27]\, Y => 
        \readData_31_am_RNO_0[24]_net_1\);
    
    \readData_31_am_RNO_0[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[2]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[2]\, D => \readData10[2]\, Y => 
        \readData_31_am_RNO_0[2]_net_1\);
    
    \readData_31_am_RNO_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[18]\, D => \readData6[18]\, Y => 
        \readData_13_1_1[16]\);
    
    block0_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem(0), Y => 
        \wen_a0_1[0]\);
    
    \readData_31_bm_1_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[0]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[0]_net_1\, Y => 
        \readData_31_bm_1_1[0]_net_1\);
    
    \readData_31_am_1_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[2]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[2]_net_1\, Y => 
        \readData_31_am_1_1[2]_net_1\);
    
    block24_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(1), Y => \wen_a24_1[1]\);
    
    block18 : RAM1K18
      port map(A_DOUT(17) => nc68, A_DOUT(16) => \readData18[16]\, 
        A_DOUT(15) => \readData18[15]\, A_DOUT(14) => 
        \readData18[14]\, A_DOUT(13) => \readData18[13]\, 
        A_DOUT(12) => \readData18[12]\, A_DOUT(11) => 
        \readData18[11]\, A_DOUT(10) => \readData18[10]\, 
        A_DOUT(9) => \readData18[9]\, A_DOUT(8) => nc3, A_DOUT(7)
         => \readData18[7]\, A_DOUT(6) => \readData18[6]\, 
        A_DOUT(5) => \readData18[5]\, A_DOUT(4) => 
        \readData18[4]\, A_DOUT(3) => \readData18[3]\, A_DOUT(2)
         => \readData18[2]\, A_DOUT(1) => \readData18[1]\, 
        A_DOUT(0) => \readData18[0]\, B_DOUT(17) => nc32, 
        B_DOUT(16) => \readData18[34]\, B_DOUT(15) => 
        \readData18[33]\, B_DOUT(14) => \readData18[32]\, 
        B_DOUT(13) => \readData18[31]\, B_DOUT(12) => 
        \readData18[30]\, B_DOUT(11) => \readData18[29]\, 
        B_DOUT(10) => \readData18[28]\, B_DOUT(9) => 
        \readData18[27]\, B_DOUT(8) => nc104, B_DOUT(7) => 
        \readData18[25]\, B_DOUT(6) => \readData18[24]\, 
        B_DOUT(5) => \readData18[23]\, B_DOUT(4) => 
        \readData18[22]\, B_DOUT(3) => \readData18[21]\, 
        B_DOUT(2) => \readData18[20]\, B_DOUT(1) => 
        \readData18[19]\, B_DOUT(0) => \readData18[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a18_1[1]\, 
        A_WEN(0) => \wen_a18_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b18_1[1]\, 
        B_WEN(0) => \wen_b18_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_1_1_RNO[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[28]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[25]\, D => \readData12[28]\, Y => 
        \readData_31_am_1_1_RNO[25]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[2]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[2]\, D => \readData9[2]\, Y => 
        \readData_31_bm_1_1_RNO_0[2]_net_1\);
    
    \readData_31_am[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[0]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[0]_net_1\, D
         => \readData_31_am_RNO_0[0]_net_1\, Y => 
        \readData_31_am[0]_net_1\);
    
    \readData_31_am_1_1_RNO_0[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[14]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[13]\, D => \readData8[14]\, Y => 
        \readData_31_am_1_1_RNO_0[13]_net_1\);
    
    \readData_31_bm_1_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[15]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[15]_net_1\, Y => 
        \readData_31_bm_1_1[15]_net_1\);
    
    block20_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(1), Y => \wen_a20_1[1]\);
    
    \readData_31_am_RNO_2[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[21]\, D => \readData2[21]\, Y => 
        \readData_10_1_1[19]\);
    
    block18_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(14), C
         => readdata_xhdl1401_1, D => sram_wen_mem(2), Y => 
        \wen_b18_1[0]\);
    
    \readData_31_bm_RNO_2[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[28]\, D => \readData3[28]\, Y => 
        \readData_25_1_1[25]\);
    
    block9_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(3), Y => \wen_b9_1[1]\);
    
    \readData_31_am_1_1_RNO_2[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[33]\, D => \readData0[33]\, Y => 
        \readData_3_1_1[30]\);
    
    \readData_31_ns[10]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[10]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[10]_net_1\, Y => 
        ram_rdata(10));
    
    \readData_31_am_RNO_2[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[15]\, D => \readData2[15]\, Y => 
        \readData_10_1_1[14]\);
    
    \readData_31_am_RNO_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[21]\, D => \readData6[21]\, Y => 
        \readData_13_1_1[19]\);
    
    \readData_31_am_1_1_RNO_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[33]\, D => \readData4[33]\, Y => 
        \readData_6_1_1[30]\);
    
    \readData_31_am[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[16]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[16]_net_1\, D
         => \readData_31_am_RNO_0[16]_net_1\, Y => 
        \readData_31_am[16]_net_1\);
    
    \readData_31_bm_1_1_RNO[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[9]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[8]\, D => \readData13[9]\, Y => 
        \readData_31_bm_1_1_RNO[8]_net_1\);
    
    \readData_31_am[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[19]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[19]_net_1\, D
         => \readData_31_am_RNO_0[19]_net_1\, Y => 
        \readData_31_am[19]_net_1\);
    
    \readData_31_am_1_1_RNO_2[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[29]\, D => \readData0[29]\, Y => 
        \readData_3_1_1[26]\);
    
    \readData_31_am_RNO_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[15]\, D => \readData6[15]\, Y => 
        \readData_13_1_1[14]\);
    
    \readData_31_bm_1_1_RNO_0[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[7]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[7]\, D => \readData9[7]\, Y => 
        \readData_31_bm_1_1_RNO_0[7]_net_1\);
    
    block2 : RAM1K18
      port map(A_DOUT(17) => nc40, A_DOUT(16) => \readData2[16]\, 
        A_DOUT(15) => \readData2[15]\, A_DOUT(14) => 
        \readData2[14]\, A_DOUT(13) => \readData2[13]\, 
        A_DOUT(12) => \readData2[12]\, A_DOUT(11) => 
        \readData2[11]\, A_DOUT(10) => \readData2[10]\, A_DOUT(9)
         => \readData2[9]\, A_DOUT(8) => nc31, A_DOUT(7) => 
        \readData2[7]\, A_DOUT(6) => \readData2[6]\, A_DOUT(5)
         => \readData2[5]\, A_DOUT(4) => \readData2[4]\, 
        A_DOUT(3) => \readData2[3]\, A_DOUT(2) => \readData2[2]\, 
        A_DOUT(1) => \readData2[1]\, A_DOUT(0) => \readData2[0]\, 
        B_DOUT(17) => nc96, B_DOUT(16) => \readData2[34]\, 
        B_DOUT(15) => \readData2[33]\, B_DOUT(14) => 
        \readData2[32]\, B_DOUT(13) => \readData2[31]\, 
        B_DOUT(12) => \readData2[30]\, B_DOUT(11) => 
        \readData2[29]\, B_DOUT(10) => \readData2[28]\, B_DOUT(9)
         => \readData2[27]\, B_DOUT(8) => nc44, B_DOUT(7) => 
        \readData2[25]\, B_DOUT(6) => \readData2[24]\, B_DOUT(5)
         => \readData2[23]\, B_DOUT(4) => \readData2[22]\, 
        B_DOUT(3) => \readData2[21]\, B_DOUT(2) => 
        \readData2[20]\, B_DOUT(1) => \readData2[19]\, B_DOUT(0)
         => \readData2[18]\, BUSY => OPEN, A_CLK => FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_21_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a2_1[1]\, 
        A_WEN(0) => \wen_a2_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b2_1[1]\, 
        B_WEN(0) => \wen_b2_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_RNO_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[9]\, D => \readData6[9]\, Y => 
        \readData_13_1_1[8]\);
    
    \readData_31_bm_1_1_RNO_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[29]\, D => \readData5[29]\, Y => 
        \readData_21_1_1[26]\);
    
    \readData_31_bm_RNO[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[0]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[0]\, D => \readData15[0]\, Y => 
        \readData_31_bm_RNO[0]_net_1\);
    
    block0 : RAM1K18
      port map(A_DOUT(17) => nc7, A_DOUT(16) => \readData0[16]\, 
        A_DOUT(15) => \readData0[15]\, A_DOUT(14) => 
        \readData0[14]\, A_DOUT(13) => \readData0[13]\, 
        A_DOUT(12) => \readData0[12]\, A_DOUT(11) => 
        \readData0[11]\, A_DOUT(10) => \readData0[10]\, A_DOUT(9)
         => \readData0[9]\, A_DOUT(8) => nc97, A_DOUT(7) => 
        \readData0[7]\, A_DOUT(6) => \readData0[6]\, A_DOUT(5)
         => \readData0[5]\, A_DOUT(4) => \readData0[4]\, 
        A_DOUT(3) => \readData0[3]\, A_DOUT(2) => \readData0[2]\, 
        A_DOUT(1) => \readData0[1]\, A_DOUT(0) => \readData0[0]\, 
        B_DOUT(17) => nc85, B_DOUT(16) => \readData0[34]\, 
        B_DOUT(15) => \readData0[33]\, B_DOUT(14) => 
        \readData0[32]\, B_DOUT(13) => \readData0[31]\, 
        B_DOUT(12) => \readData0[30]\, B_DOUT(11) => 
        \readData0[29]\, B_DOUT(10) => \readData0[28]\, B_DOUT(9)
         => \readData0[27]\, B_DOUT(8) => nc72, B_DOUT(7) => 
        \readData0[25]\, B_DOUT(6) => \readData0[24]\, B_DOUT(5)
         => \readData0[23]\, B_DOUT(4) => \readData0[22]\, 
        B_DOUT(3) => \readData0[21]\, B_DOUT(2) => 
        \readData0[20]\, B_DOUT(1) => \readData0[19]\, B_DOUT(0)
         => \readData0[18]\, BUSY => OPEN, A_CLK => FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_21_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a0_1[1]\, 
        A_WEN(0) => \wen_a0_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b0_1[1]\, 
        B_WEN(0) => \wen_b0_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[5]\, D => \readData7[5]\, Y => 
        \readData_28_1_1[5]\);
    
    \readData_31_am[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[7]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[7]_net_1\, D
         => \readData_31_am_RNO_0[7]_net_1\, Y => 
        \readData_31_am[7]_net_1\);
    
    \readData_31_am_RNO_2[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[9]\, D => \readData2[9]\, Y => 
        \readData_10_1_1[8]\);
    
    \readData_31_am_1_1_RNO_2[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[20]\, D => \readData0[20]\, Y => 
        \readData_3_1_1[18]\);
    
    \readData_31_bm_RNO_0[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[29]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[26]\, D => \readData11[29]\, Y => 
        \readData_31_bm_RNO_0[26]_net_1\);
    
    \readData_31_am_1_1_RNO_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[20]\, D => \readData4[20]\, Y => 
        \readData_6_1_1[18]\);
    
    \readData_31_ns[14]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[14]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[14]_net_1\, Y => 
        ram_rdata(14));
    
    \readData_31_bm[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[23]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[23]_net_1\, D
         => \readData_31_bm_RNO_0[23]_net_1\, Y => 
        \readData_31_bm[23]_net_1\);
    
    \readData_31_am_1_1_RNO_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[24]\, D => \readData4[24]\, Y => 
        \readData_6_1_1[22]\);
    
    block28_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(1), Y => \wen_a28_1[1]\);
    
    \readData_31_bm[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[2]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[2]_net_1\, D
         => \readData_31_bm_RNO_0[2]_net_1\, Y => 
        \readData_31_bm[2]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[27]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[24]\, D => \readData9[27]\, Y => 
        \readData_31_bm_1_1_RNO_0[24]_net_1\);
    
    \readData_31_am_1_1_RNO[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[15]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[14]\, D => \readData12[15]\, Y => 
        \readData_31_am_1_1_RNO[14]_net_1\);
    
    \readData_31_bm_RNO_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[23]\, D => \readData7[23]\, Y => 
        \readData_28_1_1[21]\);
    
    \readData_31_bm_RNO_0[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[32]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[29]\, D => \readData11[32]\, Y => 
        \readData_31_bm_RNO_0[29]_net_1\);
    
    \readData_31_am[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[15]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[15]_net_1\, D
         => \readData_31_am_RNO_0[15]_net_1\, Y => 
        \readData_31_am[15]_net_1\);
    
    block29 : RAM1K18
      port map(A_DOUT(17) => nc6, A_DOUT(16) => \readData29[16]\, 
        A_DOUT(15) => \readData29[15]\, A_DOUT(14) => 
        \readData29[14]\, A_DOUT(13) => \readData29[13]\, 
        A_DOUT(12) => \readData29[12]\, A_DOUT(11) => 
        \readData29[11]\, A_DOUT(10) => \readData29[10]\, 
        A_DOUT(9) => \readData29[9]\, A_DOUT(8) => nc71, 
        A_DOUT(7) => \readData29[7]\, A_DOUT(6) => 
        \readData29[6]\, A_DOUT(5) => \readData29[5]\, A_DOUT(4)
         => \readData29[4]\, A_DOUT(3) => \readData29[3]\, 
        A_DOUT(2) => \readData29[2]\, A_DOUT(1) => 
        \readData29[1]\, A_DOUT(0) => \readData29[0]\, B_DOUT(17)
         => nc62, B_DOUT(16) => \readData29[34]\, B_DOUT(15) => 
        \readData29[33]\, B_DOUT(14) => \readData29[32]\, 
        B_DOUT(13) => \readData29[31]\, B_DOUT(12) => 
        \readData29[30]\, B_DOUT(11) => \readData29[29]\, 
        B_DOUT(10) => \readData29[28]\, B_DOUT(9) => 
        \readData29[27]\, B_DOUT(8) => nc61, B_DOUT(7) => 
        \readData29[25]\, B_DOUT(6) => \readData29[24]\, 
        B_DOUT(5) => \readData29[23]\, B_DOUT(4) => 
        \readData29[22]\, B_DOUT(3) => \readData29[21]\, 
        B_DOUT(2) => \readData29[20]\, B_DOUT(1) => 
        \readData29[19]\, B_DOUT(0) => \readData29[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a29_1[1]\, 
        A_WEN(0) => \wen_a29_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b29_1[1]\, 
        B_WEN(0) => \wen_b29_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_1_1_RNO_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[24]\, D => \readData5[24]\, Y => 
        \readData_21_1_1[22]\);
    
    \readData_31_am_RNO_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[23]\, D => \readData6[23]\, Y => 
        \readData_13_1_1[21]\);
    
    block19_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(0), Y => \wen_a19_1[0]\);
    
    \readData_31_ns[26]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[26]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[26]_net_1\, Y => 
        ram_rdata(26));
    
    \readData_31_bm_RNO_2[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[18]\, D => \readData3[18]\, Y => 
        \readData_25_1_1[16]\);
    
    block7 : RAM1K18
      port map(A_DOUT(17) => nc125, A_DOUT(16) => \readData7[16]\, 
        A_DOUT(15) => \readData7[15]\, A_DOUT(14) => 
        \readData7[14]\, A_DOUT(13) => \readData7[13]\, 
        A_DOUT(12) => \readData7[12]\, A_DOUT(11) => 
        \readData7[11]\, A_DOUT(10) => \readData7[10]\, A_DOUT(9)
         => \readData7[9]\, A_DOUT(8) => nc115, A_DOUT(7) => 
        \readData7[7]\, A_DOUT(6) => \readData7[6]\, A_DOUT(5)
         => \readData7[5]\, A_DOUT(4) => \readData7[4]\, 
        A_DOUT(3) => \readData7[3]\, A_DOUT(2) => \readData7[2]\, 
        A_DOUT(1) => \readData7[1]\, A_DOUT(0) => \readData7[0]\, 
        B_DOUT(17) => nc102, B_DOUT(16) => \readData7[34]\, 
        B_DOUT(15) => \readData7[33]\, B_DOUT(14) => 
        \readData7[32]\, B_DOUT(13) => \readData7[31]\, 
        B_DOUT(12) => \readData7[30]\, B_DOUT(11) => 
        \readData7[29]\, B_DOUT(10) => \readData7[28]\, B_DOUT(9)
         => \readData7[27]\, B_DOUT(8) => nc19, B_DOUT(7) => 
        \readData7[25]\, B_DOUT(6) => \readData7[24]\, B_DOUT(5)
         => \readData7[23]\, B_DOUT(4) => \readData7[22]\, 
        B_DOUT(3) => \readData7[21]\, B_DOUT(2) => 
        \readData7[20]\, B_DOUT(1) => \readData7[19]\, B_DOUT(0)
         => \readData7[18]\, BUSY => OPEN, A_CLK => FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_21_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a7_1[1]\, 
        A_WEN(0) => \wen_a7_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b7_1[1]\, 
        B_WEN(0) => \wen_b7_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block25_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(1), Y => \wen_a25_1[1]\);
    
    \readData_31_bm_RNO[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[21]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[19]\, D => \readData15[21]\, Y => 
        \readData_31_bm_RNO[19]_net_1\);
    
    \readData_31_bm[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[8]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[8]_net_1\, D
         => \readData_31_bm_RNO_0[8]_net_1\, Y => 
        \readData_31_bm[8]_net_1\);
    
    block17_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(1), Y => 
        \wen_a17_1[1]\);
    
    \readData_31_am[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[24]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[24]_net_1\, D
         => \readData_31_am_RNO_0[24]_net_1\, Y => 
        \readData_31_am[24]_net_1\);
    
    \readData_31_am_RNO[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[32]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[29]\, D => \readData14[32]\, Y => 
        \readData_31_am_RNO[29]_net_1\);
    
    \readData_31_bm_RNO_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[18]\, D => \readData7[18]\, Y => 
        \readData_28_1_1[16]\);
    
    \readData_31_bm_1_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[5]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[5]_net_1\, Y => 
        \readData_31_bm_1_1[5]_net_1\);
    
    \readData_31_am_1_1_RNO_0[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[22]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[20]\, D => \readData8[22]\, Y => 
        \readData_31_am_1_1_RNO_0[20]_net_1\);
    
    \readData_31_am_1_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[4]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[4]_net_1\, Y => 
        \readData_31_am_1_1[4]_net_1\);
    
    block24 : RAM1K18
      port map(A_DOUT(17) => nc29, A_DOUT(16) => \readData24[16]\, 
        A_DOUT(15) => \readData24[15]\, A_DOUT(14) => 
        \readData24[14]\, A_DOUT(13) => \readData24[13]\, 
        A_DOUT(12) => \readData24[12]\, A_DOUT(11) => 
        \readData24[11]\, A_DOUT(10) => \readData24[10]\, 
        A_DOUT(9) => \readData24[9]\, A_DOUT(8) => nc88, 
        A_DOUT(7) => \readData24[7]\, A_DOUT(6) => 
        \readData24[6]\, A_DOUT(5) => \readData24[5]\, A_DOUT(4)
         => \readData24[4]\, A_DOUT(3) => \readData24[3]\, 
        A_DOUT(2) => \readData24[2]\, A_DOUT(1) => 
        \readData24[1]\, A_DOUT(0) => \readData24[0]\, B_DOUT(17)
         => nc53, B_DOUT(16) => \readData24[34]\, B_DOUT(15) => 
        \readData24[33]\, B_DOUT(14) => \readData24[32]\, 
        B_DOUT(13) => \readData24[31]\, B_DOUT(12) => 
        \readData24[30]\, B_DOUT(11) => \readData24[29]\, 
        B_DOUT(10) => \readData24[28]\, B_DOUT(9) => 
        \readData24[27]\, B_DOUT(8) => nc39, B_DOUT(7) => 
        \readData24[25]\, B_DOUT(6) => \readData24[24]\, 
        B_DOUT(5) => \readData24[23]\, B_DOUT(4) => 
        \readData24[22]\, B_DOUT(3) => \readData24[21]\, 
        B_DOUT(2) => \readData24[20]\, B_DOUT(1) => 
        \readData24[19]\, B_DOUT(0) => \readData24[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a24_1[1]\, 
        A_WEN(0) => \wen_a24_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b24_1[1]\, 
        B_WEN(0) => \wen_b24_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_2[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[21]\, D => \readData3[21]\, Y => 
        \readData_25_1_1[19]\);
    
    \readData_31_bm_1_1_RNO_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[5]\, D => \readData5[5]\, Y => 
        \readData_21_1_1[5]\);
    
    \readData_31_am[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[18]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[18]_net_1\, D
         => \readData_31_am_RNO_0[18]_net_1\, Y => 
        \readData_31_am[18]_net_1\);
    
    \readData_31_bm[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[29]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[29]_net_1\, D
         => \readData_31_bm_RNO_0[29]_net_1\, Y => 
        \readData_31_bm[29]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[0]\, D => \readData1[0]\, Y => 
        \readData_18_1_1[0]\);
    
    \readData_31_am_RNO_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[30]\, D => \readData6[30]\, Y => 
        \readData_13_1_1[27]\);
    
    \readData_31_ns[8]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[8]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[8]_net_1\, Y => 
        ram_rdata(8));
    
    \readData_31_am_1_1_RNO[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[5]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[5]\, D => \readData12[5]\, Y => 
        \readData_31_am_1_1_RNO[5]_net_1\);
    
    block8_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(0), Y => \wen_a8_1[0]\);
    
    \readData_31_bm_RNO_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[21]\, D => \readData7[21]\, Y => 
        \readData_28_1_1[19]\);
    
    \readData_31_ns[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[2]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[2]_net_1\, Y => 
        ram_rdata(2));
    
    \readData_31_bm_1_1_RNO_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[7]\, D => \readData5[7]\, Y => 
        \readData_21_1_1[7]\);
    
    block18_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(14), C
         => readdata_xhdl1401_1, D => sram_wen_mem(0), Y => 
        \wen_a18_1[0]\);
    
    \readData_31_am[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[22]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[22]_net_1\, D
         => \readData_31_am_RNO_0[22]_net_1\, Y => 
        \readData_31_am[22]_net_1\);
    
    \readData_31_bm_RNO_0[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[20]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[18]\, D => \readData11[20]\, Y => 
        \readData_31_bm_RNO_0[18]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[27]\, D => \readData1[27]\, Y => 
        \readData_18_1_1[24]\);
    
    \readData_31_am_1_1_RNO[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[27]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[24]\, D => \readData12[27]\, Y => 
        \readData_31_am_1_1_RNO[24]_net_1\);
    
    \readData_31_am[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_am_RNO[10]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_am_1_1[10]_net_1\, D
         => \readData_31_am_RNO_0[10]_net_1\, Y => 
        \readData_31_am[10]_net_1\);
    
    \readData_31_am_RNO_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[31]\, D => \readData6[31]\, Y => 
        \readData_13_1_1[28]\);
    
    \readData_31_am_RNO_2[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[33]\, D => \readData2[33]\, Y => 
        \readData_10_1_1[30]\);
    
    block25 : RAM1K18
      port map(A_DOUT(17) => nc8, A_DOUT(16) => \readData25[16]\, 
        A_DOUT(15) => \readData25[15]\, A_DOUT(14) => 
        \readData25[14]\, A_DOUT(13) => \readData25[13]\, 
        A_DOUT(12) => \readData25[12]\, A_DOUT(11) => 
        \readData25[11]\, A_DOUT(10) => \readData25[10]\, 
        A_DOUT(9) => \readData25[9]\, A_DOUT(8) => nc82, 
        A_DOUT(7) => \readData25[7]\, A_DOUT(6) => 
        \readData25[6]\, A_DOUT(5) => \readData25[5]\, A_DOUT(4)
         => \readData25[4]\, A_DOUT(3) => \readData25[3]\, 
        A_DOUT(2) => \readData25[2]\, A_DOUT(1) => 
        \readData25[1]\, A_DOUT(0) => \readData25[0]\, B_DOUT(17)
         => nc108, B_DOUT(16) => \readData25[34]\, B_DOUT(15) => 
        \readData25[33]\, B_DOUT(14) => \readData25[32]\, 
        B_DOUT(13) => \readData25[31]\, B_DOUT(12) => 
        \readData25[30]\, B_DOUT(11) => \readData25[29]\, 
        B_DOUT(10) => \readData25[28]\, B_DOUT(9) => 
        \readData25[27]\, B_DOUT(8) => nc81, B_DOUT(7) => 
        \readData25[25]\, B_DOUT(6) => \readData25[24]\, 
        B_DOUT(5) => \readData25[23]\, B_DOUT(4) => 
        \readData25[22]\, B_DOUT(3) => \readData25[21]\, 
        B_DOUT(2) => \readData25[20]\, B_DOUT(1) => 
        \readData25[19]\, B_DOUT(0) => \readData25[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a25_1[1]\, 
        A_WEN(0) => \wen_a25_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b25_1[1]\, 
        B_WEN(0) => \wen_b25_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block1_RNO_1 : CFG4
      generic map(INIT => x"0080")

      port map(A => readdata_xhdl1419_0_a2_0, B => 
        sram_wen_mem(2), C => ahbsram_addr(11), D => 
        ahbsram_addr(15), Y => \wen_b1_1[0]\);
    
    \readData_31_bm_RNO_0[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[25]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[23]\, D => \readData11[25]\, Y => 
        \readData_31_bm_RNO_0[23]_net_1\);
    
    \readData_31_am_1_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[14]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[14]_net_1\, Y => 
        \readData_31_am_1_1[14]_net_1\);
    
    block6_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(0), Y => \wen_a6_1[0]\);
    
    \readData_31_bm_1_1_RNO[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[3]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[3]\, D => \readData13[3]\, Y => 
        \readData_31_bm_1_1_RNO[3]_net_1\);
    
    \readData_31_am_1_1_RNO_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[29]\, D => \readData4[29]\, Y => 
        \readData_6_1_1[26]\);
    
    \readData_31_bm_RNO_0[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[22]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[20]\, D => \readData11[22]\, Y => 
        \readData_31_bm_RNO_0[20]_net_1\);
    
    \readData_31_bm[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[22]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[22]_net_1\, D
         => \readData_31_bm_RNO_0[22]_net_1\, Y => 
        \readData_31_bm[22]_net_1\);
    
    \readData_31_am_1_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[20]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[20]_net_1\, Y => 
        \readData_31_am_1_1[20]_net_1\);
    
    block19_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(1), Y => \wen_a19_1[1]\);
    
    \readData_31_am_1_1_RNO_2[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[14]\, D => \readData0[14]\, Y => 
        \readData_3_1_1[13]\);
    
    block21_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(1), Y => \wen_a21_1[1]\);
    
    block16 : RAM1K18
      port map(A_DOUT(17) => nc79, A_DOUT(16) => \readData16[16]\, 
        A_DOUT(15) => \readData16[15]\, A_DOUT(14) => 
        \readData16[14]\, A_DOUT(13) => \readData16[13]\, 
        A_DOUT(12) => \readData16[12]\, A_DOUT(11) => 
        \readData16[11]\, A_DOUT(10) => \readData16[10]\, 
        A_DOUT(9) => \readData16[9]\, A_DOUT(8) => nc43, 
        A_DOUT(7) => \readData16[7]\, A_DOUT(6) => 
        \readData16[6]\, A_DOUT(5) => \readData16[5]\, A_DOUT(4)
         => \readData16[4]\, A_DOUT(3) => \readData16[3]\, 
        A_DOUT(2) => \readData16[2]\, A_DOUT(1) => 
        \readData16[1]\, A_DOUT(0) => \readData16[0]\, B_DOUT(17)
         => nc69, B_DOUT(16) => \readData16[34]\, B_DOUT(15) => 
        \readData16[33]\, B_DOUT(14) => \readData16[32]\, 
        B_DOUT(13) => \readData16[31]\, B_DOUT(12) => 
        \readData16[30]\, B_DOUT(11) => \readData16[29]\, 
        B_DOUT(10) => \readData16[28]\, B_DOUT(9) => 
        \readData16[27]\, B_DOUT(8) => nc56, B_DOUT(7) => 
        \readData16[25]\, B_DOUT(6) => \readData16[24]\, 
        B_DOUT(5) => \readData16[23]\, B_DOUT(4) => 
        \readData16[22]\, B_DOUT(3) => \readData16[21]\, 
        B_DOUT(2) => \readData16[20]\, B_DOUT(1) => 
        \readData16[19]\, B_DOUT(0) => \readData16[18]\, BUSY => 
        OPEN, A_CLK => FAB_CCC_GL0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_21_i_0, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a16_1[1]\, 
        A_WEN(0) => \wen_a16_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b16_1[1]\, 
        B_WEN(0) => \wen_b16_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_1_1_RNO[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[10]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[9]\, D => \readData13[10]\, Y => 
        \readData_31_bm_1_1_RNO[9]_net_1\);
    
    \readData_31_bm[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[11]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[11]_net_1\, D
         => \readData_31_bm_RNO_0[11]_net_1\, Y => 
        \readData_31_bm[11]_net_1\);
    
    \readData_31_am_1_1_RNO_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[14]\, D => \readData4[14]\, Y => 
        \readData_6_1_1[13]\);
    
    \readData_31_bm_1_1_RNO[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[19]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[17]\, D => \readData13[19]\, Y => 
        \readData_31_bm_1_1_RNO[17]_net_1\);
    
    \readData_31_bm_1_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[23]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[23]_net_1\, Y => 
        \readData_31_bm_1_1[23]_net_1\);
    
    \readData_31_bm_1_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[12]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[12]_net_1\, Y => 
        \readData_31_bm_1_1[12]_net_1\);
    
    \readData_31_am_1_1_RNO_2[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[22]\, D => \readData0[22]\, Y => 
        \readData_3_1_1[20]\);
    
    \readData_31_am_1_1_RNO[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[2]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[2]\, D => \readData12[2]\, Y => 
        \readData_31_am_1_1_RNO[2]_net_1\);
    
    \readData_31_bm_1_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[6]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[6]_net_1\, Y => 
        \readData_31_bm_1_1[6]_net_1\);
    
    block4_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(1), Y => \wen_a4_1[1]\);
    
    block16_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(0), Y => 
        \wen_a16_1[0]\);
    
    \readData_31_bm_RNO_2[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[31]\, D => \readData3[31]\, Y => 
        \readData_25_1_1[28]\);
    
    \readData_31_bm_RNO_2[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[14]\, D => \readData3[14]\, Y => 
        \readData_25_1_1[13]\);
    
    \readData_31_bm[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[30]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[30]_net_1\, D
         => \readData_31_bm_RNO_0[30]_net_1\, Y => 
        \readData_31_bm[30]_net_1\);
    
    block9 : RAM1K18
      port map(A_DOUT(17) => nc20, A_DOUT(16) => \readData9[16]\, 
        A_DOUT(15) => \readData9[15]\, A_DOUT(14) => 
        \readData9[14]\, A_DOUT(13) => \readData9[13]\, 
        A_DOUT(12) => \readData9[12]\, A_DOUT(11) => 
        \readData9[11]\, A_DOUT(10) => \readData9[10]\, A_DOUT(9)
         => \readData9[9]\, A_DOUT(8) => nc10, A_DOUT(7) => 
        \readData9[7]\, A_DOUT(6) => \readData9[6]\, A_DOUT(5)
         => \readData9[5]\, A_DOUT(4) => \readData9[4]\, 
        A_DOUT(3) => \readData9[3]\, A_DOUT(2) => \readData9[2]\, 
        A_DOUT(1) => \readData9[1]\, A_DOUT(0) => \readData9[0]\, 
        B_DOUT(17) => nc57, B_DOUT(16) => \readData9[34]\, 
        B_DOUT(15) => \readData9[33]\, B_DOUT(14) => 
        \readData9[32]\, B_DOUT(13) => \readData9[31]\, 
        B_DOUT(12) => \readData9[30]\, B_DOUT(11) => 
        \readData9[29]\, B_DOUT(10) => \readData9[28]\, B_DOUT(9)
         => \readData9[27]\, B_DOUT(8) => nc95, B_DOUT(7) => 
        \readData9[25]\, B_DOUT(6) => \readData9[24]\, B_DOUT(5)
         => \readData9[23]\, B_DOUT(4) => \readData9[22]\, 
        B_DOUT(3) => \readData9[21]\, B_DOUT(2) => 
        \readData9[20]\, B_DOUT(1) => \readData9[19]\, B_DOUT(0)
         => \readData9[18]\, BUSY => OPEN, A_CLK => FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_21_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a9_1[1]\, 
        A_WEN(0) => \wen_a9_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b9_1[1]\, 
        B_WEN(0) => \wen_b9_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_2[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[11]\, D => \readData3[11]\, Y => 
        \readData_25_1_1[10]\);
    
    \readData_31_am_1_1_RNO_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[4]\, D => \readData4[4]\, Y => 
        \readData_6_1_1[4]\);
    
    \readData_31_am_RNO_0[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[5]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[5]\, D => \readData10[5]\, Y => 
        \readData_31_am_RNO_0[5]_net_1\);
    
    \readData_31_am_1_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[27]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[27]_net_1\, Y => 
        \readData_31_am_1_1[27]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[14]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[13]\, D => \readData9[14]\, Y => 
        \readData_31_bm_1_1_RNO_0[13]_net_1\);
    
    \readData_31_bm_RNO_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[14]\, D => \readData7[14]\, Y => 
        \readData_28_1_1[13]\);
    
    block17_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(3), Y => 
        \wen_b17_1[1]\);
    
    \readData_31_bm_RNO_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[4]\, D => \readData7[4]\, Y => 
        \readData_28_1_1[4]\);
    
    \readData_31_am_1_1_RNO_0[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[34]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[31]\, D => \readData8[34]\, Y => 
        \readData_31_am_1_1_RNO_0[31]_net_1\);
    
    block21_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(3), Y => \wen_b_m[1]\);
    
    \readData_31_am_1_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[30]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[30]_net_1\, Y => 
        \readData_31_am_1_1[30]_net_1\);
    
    \readData_31_bm_RNO_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[11]\, D => \readData7[11]\, Y => 
        \readData_28_1_1[10]\);
    
    \readData_31_am_1_1_RNO_0[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[6]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[6]\, D => \readData8[6]\, Y => 
        \readData_31_am_1_1_RNO_0[6]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[33]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[30]\, D => \readData9[33]\, Y => 
        \readData_31_bm_1_1_RNO_0[30]_net_1\);
    
    \readData_31_bm[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[0]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[0]_net_1\, D
         => \readData_31_bm_RNO_0[0]_net_1\, Y => 
        \readData_31_bm[0]_net_1\);
    
    \readData_31_bm_RNO_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[6]\, D => \readData7[6]\, Y => 
        \readData_28_1_1[6]\);
    
    \readData_31_am_1_1_RNO[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[4]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[4]\, D => \readData12[4]\, Y => 
        \readData_31_am_1_1_RNO[4]_net_1\);
    
    block17_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(2), Y => 
        \wen_b17_1[0]\);
    
    \readData_31_bm_RNO_0[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[7]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[7]\, D => \readData11[7]\, Y => 
        \readData_31_bm_RNO_0[7]_net_1\);
    
    \readData_31_bm_1_1_RNO[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[30]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[27]\, D => \readData13[30]\, Y => 
        \readData_31_bm_1_1_RNO[27]_net_1\);
    
    \readData_31_am_1_1_RNO_0[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[21]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[19]\, D => \readData8[21]\, Y => 
        \readData_31_am_1_1_RNO_0[19]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[34]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[31]\, D => \readData9[34]\, Y => 
        \readData_31_bm_1_1_RNO_0[31]_net_1\);
    
    \readData_31_am_1_1_RNO[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[6]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[6]\, D => \readData12[6]\, Y => 
        \readData_31_am_1_1_RNO[6]_net_1\);
    
    block30_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(3), Y => \wen_b30_1[1]\);
    
    \readData_31_bm_1_1_RNO[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[33]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[30]\, D => \readData13[33]\, Y => 
        \readData_31_bm_1_1_RNO[30]_net_1\);
    
    block3 : RAM1K18
      port map(A_DOUT(17) => nc24, A_DOUT(16) => \readData3[16]\, 
        A_DOUT(15) => \readData3[15]\, A_DOUT(14) => 
        \readData3[14]\, A_DOUT(13) => \readData3[13]\, 
        A_DOUT(12) => \readData3[12]\, A_DOUT(11) => 
        \readData3[11]\, A_DOUT(10) => \readData3[10]\, A_DOUT(9)
         => \readData3[9]\, A_DOUT(8) => nc14, A_DOUT(7) => 
        \readData3[7]\, A_DOUT(6) => \readData3[6]\, A_DOUT(5)
         => \readData3[5]\, A_DOUT(4) => \readData3[4]\, 
        A_DOUT(3) => \readData3[3]\, A_DOUT(2) => \readData3[2]\, 
        A_DOUT(1) => \readData3[1]\, A_DOUT(0) => \readData3[0]\, 
        B_DOUT(17) => nc46, B_DOUT(16) => \readData3[34]\, 
        B_DOUT(15) => \readData3[33]\, B_DOUT(14) => 
        \readData3[32]\, B_DOUT(13) => \readData3[31]\, 
        B_DOUT(12) => \readData3[30]\, B_DOUT(11) => 
        \readData3[29]\, B_DOUT(10) => \readData3[28]\, B_DOUT(9)
         => \readData3[27]\, B_DOUT(8) => nc30, B_DOUT(7) => 
        \readData3[25]\, B_DOUT(6) => \readData3[24]\, B_DOUT(5)
         => \readData3[23]\, B_DOUT(4) => \readData3[22]\, 
        B_DOUT(3) => \readData3[21]\, B_DOUT(2) => 
        \readData3[20]\, B_DOUT(1) => \readData3[19]\, B_DOUT(0)
         => \readData3[18]\, BUSY => OPEN, A_CLK => FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_21_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), A_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), A_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), A_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), A_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), A_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), A_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), A_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), A_DIN(8) => GND_net_1, 
        A_DIN(7) => CoreAHBLite_0_AHBmslave3_HWDATA(7), A_DIN(6)
         => CoreAHBLite_0_AHBmslave3_HWDATA(6), A_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), A_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), A_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), A_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), A_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), A_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a3_1[1]\, 
        A_WEN(0) => \wen_a3_1[0]\, B_CLK => FAB_CCC_GL0, 
        B_DOUT_CLK => VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN
         => VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => 
        VCC_net_1, B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => 
        VCC_net_1, B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => 
        GND_net_1, B_DIN(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), B_DIN(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), B_DIN(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), B_DIN(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), B_DIN(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), B_DIN(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), B_DIN(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), B_DIN(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), B_DIN(8) => 
        GND_net_1, B_DIN(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), B_DIN(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), B_DIN(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), B_DIN(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), B_DIN(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), B_DIN(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), B_DIN(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), B_DIN(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b3_1[1]\, 
        B_WEN(0) => \wen_b3_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_ns[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[0]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[0]_net_1\, Y => 
        ram_rdata(0));
    
    \readData_31_am_1_1_RNO[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[34]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[31]\, D => \readData12[34]\, Y => 
        \readData_31_am_1_1_RNO[31]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[21]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[19]\, D => \readData9[21]\, Y => 
        \readData_31_bm_1_1_RNO_0[19]_net_1\);
    
    \readData_31_bm[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData_31_bm_RNO[7]_net_1\, B => 
        ahbsram_addr(12), C => \readData_31_bm_1_1[7]_net_1\, D
         => \readData_31_bm_RNO_0[7]_net_1\, Y => 
        \readData_31_bm[7]_net_1\);
    
    \readData_31_am_RNO_2[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[2]\, D => \readData2[2]\, Y => 
        \readData_10_1_1[2]\);
    
    \readData_31_bm_1_1_RNO_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[27]\, D => \readData5[27]\, Y => 
        \readData_21_1_1[24]\);
    
    \readData_31_bm_RNO[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[15]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[14]\, D => \readData15[15]\, Y => 
        \readData_31_bm_RNO[14]_net_1\);
    
    \readData_31_am_RNO_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[10]\, D => \readData6[10]\, Y => 
        \readData_13_1_1[9]\);
    
    \readData_31_bm_1_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[18]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[18]_net_1\, Y => 
        \readData_31_bm_1_1[18]_net_1\);
    
    \readData_31_am_1_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_am_1_1_RNO[3]_net_1\, D => 
        \readData_31_am_1_1_RNO_0[3]_net_1\, Y => 
        \readData_31_am_1_1[3]_net_1\);
    
    \readData_31_am_1_1_RNO_2[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[9]\, D => \readData0[9]\, Y => 
        \readData_3_1_1[8]\);
    
    \readData_31_am_1_1_RNO_0[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[27]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[24]\, D => \readData8[27]\, Y => 
        \readData_31_am_1_1_RNO_0[24]_net_1\);
    
    \readData_31_bm_1_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => \readData_31_bm_1_1_RNO[26]_net_1\, D => 
        \readData_31_bm_1_1_RNO_0[26]_net_1\, Y => 
        \readData_31_bm_1_1[26]_net_1\);
    
    \wen_a_m_12_0_a2_0[1]\ : CFG3
      generic map(INIT => x"08")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1147);
    
    block29_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(0), Y => \wen_a29_1[0]\);
    
    block3_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(2), Y => \wen_b3_1[0]\);
    
    \readData_31_ns[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[3]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[3]_net_1\, Y => 
        ram_rdata(3));
    
    \readData_31_am_1_1_RNO_0[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[28]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[25]\, D => \readData8[28]\, Y => 
        \readData_31_am_1_1_RNO_0[25]_net_1\);
    
    \readData_31_am_1_1_RNO[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[1]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[1]\, D => \readData12[1]\, Y => 
        \readData_31_am_1_1_RNO[1]_net_1\);
    
    \readData_31_am_RNO[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[20]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[18]\, D => \readData14[20]\, Y => 
        \readData_31_am_RNO[18]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf is

    port( CoreAHBLite_0_AHBmslave3_HRDATA : out   std_logic_vector(31 downto 0);
          sramcurr_state                  : out   std_logic_vector(1 downto 0);
          ahbsram_size                    : in    std_logic_vector(1 downto 0);
          ahbcurr_state                   : in    std_logic_vector(1 downto 0);
          ahbsram_addr                    : in    std_logic_vector(15 downto 0);
          CoreAHBLite_0_AHBmslave3_HWDATA : in    std_logic_vector(31 downto 0);
          MSS_READY                       : in    std_logic;
          FAB_CCC_GL0                     : in    std_logic;
          sram_done                       : out   std_logic;
          ahbsram_req_d1                  : in    std_logic;
          HWRITE_d                        : in    std_logic
        );

end CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf;

architecture DEF_ARCH of 
        CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component 
        CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8
    port( ram_rdata                       : out   std_logic_vector(31 downto 0);
          sram_wen_mem                    : in    std_logic_vector(3 downto 0) := (others => 'U');
          ahbsram_addr                    : in    std_logic_vector(15 downto 2) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HWDATA : in    std_logic_vector(31 downto 0) := (others => 'U');
          FAB_CCC_GL0                     : in    std_logic := 'U';
          MSS_READY                       : in    std_logic := 'U';
          N_21_i_0                        : in    std_logic := 'U'
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \ram_rdata[20]\, \sram_ren_d\, GND_net_1, 
        \ram_rdata[21]\, \ram_rdata[22]\, \ram_rdata[23]\, 
        \ram_rdata[24]\, \ram_rdata[25]\, \ram_rdata[26]\, 
        \ram_rdata[27]\, \ram_rdata[28]\, \ram_rdata[29]\, 
        \ram_rdata[30]\, \ram_rdata[31]\, \ram_rdata[5]\, 
        \ram_rdata[6]\, \ram_rdata[7]\, \ram_rdata[8]\, 
        \ram_rdata[9]\, \ram_rdata[10]\, \ram_rdata[11]\, 
        \ram_rdata[12]\, \ram_rdata[13]\, \ram_rdata[14]\, 
        \ram_rdata[15]\, \ram_rdata[16]\, \ram_rdata[17]\, 
        \ram_rdata[18]\, \ram_rdata[19]\, \ram_rdata[0]\, 
        \ram_rdata[1]\, \ram_rdata[2]\, \ram_rdata[3]\, 
        \ram_rdata[4]\, \sramcurr_state[0]_net_1\, N_20_i_0, 
        \sramcurr_state[1]_net_1\, N_44_i_0, sram_done_net_1, 
        N_50_i_0, N_21_i_0, N_121, N_116, N_83, N_104, N_96, 
        N_107, \sram_wen_mem[0]_net_1\, \sram_wen_mem[1]_net_1\, 
        \sram_wen_mem[2]\, \sram_wen_mem[3]\ : std_logic;

    for all : CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8
	Use entity work.
        CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8(DEF_ARCH);
begin 

    sramcurr_state(1) <= \sramcurr_state[1]_net_1\;
    sramcurr_state(0) <= \sramcurr_state[0]_net_1\;
    sram_done <= sram_done_net_1;

    \sramahb_rdata_xhdl2[25]\ : SLE
      port map(D => \ram_rdata[25]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(25));
    
    \sramahb_rdata_xhdl2[16]\ : SLE
      port map(D => \ram_rdata[16]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(16));
    
    \sramahb_rdata_xhdl2[24]\ : SLE
      port map(D => \ram_rdata[24]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(24));
    
    \sram_wen_mem_m3[3]\ : CFG4
      generic map(INIT => x"080F")

      port map(A => ahbsram_addr(1), B => ahbsram_addr(0), C => 
        N_96, D => N_116, Y => \sram_wen_mem[3]\);
    
    \sramahb_rdata_xhdl2[8]\ : SLE
      port map(D => \ram_rdata[8]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(8));
    
    \sramahb_rdata_xhdl2[13]\ : SLE
      port map(D => \ram_rdata[13]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(13));
    
    sram_ren_1_sqmuxa_0_a2_i_o3_RNIK3121 : CFG3
      generic map(INIT => x"01")

      port map(A => \sramcurr_state[0]_net_1\, B => N_104, C => 
        \sramcurr_state[1]_net_1\, Y => N_21_i_0);
    
    \sramahb_rdata_xhdl2[9]\ : SLE
      port map(D => \ram_rdata[9]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(9));
    
    \sramcurr_state_ns_1_0_.m4_i_m4\ : CFG4
      generic map(INIT => x"303A")

      port map(A => HWRITE_d, B => sram_done_net_1, C => 
        \sramcurr_state[0]_net_1\, D => N_83, Y => N_107);
    
    \sramahb_rdata_xhdl2[2]\ : SLE
      port map(D => \ram_rdata[2]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(2));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sramahb_rdata_xhdl2[22]\ : SLE
      port map(D => \ram_rdata[22]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(22));
    
    \sram_wen_mem[0]\ : CFG4
      generic map(INIT => x"010F")

      port map(A => ahbsram_addr(1), B => ahbsram_addr(0), C => 
        N_96, D => N_121, Y => \sram_wen_mem[0]_net_1\);
    
    \sramahb_rdata_xhdl2[5]\ : SLE
      port map(D => \ram_rdata[5]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(5));
    
    \sramahb_rdata_xhdl2[19]\ : SLE
      port map(D => \ram_rdata[19]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(19));
    
    \sramahb_rdata_xhdl2[4]\ : SLE
      port map(D => \ram_rdata[4]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(4));
    
    \sramahb_rdata_xhdl2[21]\ : SLE
      port map(D => \ram_rdata[21]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(21));
    
    \sramahb_rdata_xhdl2[18]\ : SLE
      port map(D => \ram_rdata[18]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(18));
    
    \sramahb_rdata_xhdl2[20]\ : SLE
      port map(D => \ram_rdata[20]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(20));
    
    \sramahb_rdata_xhdl2[15]\ : SLE
      port map(D => \ram_rdata[15]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(15));
    
    \sramcurr_state[0]\ : SLE
      port map(D => N_20_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sramcurr_state[0]_net_1\);
    
    \sramahb_rdata_xhdl2[14]\ : SLE
      port map(D => \ram_rdata[14]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(14));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sram_done\ : SLE
      port map(D => N_50_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => sram_done_net_1);
    
    \sramahb_rdata_xhdl2[0]\ : SLE
      port map(D => \ram_rdata[0]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(0));
    
    sram_done_RNO : CFG3
      generic map(INIT => x"01")

      port map(A => \sramcurr_state[0]_net_1\, B => N_83, C => 
        \sramcurr_state[1]_net_1\, Y => N_50_i_0);
    
    \sram_wen_mem_m3[2]\ : CFG4
      generic map(INIT => x"020F")

      port map(A => ahbsram_addr(1), B => ahbsram_addr(0), C => 
        N_96, D => N_116, Y => \sram_wen_mem[2]\);
    
    \sramahb_rdata_xhdl2[27]\ : SLE
      port map(D => \ram_rdata[27]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(27));
    
    \S0.byte_0\ : 
        CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8
      port map(ram_rdata(31) => \ram_rdata[31]\, ram_rdata(30)
         => \ram_rdata[30]\, ram_rdata(29) => \ram_rdata[29]\, 
        ram_rdata(28) => \ram_rdata[28]\, ram_rdata(27) => 
        \ram_rdata[27]\, ram_rdata(26) => \ram_rdata[26]\, 
        ram_rdata(25) => \ram_rdata[25]\, ram_rdata(24) => 
        \ram_rdata[24]\, ram_rdata(23) => \ram_rdata[23]\, 
        ram_rdata(22) => \ram_rdata[22]\, ram_rdata(21) => 
        \ram_rdata[21]\, ram_rdata(20) => \ram_rdata[20]\, 
        ram_rdata(19) => \ram_rdata[19]\, ram_rdata(18) => 
        \ram_rdata[18]\, ram_rdata(17) => \ram_rdata[17]\, 
        ram_rdata(16) => \ram_rdata[16]\, ram_rdata(15) => 
        \ram_rdata[15]\, ram_rdata(14) => \ram_rdata[14]\, 
        ram_rdata(13) => \ram_rdata[13]\, ram_rdata(12) => 
        \ram_rdata[12]\, ram_rdata(11) => \ram_rdata[11]\, 
        ram_rdata(10) => \ram_rdata[10]\, ram_rdata(9) => 
        \ram_rdata[9]\, ram_rdata(8) => \ram_rdata[8]\, 
        ram_rdata(7) => \ram_rdata[7]\, ram_rdata(6) => 
        \ram_rdata[6]\, ram_rdata(5) => \ram_rdata[5]\, 
        ram_rdata(4) => \ram_rdata[4]\, ram_rdata(3) => 
        \ram_rdata[3]\, ram_rdata(2) => \ram_rdata[2]\, 
        ram_rdata(1) => \ram_rdata[1]\, ram_rdata(0) => 
        \ram_rdata[0]\, sram_wen_mem(3) => \sram_wen_mem[3]\, 
        sram_wen_mem(2) => \sram_wen_mem[2]\, sram_wen_mem(1) => 
        \sram_wen_mem[1]_net_1\, sram_wen_mem(0) => 
        \sram_wen_mem[0]_net_1\, ahbsram_addr(15) => 
        ahbsram_addr(15), ahbsram_addr(14) => ahbsram_addr(14), 
        ahbsram_addr(13) => ahbsram_addr(13), ahbsram_addr(12)
         => ahbsram_addr(12), ahbsram_addr(11) => 
        ahbsram_addr(11), ahbsram_addr(10) => ahbsram_addr(10), 
        ahbsram_addr(9) => ahbsram_addr(9), ahbsram_addr(8) => 
        ahbsram_addr(8), ahbsram_addr(7) => ahbsram_addr(7), 
        ahbsram_addr(6) => ahbsram_addr(6), ahbsram_addr(5) => 
        ahbsram_addr(5), ahbsram_addr(4) => ahbsram_addr(4), 
        ahbsram_addr(3) => ahbsram_addr(3), ahbsram_addr(2) => 
        ahbsram_addr(2), CoreAHBLite_0_AHBmslave3_HWDATA(31) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), 
        CoreAHBLite_0_AHBmslave3_HWDATA(30) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), 
        CoreAHBLite_0_AHBmslave3_HWDATA(29) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), 
        CoreAHBLite_0_AHBmslave3_HWDATA(28) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), 
        CoreAHBLite_0_AHBmslave3_HWDATA(27) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), 
        CoreAHBLite_0_AHBmslave3_HWDATA(26) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), 
        CoreAHBLite_0_AHBmslave3_HWDATA(25) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), 
        CoreAHBLite_0_AHBmslave3_HWDATA(24) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), 
        CoreAHBLite_0_AHBmslave3_HWDATA(23) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), 
        CoreAHBLite_0_AHBmslave3_HWDATA(22) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), 
        CoreAHBLite_0_AHBmslave3_HWDATA(21) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), 
        CoreAHBLite_0_AHBmslave3_HWDATA(20) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), 
        CoreAHBLite_0_AHBmslave3_HWDATA(19) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), 
        CoreAHBLite_0_AHBmslave3_HWDATA(18) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), 
        CoreAHBLite_0_AHBmslave3_HWDATA(17) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), 
        CoreAHBLite_0_AHBmslave3_HWDATA(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), 
        CoreAHBLite_0_AHBmslave3_HWDATA(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), 
        CoreAHBLite_0_AHBmslave3_HWDATA(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), 
        CoreAHBLite_0_AHBmslave3_HWDATA(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), 
        CoreAHBLite_0_AHBmslave3_HWDATA(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), 
        CoreAHBLite_0_AHBmslave3_HWDATA(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), 
        CoreAHBLite_0_AHBmslave3_HWDATA(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), 
        CoreAHBLite_0_AHBmslave3_HWDATA(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), 
        CoreAHBLite_0_AHBmslave3_HWDATA(8) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), 
        CoreAHBLite_0_AHBmslave3_HWDATA(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(7), 
        CoreAHBLite_0_AHBmslave3_HWDATA(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(6), 
        CoreAHBLite_0_AHBmslave3_HWDATA(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), 
        CoreAHBLite_0_AHBmslave3_HWDATA(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), 
        CoreAHBLite_0_AHBmslave3_HWDATA(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), 
        CoreAHBLite_0_AHBmslave3_HWDATA(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), 
        CoreAHBLite_0_AHBmslave3_HWDATA(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), 
        CoreAHBLite_0_AHBmslave3_HWDATA(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), FAB_CCC_GL0 => 
        FAB_CCC_GL0, MSS_READY => MSS_READY, N_21_i_0 => N_21_i_0);
    
    sram_wen_mems2_i_a3 : CFG3
      generic map(INIT => x"51")

      port map(A => ahbsram_size(1), B => ahbsram_size(0), C => 
        ahbsram_addr(1), Y => N_121);
    
    \sramahb_rdata_xhdl2[26]\ : SLE
      port map(D => \ram_rdata[26]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(26));
    
    \sramcurr_state_ns_1_0_.N_20_i\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_107, B => \sramcurr_state[1]_net_1\, Y => 
        N_20_i_0);
    
    \sram_wen_mem_m3_i_o3[0]\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => HWRITE_d, B => \sramcurr_state[1]_net_1\, C
         => \sramcurr_state[0]_net_1\, D => N_83, Y => N_96);
    
    \sramahb_rdata_xhdl2[12]\ : SLE
      port map(D => \ram_rdata[12]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(12));
    
    \sramahb_rdata_xhdl2[31]\ : SLE
      port map(D => \ram_rdata[31]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(31));
    
    \sramahb_rdata_xhdl2[23]\ : SLE
      port map(D => \ram_rdata[23]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(23));
    
    \sramahb_rdata_xhdl2[30]\ : SLE
      port map(D => \ram_rdata[30]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(30));
    
    \sram_wen_mem[1]\ : CFG4
      generic map(INIT => x"040F")

      port map(A => ahbsram_addr(1), B => ahbsram_addr(0), C => 
        N_96, D => N_121, Y => \sram_wen_mem[1]_net_1\);
    
    sram_ren_d : SLE
      port map(D => N_21_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sram_ren_d\);
    
    sram_ren_1_sqmuxa_0_a2_i_o3 : CFG2
      generic map(INIT => x"E")

      port map(A => N_83, B => HWRITE_d, Y => N_104);
    
    \sramahb_rdata_xhdl2[11]\ : SLE
      port map(D => \ram_rdata[11]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(11));
    
    \sramcurr_state_ns_1_0_.N_44_i\ : CFG4
      generic map(INIT => x"0407")

      port map(A => sram_done_net_1, B => 
        \sramcurr_state[1]_net_1\, C => \sramcurr_state[0]_net_1\, 
        D => N_104, Y => N_44_i_0);
    
    \sramahb_rdata_xhdl2[10]\ : SLE
      port map(D => \ram_rdata[10]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(10));
    
    \sramcurr_state[1]\ : SLE
      port map(D => N_44_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sramcurr_state[1]_net_1\);
    
    \sramahb_rdata_xhdl2[6]\ : SLE
      port map(D => \ram_rdata[6]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(6));
    
    \sramahb_rdata_xhdl2[7]\ : SLE
      port map(D => \ram_rdata[7]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(7));
    
    \sramahb_rdata_xhdl2[1]\ : SLE
      port map(D => \ram_rdata[1]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(1));
    
    sram_wen_mem_ss3_i_0_a3 : CFG3
      generic map(INIT => x"15")

      port map(A => ahbsram_size(1), B => ahbsram_size(0), C => 
        ahbsram_addr(1), Y => N_116);
    
    \sramahb_rdata_xhdl2[29]\ : SLE
      port map(D => \ram_rdata[29]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(29));
    
    \sramahb_rdata_xhdl2[28]\ : SLE
      port map(D => \ram_rdata[28]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(28));
    
    \sramahb_rdata_xhdl2[17]\ : SLE
      port map(D => \ram_rdata[17]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(17));
    
    sram_ren_0_sqmuxa_0_a2_i_o3 : CFG3
      generic map(INIT => x"AB")

      port map(A => ahbsram_req_d1, B => ahbcurr_state(1), C => 
        ahbcurr_state(0), Y => N_83);
    
    \sramahb_rdata_xhdl2[3]\ : SLE
      port map(D => \ram_rdata[3]\, CLK => FAB_CCC_GL0, EN => 
        \sram_ren_d\, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf is

    port( ahbsram_size                            : out   std_logic_vector(1 downto 0);
          M0GATEDHSIZE                            : in    std_logic_vector(1 downto 0);
          ahbsram_addr                            : out   std_logic_vector(15 downto 0);
          M0GATEDHADDR                            : in    std_logic_vector(15 downto 0);
          ahbcurr_state                           : out   std_logic_vector(1 downto 0);
          MASTERADDRINPROG_i_a2_0_a3_0            : in    std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_d_d          : in    std_logic_vector(0 to 0);
          sramcurr_state                          : in    std_logic_vector(1 downto 0);
          MSS_READY                               : in    std_logic;
          FAB_CCC_GL0                             : in    std_logic;
          N_25_i_0                                : in    std_logic;
          HWRITE_d                                : out   std_logic;
          N_7_i_0                                 : in    std_logic;
          ahbsram_req_d1                          : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1     : out   std_logic;
          M0GATEDHWRITE                           : in    std_logic;
          defSlaveSMNextState_m                   : in    std_logic;
          sram_done                               : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3         : in    std_logic;
          defSlaveSMCurrentState                  : in    std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_2         : in    std_logic
        );

end CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf;

architecture DEF_ARCH of 
        CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \count[3]_net_1\, VCC_net_1, N_94_i_0, counte, 
        GND_net_1, \count[4]_net_1\, N_103_i_i_0, 
        \count[1]_net_1\, N_5_i_0, \count[2]_net_1\, N_93_i_0, 
        \count[0]_net_1\, N_119, \burst_count_reg[0]_net_1\, 
        N_24_i_0, \ahbcurr_state[1]_net_1\, N_23_i_0, 
        \ahbcurr_state[0]_net_1\, \ahbcurr_state_ns[0]\, 
        ahbsram_req_d1_net_1, 
        \CoreAHBLite_0_AHBmslave3_HREADY_i_1\, N_23_i_1, 
        m9_i_a3_1_0, m9_i_a3_0_0, m6_0_a2_4_0, N_78_i, N_85, 
        N_126, m6_0_a3_0, m6_0_a2_1, un1_sramahb_ack_i_i_0, N_80, 
        N_131, N_151, m6_0_a3_2 : std_logic;

begin 

    ahbcurr_state(1) <= \ahbcurr_state[1]_net_1\;
    ahbcurr_state(0) <= \ahbcurr_state[0]_net_1\;
    ahbsram_req_d1 <= ahbsram_req_d1_net_1;
    CoreAHBLite_0_AHBmslave3_HREADY_i_1 <= 
        \CoreAHBLite_0_AHBmslave3_HREADY_i_1\;

    \HWRITE_d\ : SLE
      port map(D => N_7_i_0, CLK => FAB_CCC_GL0, EN => N_25_i_0, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => HWRITE_d);
    
    \count[1]\ : SLE
      port map(D => N_5_i_0, CLK => FAB_CCC_GL0, EN => counte, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \count[1]_net_1\);
    
    \HADDR_d[1]\ : SLE
      port map(D => M0GATEDHADDR(1), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(1));
    
    \HADDR_d[15]\ : SLE
      port map(D => M0GATEDHADDR(15), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(15));
    
    \count[0]\ : SLE
      port map(D => N_119, CLK => FAB_CCC_GL0, EN => counte, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \count[0]_net_1\);
    
    \ahbcurr_state_ns_1_0_.m6_0_a3_2\ : CFG4
      generic map(INIT => x"C0C4")

      port map(A => un1_hready_m_xhdl342_1_i_0_o3_3, B => 
        m6_0_a3_0, C => defSlaveSMCurrentState, D => 
        un1_hready_m_xhdl342_1_i_0_o3_2, Y => m6_0_a3_2);
    
    \ahbcurr_state_ns_1_0_.m6_0_a3_0\ : CFG3
      generic map(INIT => x"04")

      port map(A => \ahbcurr_state[0]_net_1\, B => M0GATEDHWRITE, 
        C => \ahbcurr_state[1]_net_1\, Y => m6_0_a3_0);
    
    \HADDR_d[14]\ : SLE
      port map(D => M0GATEDHADDR(14), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(14));
    
    \burst_count_reg_RNIEB7I[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \count[0]_net_1\, B => 
        \burst_count_reg[0]_net_1\, Y => N_78_i);
    
    \HSIZE_d[1]\ : SLE
      port map(D => M0GATEDHSIZE(1), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_size(1));
    
    \count_RNO[2]\ : CFG2
      generic map(INIT => x"9")

      port map(A => N_85, B => \count[2]_net_1\, Y => N_93_i_0);
    
    \ahbcurr_state_ns_1_0_.N_23_i_1\ : CFG4
      generic map(INIT => x"4445")

      port map(A => m9_i_a3_1_0, B => \ahbcurr_state[1]_net_1\, C
         => M0GATEDHWRITE, D => defSlaveSMNextState_m, Y => 
        N_23_i_1);
    
    ahbsram_req_d1_RNIPK2R3 : CFG4
      generic map(INIT => x"FFCE")

      port map(A => N_80, B => un1_sramahb_ack_i_i_0, C => 
        ahbsram_req_d1_net_1, D => N_126, Y => counte);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \count_RNO[4]\ : CFG4
      generic map(INIT => x"D2F0")

      port map(A => \count[2]_net_1\, B => N_85, C => 
        \count[4]_net_1\, D => \count[3]_net_1\, Y => N_103_i_i_0);
    
    \ahbcurr_state_ns_1_0_.m6_0_o4\ : CFG3
      generic map(INIT => x"FD")

      port map(A => \ahbcurr_state[0]_net_1\, B => N_131, C => 
        \ahbcurr_state[1]_net_1\, Y => N_151);
    
    \ahbcurr_state[0]\ : SLE
      port map(D => \ahbcurr_state_ns[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ahbcurr_state[0]_net_1\);
    
    \ahbsram_req_d1\ : SLE
      port map(D => \CoreAHBLite_0_AHBmslave3_HREADY_i_1\, CLK
         => FAB_CCC_GL0, EN => VCC_net_1, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ahbsram_req_d1_net_1);
    
    \HADDR_d[9]\ : SLE
      port map(D => M0GATEDHADDR(9), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(9));
    
    \count_RNO[3]\ : CFG3
      generic map(INIT => x"D2")

      port map(A => \count[2]_net_1\, B => N_85, C => 
        \count[3]_net_1\, Y => N_94_i_0);
    
    \ahbcurr_state_ns_1_0_.m6_0_a2_4_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \count[2]_net_1\, B => \count[4]_net_1\, Y
         => m6_0_a2_4_0);
    
    \count_RNO[1]\ : CFG3
      generic map(INIT => x"12")

      port map(A => \count[0]_net_1\, B => un1_sramahb_ack_i_i_0, 
        C => \count[1]_net_1\, Y => N_5_i_0);
    
    \HADDR_d[8]\ : SLE
      port map(D => M0GATEDHADDR(8), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(8));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \count_RNIS3IO1[1]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => m6_0_a2_4_0, B => N_78_i, C => 
        \count[3]_net_1\, D => \count[1]_net_1\, Y => 
        un1_sramahb_ack_i_i_0);
    
    \count[2]\ : SLE
      port map(D => N_93_i_0, CLK => FAB_CCC_GL0, EN => counte, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \count[2]_net_1\);
    
    \ahbcurr_state[1]\ : SLE
      port map(D => N_23_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ahbcurr_state[1]_net_1\);
    
    \ahbcurr_state_RNI75PQ3_0[0]\ : CFG4
      generic map(INIT => x"030B")

      port map(A => sram_done, B => \ahbcurr_state[0]_net_1\, C
         => N_80, D => un1_sramahb_ack_i_i_0, Y => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0);
    
    \ahbcurr_state_ns_1_0_.m6_0\ : CFG4
      generic map(INIT => x"5755")

      port map(A => N_151, B => MASTERADDRINPROG_i_a2_0_a3_d_d(0), 
        C => MASTERADDRINPROG_i_a2_0_a3_0(0), D => m6_0_a3_2, Y
         => \ahbcurr_state_ns[0]\);
    
    \HADDR_d[12]\ : SLE
      port map(D => M0GATEDHADDR(12), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(12));
    
    \ahbcurr_state_ns_1_0_.m9_i_a3_1_0\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => sramcurr_state(0), B => sramcurr_state(1), C
         => m9_i_a3_0_0, D => \ahbcurr_state[0]_net_1\, Y => 
        m9_i_a3_1_0);
    
    ahbsram_req_d1_RNIIP8P : CFG3
      generic map(INIT => x"04")

      port map(A => sram_done, B => \ahbcurr_state[0]_net_1\, C
         => ahbsram_req_d1_net_1, Y => N_126);
    
    \HADDR_d[13]\ : SLE
      port map(D => M0GATEDHADDR(13), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(13));
    
    \HADDR_d[3]\ : SLE
      port map(D => M0GATEDHADDR(3), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(3));
    
    \ahbcurr_state_ns_1_0_.N_23_i\ : CFG4
      generic map(INIT => x"888A")

      port map(A => N_23_i_1, B => \ahbcurr_state[1]_net_1\, C
         => MASTERADDRINPROG_i_a2_0_a3_0(0), D => 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0), Y => N_23_i_0);
    
    \HADDR_d[10]\ : SLE
      port map(D => M0GATEDHADDR(10), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(10));
    
    \count[3]\ : SLE
      port map(D => N_94_i_0, CLK => FAB_CCC_GL0, EN => counte, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \count[3]_net_1\);
    
    \HSIZE_d[0]\ : SLE
      port map(D => M0GATEDHSIZE(0), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_size(0));
    
    count_n2_i_o4 : CFG2
      generic map(INIT => x"7")

      port map(A => \count[0]_net_1\, B => \count[1]_net_1\, Y
         => N_85);
    
    \burst_count_reg[0]\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => N_24_i_0, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \burst_count_reg[0]_net_1\);
    
    count_n0_i_a3 : CFG2
      generic map(INIT => x"1")

      port map(A => un1_sramahb_ack_i_i_0, B => \count[0]_net_1\, 
        Y => N_119);
    
    \ahbcurr_state_RNI75PQ3[0]\ : CFG4
      generic map(INIT => x"FCF4")

      port map(A => sram_done, B => \ahbcurr_state[0]_net_1\, C
         => N_80, D => un1_sramahb_ack_i_i_0, Y => 
        \CoreAHBLite_0_AHBmslave3_HREADY_i_1\);
    
    \ahbcurr_state_ns_1_0_.m6_0_a2_1_0\ : CFG4
      generic map(INIT => x"00A8")

      port map(A => sram_done, B => sramcurr_state(1), C => 
        sramcurr_state(0), D => N_78_i, Y => m6_0_a2_1);
    
    \ahbcurr_state_ns_1_0_.m6_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \count[3]_net_1\, B => \count[1]_net_1\, C
         => m6_0_a2_4_0, D => m6_0_a2_1, Y => N_131);
    
    \ahbcurr_state_ns_1_0_.m9_i_a3_0_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \ahbcurr_state[1]_net_1\, B => sram_done, Y
         => m9_i_a3_0_0);
    
    \HADDR_d[7]\ : SLE
      port map(D => M0GATEDHADDR(7), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(7));
    
    \HADDR_d[6]\ : SLE
      port map(D => M0GATEDHADDR(6), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(6));
    
    \burst_count_reg_RNO[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => MASTERADDRINPROG_i_a2_0_a3_d_d(0), B => 
        MASTERADDRINPROG_i_a2_0_a3_0(0), C => 
        \CoreAHBLite_0_AHBmslave3_HREADY_i_1\, D => 
        defSlaveSMNextState_m, Y => N_24_i_0);
    
    \HADDR_d[2]\ : SLE
      port map(D => M0GATEDHADDR(2), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(2));
    
    \HADDR_d[4]\ : SLE
      port map(D => M0GATEDHADDR(4), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(4));
    
    \HADDR_d[5]\ : SLE
      port map(D => M0GATEDHADDR(5), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(5));
    
    \HADDR_d[0]\ : SLE
      port map(D => M0GATEDHADDR(0), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(0));
    
    \count[4]\ : SLE
      port map(D => N_103_i_i_0, CLK => FAB_CCC_GL0, EN => counte, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \count[4]_net_1\);
    
    \HADDR_d[11]\ : SLE
      port map(D => M0GATEDHADDR(11), CLK => FAB_CCC_GL0, EN => 
        N_25_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_addr(11));
    
    \ahbcurr_state_RNIIV291[1]\ : CFG4
      generic map(INIT => x"CCDC")

      port map(A => sramcurr_state(1), B => 
        \ahbcurr_state[1]_net_1\, C => \ahbcurr_state[0]_net_1\, 
        D => sramcurr_state(0), Y => N_80);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM is

    port( M0GATEDHSIZE                            : in    std_logic_vector(1 downto 0);
          M0GATEDHADDR                            : in    std_logic_vector(15 downto 0);
          MASTERADDRINPROG_i_a2_0_a3_0            : in    std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_d_d          : in    std_logic_vector(0 to 0);
          CoreAHBLite_0_AHBmslave3_HRDATA         : out   std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave3_HWDATA         : in    std_logic_vector(31 downto 0);
          MSS_READY                               : in    std_logic;
          FAB_CCC_GL0                             : in    std_logic;
          N_25_i_0                                : in    std_logic;
          N_7_i_0                                 : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1     : out   std_logic;
          M0GATEDHWRITE                           : in    std_logic;
          defSlaveSMNextState_m                   : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3         : in    std_logic;
          defSlaveSMCurrentState                  : in    std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_2         : in    std_logic
        );

end CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM;

architecture DEF_ARCH of 
        CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf
    port( CoreAHBLite_0_AHBmslave3_HRDATA : out   std_logic_vector(31 downto 0);
          sramcurr_state                  : out   std_logic_vector(1 downto 0);
          ahbsram_size                    : in    std_logic_vector(1 downto 0) := (others => 'U');
          ahbcurr_state                   : in    std_logic_vector(1 downto 0) := (others => 'U');
          ahbsram_addr                    : in    std_logic_vector(15 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HWDATA : in    std_logic_vector(31 downto 0) := (others => 'U');
          MSS_READY                       : in    std_logic := 'U';
          FAB_CCC_GL0                     : in    std_logic := 'U';
          sram_done                       : out   std_logic;
          ahbsram_req_d1                  : in    std_logic := 'U';
          HWRITE_d                        : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf
    port( ahbsram_size                            : out   std_logic_vector(1 downto 0);
          M0GATEDHSIZE                            : in    std_logic_vector(1 downto 0) := (others => 'U');
          ahbsram_addr                            : out   std_logic_vector(15 downto 0);
          M0GATEDHADDR                            : in    std_logic_vector(15 downto 0) := (others => 'U');
          ahbcurr_state                           : out   std_logic_vector(1 downto 0);
          MASTERADDRINPROG_i_a2_0_a3_0            : in    std_logic_vector(0 to 0) := (others => 'U');
          MASTERADDRINPROG_i_a2_0_a3_d_d          : in    std_logic_vector(0 to 0) := (others => 'U');
          sramcurr_state                          : in    std_logic_vector(1 downto 0) := (others => 'U');
          MSS_READY                               : in    std_logic := 'U';
          FAB_CCC_GL0                             : in    std_logic := 'U';
          N_25_i_0                                : in    std_logic := 'U';
          HWRITE_d                                : out   std_logic;
          N_7_i_0                                 : in    std_logic := 'U';
          ahbsram_req_d1                          : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1     : out   std_logic;
          M0GATEDHWRITE                           : in    std_logic := 'U';
          defSlaveSMNextState_m                   : in    std_logic := 'U';
          sram_done                               : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3         : in    std_logic := 'U';
          defSlaveSMCurrentState                  : in    std_logic := 'U';
          un1_hready_m_xhdl342_1_i_0_o3_2         : in    std_logic := 'U'
        );
  end component;

    signal \ahbsram_size[0]\, \ahbsram_size[1]\, 
        \ahbsram_addr[0]\, \ahbsram_addr[1]\, \ahbsram_addr[2]\, 
        \ahbsram_addr[3]\, \ahbsram_addr[4]\, \ahbsram_addr[5]\, 
        \ahbsram_addr[6]\, \ahbsram_addr[7]\, \ahbsram_addr[8]\, 
        \ahbsram_addr[9]\, \ahbsram_addr[10]\, \ahbsram_addr[11]\, 
        \ahbsram_addr[12]\, \ahbsram_addr[13]\, 
        \ahbsram_addr[14]\, \ahbsram_addr[15]\, 
        \ahbcurr_state[0]\, \ahbcurr_state[1]\, 
        \sramcurr_state[0]\, \sramcurr_state[1]\, HWRITE_d, 
        ahbsram_req_d1, sram_done, GND_net_1, VCC_net_1
         : std_logic;

    for all : CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf
	Use entity work.
        CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf(DEF_ARCH);
    for all : CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf
	Use entity work.
        CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    U_SramCtrlIf : 
        CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf
      port map(CoreAHBLite_0_AHBmslave3_HRDATA(31) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(31), 
        CoreAHBLite_0_AHBmslave3_HRDATA(30) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(30), 
        CoreAHBLite_0_AHBmslave3_HRDATA(29) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(29), 
        CoreAHBLite_0_AHBmslave3_HRDATA(28) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(28), 
        CoreAHBLite_0_AHBmslave3_HRDATA(27) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(27), 
        CoreAHBLite_0_AHBmslave3_HRDATA(26) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(26), 
        CoreAHBLite_0_AHBmslave3_HRDATA(25) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(25), 
        CoreAHBLite_0_AHBmslave3_HRDATA(24) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(24), 
        CoreAHBLite_0_AHBmslave3_HRDATA(23) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(23), 
        CoreAHBLite_0_AHBmslave3_HRDATA(22) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(22), 
        CoreAHBLite_0_AHBmslave3_HRDATA(21) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(21), 
        CoreAHBLite_0_AHBmslave3_HRDATA(20) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(20), 
        CoreAHBLite_0_AHBmslave3_HRDATA(19) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(19), 
        CoreAHBLite_0_AHBmslave3_HRDATA(18) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(18), 
        CoreAHBLite_0_AHBmslave3_HRDATA(17) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(17), 
        CoreAHBLite_0_AHBmslave3_HRDATA(16) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(16), 
        CoreAHBLite_0_AHBmslave3_HRDATA(15) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(15), 
        CoreAHBLite_0_AHBmslave3_HRDATA(14) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(14), 
        CoreAHBLite_0_AHBmslave3_HRDATA(13) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(13), 
        CoreAHBLite_0_AHBmslave3_HRDATA(12) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(12), 
        CoreAHBLite_0_AHBmslave3_HRDATA(11) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(11), 
        CoreAHBLite_0_AHBmslave3_HRDATA(10) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(10), 
        CoreAHBLite_0_AHBmslave3_HRDATA(9) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(9), 
        CoreAHBLite_0_AHBmslave3_HRDATA(8) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(8), 
        CoreAHBLite_0_AHBmslave3_HRDATA(7) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(7), 
        CoreAHBLite_0_AHBmslave3_HRDATA(6) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(6), 
        CoreAHBLite_0_AHBmslave3_HRDATA(5) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(5), 
        CoreAHBLite_0_AHBmslave3_HRDATA(4) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(4), 
        CoreAHBLite_0_AHBmslave3_HRDATA(3) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(3), 
        CoreAHBLite_0_AHBmslave3_HRDATA(2) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(2), 
        CoreAHBLite_0_AHBmslave3_HRDATA(1) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(1), 
        CoreAHBLite_0_AHBmslave3_HRDATA(0) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(0), sramcurr_state(1) => 
        \sramcurr_state[1]\, sramcurr_state(0) => 
        \sramcurr_state[0]\, ahbsram_size(1) => \ahbsram_size[1]\, 
        ahbsram_size(0) => \ahbsram_size[0]\, ahbcurr_state(1)
         => \ahbcurr_state[1]\, ahbcurr_state(0) => 
        \ahbcurr_state[0]\, ahbsram_addr(15) => 
        \ahbsram_addr[15]\, ahbsram_addr(14) => 
        \ahbsram_addr[14]\, ahbsram_addr(13) => 
        \ahbsram_addr[13]\, ahbsram_addr(12) => 
        \ahbsram_addr[12]\, ahbsram_addr(11) => 
        \ahbsram_addr[11]\, ahbsram_addr(10) => 
        \ahbsram_addr[10]\, ahbsram_addr(9) => \ahbsram_addr[9]\, 
        ahbsram_addr(8) => \ahbsram_addr[8]\, ahbsram_addr(7) => 
        \ahbsram_addr[7]\, ahbsram_addr(6) => \ahbsram_addr[6]\, 
        ahbsram_addr(5) => \ahbsram_addr[5]\, ahbsram_addr(4) => 
        \ahbsram_addr[4]\, ahbsram_addr(3) => \ahbsram_addr[3]\, 
        ahbsram_addr(2) => \ahbsram_addr[2]\, ahbsram_addr(1) => 
        \ahbsram_addr[1]\, ahbsram_addr(0) => \ahbsram_addr[0]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(31) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(31), 
        CoreAHBLite_0_AHBmslave3_HWDATA(30) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(30), 
        CoreAHBLite_0_AHBmslave3_HWDATA(29) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(29), 
        CoreAHBLite_0_AHBmslave3_HWDATA(28) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(28), 
        CoreAHBLite_0_AHBmslave3_HWDATA(27) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(27), 
        CoreAHBLite_0_AHBmslave3_HWDATA(26) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(26), 
        CoreAHBLite_0_AHBmslave3_HWDATA(25) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(25), 
        CoreAHBLite_0_AHBmslave3_HWDATA(24) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(24), 
        CoreAHBLite_0_AHBmslave3_HWDATA(23) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(23), 
        CoreAHBLite_0_AHBmslave3_HWDATA(22) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(22), 
        CoreAHBLite_0_AHBmslave3_HWDATA(21) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(21), 
        CoreAHBLite_0_AHBmslave3_HWDATA(20) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(20), 
        CoreAHBLite_0_AHBmslave3_HWDATA(19) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(19), 
        CoreAHBLite_0_AHBmslave3_HWDATA(18) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(18), 
        CoreAHBLite_0_AHBmslave3_HWDATA(17) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(17), 
        CoreAHBLite_0_AHBmslave3_HWDATA(16) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(16), 
        CoreAHBLite_0_AHBmslave3_HWDATA(15) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(15), 
        CoreAHBLite_0_AHBmslave3_HWDATA(14) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(14), 
        CoreAHBLite_0_AHBmslave3_HWDATA(13) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(13), 
        CoreAHBLite_0_AHBmslave3_HWDATA(12) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(12), 
        CoreAHBLite_0_AHBmslave3_HWDATA(11) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(11), 
        CoreAHBLite_0_AHBmslave3_HWDATA(10) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(10), 
        CoreAHBLite_0_AHBmslave3_HWDATA(9) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(9), 
        CoreAHBLite_0_AHBmslave3_HWDATA(8) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(8), 
        CoreAHBLite_0_AHBmslave3_HWDATA(7) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(7), 
        CoreAHBLite_0_AHBmslave3_HWDATA(6) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(6), 
        CoreAHBLite_0_AHBmslave3_HWDATA(5) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(5), 
        CoreAHBLite_0_AHBmslave3_HWDATA(4) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(4), 
        CoreAHBLite_0_AHBmslave3_HWDATA(3) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(3), 
        CoreAHBLite_0_AHBmslave3_HWDATA(2) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(2), 
        CoreAHBLite_0_AHBmslave3_HWDATA(1) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(1), 
        CoreAHBLite_0_AHBmslave3_HWDATA(0) => 
        CoreAHBLite_0_AHBmslave3_HWDATA(0), MSS_READY => 
        MSS_READY, FAB_CCC_GL0 => FAB_CCC_GL0, sram_done => 
        sram_done, ahbsram_req_d1 => ahbsram_req_d1, HWRITE_d => 
        HWRITE_d);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    U_CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf : 
        CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf
      port map(ahbsram_size(1) => \ahbsram_size[1]\, 
        ahbsram_size(0) => \ahbsram_size[0]\, M0GATEDHSIZE(1) => 
        M0GATEDHSIZE(1), M0GATEDHSIZE(0) => M0GATEDHSIZE(0), 
        ahbsram_addr(15) => \ahbsram_addr[15]\, ahbsram_addr(14)
         => \ahbsram_addr[14]\, ahbsram_addr(13) => 
        \ahbsram_addr[13]\, ahbsram_addr(12) => 
        \ahbsram_addr[12]\, ahbsram_addr(11) => 
        \ahbsram_addr[11]\, ahbsram_addr(10) => 
        \ahbsram_addr[10]\, ahbsram_addr(9) => \ahbsram_addr[9]\, 
        ahbsram_addr(8) => \ahbsram_addr[8]\, ahbsram_addr(7) => 
        \ahbsram_addr[7]\, ahbsram_addr(6) => \ahbsram_addr[6]\, 
        ahbsram_addr(5) => \ahbsram_addr[5]\, ahbsram_addr(4) => 
        \ahbsram_addr[4]\, ahbsram_addr(3) => \ahbsram_addr[3]\, 
        ahbsram_addr(2) => \ahbsram_addr[2]\, ahbsram_addr(1) => 
        \ahbsram_addr[1]\, ahbsram_addr(0) => \ahbsram_addr[0]\, 
        M0GATEDHADDR(15) => M0GATEDHADDR(15), M0GATEDHADDR(14)
         => M0GATEDHADDR(14), M0GATEDHADDR(13) => 
        M0GATEDHADDR(13), M0GATEDHADDR(12) => M0GATEDHADDR(12), 
        M0GATEDHADDR(11) => M0GATEDHADDR(11), M0GATEDHADDR(10)
         => M0GATEDHADDR(10), M0GATEDHADDR(9) => M0GATEDHADDR(9), 
        M0GATEDHADDR(8) => M0GATEDHADDR(8), M0GATEDHADDR(7) => 
        M0GATEDHADDR(7), M0GATEDHADDR(6) => M0GATEDHADDR(6), 
        M0GATEDHADDR(5) => M0GATEDHADDR(5), M0GATEDHADDR(4) => 
        M0GATEDHADDR(4), M0GATEDHADDR(3) => M0GATEDHADDR(3), 
        M0GATEDHADDR(2) => M0GATEDHADDR(2), M0GATEDHADDR(1) => 
        M0GATEDHADDR(1), M0GATEDHADDR(0) => M0GATEDHADDR(0), 
        ahbcurr_state(1) => \ahbcurr_state[1]\, ahbcurr_state(0)
         => \ahbcurr_state[0]\, MASTERADDRINPROG_i_a2_0_a3_0(0)
         => MASTERADDRINPROG_i_a2_0_a3_0(0), 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0) => 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0), sramcurr_state(1) => 
        \sramcurr_state[1]\, sramcurr_state(0) => 
        \sramcurr_state[0]\, MSS_READY => MSS_READY, FAB_CCC_GL0
         => FAB_CCC_GL0, N_25_i_0 => N_25_i_0, HWRITE_d => 
        HWRITE_d, N_7_i_0 => N_7_i_0, ahbsram_req_d1 => 
        ahbsram_req_d1, CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, M0GATEDHWRITE => 
        M0GATEDHWRITE, defSlaveSMNextState_m => 
        defSlaveSMNextState_m, sram_done => sram_done, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, 
        un1_hready_m_xhdl342_1_i_0_o3_3 => 
        un1_hready_m_xhdl342_1_i_0_o3_3, defSlaveSMCurrentState
         => defSlaveSMCurrentState, 
        un1_hready_m_xhdl342_1_i_0_o3_2 => 
        un1_hready_m_xhdl342_1_i_0_o3_2);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb is

    port( DEVRST_N     : in    std_logic;
          SPI_0_SS0    : inout std_logic := 'Z';
          SPI_0_DO     : out   std_logic;
          SPI_0_DI     : in    std_logic;
          SPI_0_CLK    : inout std_logic := 'Z';
          MMUART_1_TXD : out   std_logic;
          MMUART_1_RXD : in    std_logic;
          GPIO_0_M2F_c : out   std_logic
        );

end CertificationSystem_sb;

architecture DEF_ARCH of CertificationSystem_sb is 

  component CertificationSystem_sb_FABOSC_0_OSC
    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );
  end component;

  component CoreResetP
    port( MSS_READY                                             : out   std_logic;
          FAB_CCC_GL0                                           : in    std_logic := 'U';
          POWER_ON_RESET_N                                      : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic := 'U'
        );
  end component;

  component CoreAHBLite
    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0) := (others => 'U');
          xhdl1250_i_m_1                                             : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : in    std_logic_vector(1 to 1) := (others => 'U');
          M0GATEDHSIZE                                               : out   std_logic_vector(1 downto 0);
          M0GATEDHADDR                                               : out   std_logic_vector(15 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HWDATA                            : out   std_logic_vector(31 downto 0);
          MASTERADDRINPROG_i_a2_0_a3_d_d                             : out   std_logic_vector(0 to 0);
          MASTERADDRINPROG_i_a2_0_a3_0                               : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28 : in    std_logic := 'U';
          MSS_READY                                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                                : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                        : in    std_logic := 'U';
          M0GATEDHWRITE                                              : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_2                            : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3                            : out   std_logic;
          defSlaveSMCurrentState                                     : out   std_logic;
          HREADY_M_iv_i_0                                            : out   std_logic;
          defSlaveSMNextState_m                                      : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                    : in    std_logic := 'U';
          N_7_i_0                                                    : out   std_logic;
          N_25_i_0                                                   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CertificationSystem_sb_MSS
    port( xhdl1250_i_m_1                                             : in    std_logic_vector(0 to 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HRDATA                            : in    std_logic_vector(31 downto 0) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE    : out   std_logic_vector(1 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS   : out   std_logic_vector(1 to 1);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA   : out   std_logic_vector(31 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP    : in    std_logic_vector(0 to 0) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31 : out   std_logic;
          SPI_0_SS0                                                  : inout   std_logic;
          SPI_0_DO                                                   : out   std_logic;
          SPI_0_DI                                                   : in    std_logic := 'U';
          SPI_0_CLK                                                  : inout   std_logic;
          MMUART_1_TXD                                               : out   std_logic;
          MMUART_1_RXD                                               : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N      : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F           : out   std_logic;
          GPIO_0_M2F_c                                               : out   std_logic;
          HREADY_M_iv_i_0                                            : in    std_logic := 'U';
          FAB_CCC_LOCK                                               : in    std_logic := 'U';
          FAB_CCC_GL0                                                : in    std_logic := 'U'
        );
  end component;

  component CertificationSystem_sb_CCC_0_FCCC
    port( FAB_CCC_GL0                                        : out   std_logic;
          FAB_CCC_LOCK                                       : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

  component CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM
    port( M0GATEDHSIZE                            : in    std_logic_vector(1 downto 0) := (others => 'U');
          M0GATEDHADDR                            : in    std_logic_vector(15 downto 0) := (others => 'U');
          MASTERADDRINPROG_i_a2_0_a3_0            : in    std_logic_vector(0 to 0) := (others => 'U');
          MASTERADDRINPROG_i_a2_0_a3_d_d          : in    std_logic_vector(0 to 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HRDATA         : out   std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave3_HWDATA         : in    std_logic_vector(31 downto 0) := (others => 'U');
          MSS_READY                               : in    std_logic := 'U';
          FAB_CCC_GL0                             : in    std_logic := 'U';
          N_25_i_0                                : in    std_logic := 'U';
          N_7_i_0                                 : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1     : out   std_logic;
          M0GATEDHWRITE                           : in    std_logic := 'U';
          defSlaveSMNextState_m                   : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 : out   std_logic;
          un1_hready_m_xhdl342_1_i_0_o3_3         : in    std_logic := 'U';
          defSlaveSMCurrentState                  : in    std_logic := 'U';
          un1_hready_m_xhdl342_1_i_0_o3_2         : in    std_logic := 'U'
        );
  end component;

    signal POWER_ON_RESET_N, FAB_CCC_GL0, FAB_CCC_LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        \xhdl1250_i_m_1[0]\, \CoreAHBLite_0_AHBmslave3_HRDATA[0]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[1]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[2]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[3]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[4]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[5]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[6]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[7]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[8]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[9]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[10]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[11]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[12]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[13]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[14]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[15]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[16]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[17]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[18]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[19]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[20]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[21]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[22]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[23]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[24]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[25]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[26]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[27]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[28]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[29]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[30]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[31]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[0]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[1]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[6]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[7]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[8]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[9]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[10]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[11]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[12]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[13]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[14]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[15]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[28]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[29]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[30]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[31]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[0]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[1]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        HREADY_M_iv_i_0, \M0GATEDHSIZE[0]\, \M0GATEDHSIZE[1]\, 
        \M0GATEDHADDR[0]\, \M0GATEDHADDR[1]\, \M0GATEDHADDR[2]\, 
        \M0GATEDHADDR[3]\, \M0GATEDHADDR[4]\, \M0GATEDHADDR[5]\, 
        \M0GATEDHADDR[6]\, \M0GATEDHADDR[7]\, \M0GATEDHADDR[8]\, 
        \M0GATEDHADDR[9]\, \M0GATEDHADDR[10]\, \M0GATEDHADDR[11]\, 
        \M0GATEDHADDR[12]\, \M0GATEDHADDR[13]\, 
        \M0GATEDHADDR[14]\, \M0GATEDHADDR[15]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[0]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[1]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[2]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[3]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[4]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[5]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[6]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[7]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[8]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[9]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[10]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[11]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[12]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[13]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[14]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[15]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[16]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[17]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[18]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[19]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[20]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[21]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[22]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[23]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[24]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[25]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[26]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[27]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[28]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[29]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[30]\, 
        \CoreAHBLite_0_AHBmslave3_HWDATA[31]\, 
        \MASTERADDRINPROG_i_a2_0_a3_d_d[0]\, 
        \MASTERADDRINPROG_i_a2_0_a3_0[0]\, MSS_READY, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, M0GATEDHWRITE, 
        un1_hready_m_xhdl342_1_i_0_o3_2, 
        un1_hready_m_xhdl342_1_i_0_o3_3, defSlaveSMCurrentState, 
        defSlaveSMNextState_m, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, N_7_i_0, 
        N_25_i_0, GND_net_1, VCC_net_1 : std_logic;

    for all : CertificationSystem_sb_FABOSC_0_OSC
	Use entity work.CertificationSystem_sb_FABOSC_0_OSC(DEF_ARCH);
    for all : CoreResetP
	Use entity work.CoreResetP(DEF_ARCH);
    for all : CoreAHBLite
	Use entity work.CoreAHBLite(DEF_ARCH);
    for all : CertificationSystem_sb_MSS
	Use entity work.CertificationSystem_sb_MSS(DEF_ARCH);
    for all : CertificationSystem_sb_CCC_0_FCCC
	Use entity work.CertificationSystem_sb_CCC_0_FCCC(DEF_ARCH);
    for all : CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM
	Use entity work.
        CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM(DEF_ARCH);
begin 


    FABOSC_0 : CertificationSystem_sb_FABOSC_0_OSC
      port map(FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
         => FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    CORERESETP_0 : CoreResetP
      port map(MSS_READY => MSS_READY, FAB_CCC_GL0 => FAB_CCC_GL0, 
        POWER_ON_RESET_N => POWER_ON_RESET_N, 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N);
    
    CoreAHBLite_0 : CoreAHBLite
      port map(
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[0]\, 
        xhdl1250_i_m_1(0) => \xhdl1250_i_m_1[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        M0GATEDHSIZE(1) => \M0GATEDHSIZE[1]\, M0GATEDHSIZE(0) => 
        \M0GATEDHSIZE[0]\, M0GATEDHADDR(15) => \M0GATEDHADDR[15]\, 
        M0GATEDHADDR(14) => \M0GATEDHADDR[14]\, M0GATEDHADDR(13)
         => \M0GATEDHADDR[13]\, M0GATEDHADDR(12) => 
        \M0GATEDHADDR[12]\, M0GATEDHADDR(11) => 
        \M0GATEDHADDR[11]\, M0GATEDHADDR(10) => 
        \M0GATEDHADDR[10]\, M0GATEDHADDR(9) => \M0GATEDHADDR[9]\, 
        M0GATEDHADDR(8) => \M0GATEDHADDR[8]\, M0GATEDHADDR(7) => 
        \M0GATEDHADDR[7]\, M0GATEDHADDR(6) => \M0GATEDHADDR[6]\, 
        M0GATEDHADDR(5) => \M0GATEDHADDR[5]\, M0GATEDHADDR(4) => 
        \M0GATEDHADDR[4]\, M0GATEDHADDR(3) => \M0GATEDHADDR[3]\, 
        M0GATEDHADDR(2) => \M0GATEDHADDR[2]\, M0GATEDHADDR(1) => 
        \M0GATEDHADDR[1]\, M0GATEDHADDR(0) => \M0GATEDHADDR[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(31) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[31]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(30) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[30]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(29) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[29]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(28) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[28]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(27) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[27]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(26) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[26]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(25) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[25]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(24) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[24]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(23) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[23]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(22) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[22]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(21) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[21]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(20) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[20]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(19) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[19]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(18) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[18]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(17) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[17]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(16) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[16]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(15) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[15]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(14) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[14]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(13) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[13]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(12) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[12]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(11) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[11]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(10) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[10]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(9) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[9]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(8) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[8]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(7) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[7]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(6) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[6]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(5) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[5]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(4) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[4]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(3) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[3]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(2) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[2]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(1) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[1]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(0) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[0]\, 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0) => 
        \MASTERADDRINPROG_i_a2_0_a3_d_d[0]\, 
        MASTERADDRINPROG_i_a2_0_a3_0(0) => 
        \MASTERADDRINPROG_i_a2_0_a3_0[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[12]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[14]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[6]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[7]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[8]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[9]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[10]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[11]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[31]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[30]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[29]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[28]\, 
        MSS_READY => MSS_READY, FAB_CCC_GL0 => FAB_CCC_GL0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, M0GATEDHWRITE => 
        M0GATEDHWRITE, un1_hready_m_xhdl342_1_i_0_o3_2 => 
        un1_hready_m_xhdl342_1_i_0_o3_2, 
        un1_hready_m_xhdl342_1_i_0_o3_3 => 
        un1_hready_m_xhdl342_1_i_0_o3_3, defSlaveSMCurrentState
         => defSlaveSMCurrentState, HREADY_M_iv_i_0 => 
        HREADY_M_iv_i_0, defSlaveSMNextState_m => 
        defSlaveSMNextState_m, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, N_7_i_0 => 
        N_7_i_0, N_25_i_0 => N_25_i_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    CertificationSystem_sb_MSS_0 : CertificationSystem_sb_MSS
      port map(xhdl1250_i_m_1(0) => \xhdl1250_i_m_1[0]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(31) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[31]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(30) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[30]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(29) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[29]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(28) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[28]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(27) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[27]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(26) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[26]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(25) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[25]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(24) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[24]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(23) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[23]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(22) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[22]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(21) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[21]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(20) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[20]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(19) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[19]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(18) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[18]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(17) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[17]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(16) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[16]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(15) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[15]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(14) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[14]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(13) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[13]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(12) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[12]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(11) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[11]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(10) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[10]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(9) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[9]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(8) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[8]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(7) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[7]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(6) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[6]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(5) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[5]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(4) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[4]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(3) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[3]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(2) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[2]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(1) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[1]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(0) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[6]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[7]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[8]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[9]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[10]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[11]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[12]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[14]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[28]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[29]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[30]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[31]\, 
        SPI_0_SS0 => SPI_0_SS0, SPI_0_DO => SPI_0_DO, SPI_0_DI
         => SPI_0_DI, SPI_0_CLK => SPI_0_CLK, MMUART_1_TXD => 
        MMUART_1_TXD, MMUART_1_RXD => MMUART_1_RXD, 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        GPIO_0_M2F_c => GPIO_0_M2F_c, HREADY_M_iv_i_0 => 
        HREADY_M_iv_i_0, FAB_CCC_LOCK => FAB_CCC_LOCK, 
        FAB_CCC_GL0 => FAB_CCC_GL0);
    
    CCC_0 : CertificationSystem_sb_CCC_0_FCCC
      port map(FAB_CCC_GL0 => FAB_CCC_GL0, FAB_CCC_LOCK => 
        FAB_CCC_LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => POWER_ON_RESET_N, DEVRST_N => 
        DEVRST_N);
    
    COREAHBLSRAM_0_0 : 
        CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM
      port map(M0GATEDHSIZE(1) => \M0GATEDHSIZE[1]\, 
        M0GATEDHSIZE(0) => \M0GATEDHSIZE[0]\, M0GATEDHADDR(15)
         => \M0GATEDHADDR[15]\, M0GATEDHADDR(14) => 
        \M0GATEDHADDR[14]\, M0GATEDHADDR(13) => 
        \M0GATEDHADDR[13]\, M0GATEDHADDR(12) => 
        \M0GATEDHADDR[12]\, M0GATEDHADDR(11) => 
        \M0GATEDHADDR[11]\, M0GATEDHADDR(10) => 
        \M0GATEDHADDR[10]\, M0GATEDHADDR(9) => \M0GATEDHADDR[9]\, 
        M0GATEDHADDR(8) => \M0GATEDHADDR[8]\, M0GATEDHADDR(7) => 
        \M0GATEDHADDR[7]\, M0GATEDHADDR(6) => \M0GATEDHADDR[6]\, 
        M0GATEDHADDR(5) => \M0GATEDHADDR[5]\, M0GATEDHADDR(4) => 
        \M0GATEDHADDR[4]\, M0GATEDHADDR(3) => \M0GATEDHADDR[3]\, 
        M0GATEDHADDR(2) => \M0GATEDHADDR[2]\, M0GATEDHADDR(1) => 
        \M0GATEDHADDR[1]\, M0GATEDHADDR(0) => \M0GATEDHADDR[0]\, 
        MASTERADDRINPROG_i_a2_0_a3_0(0) => 
        \MASTERADDRINPROG_i_a2_0_a3_0[0]\, 
        MASTERADDRINPROG_i_a2_0_a3_d_d(0) => 
        \MASTERADDRINPROG_i_a2_0_a3_d_d[0]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(31) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[31]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(30) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[30]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(29) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[29]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(28) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[28]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(27) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[27]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(26) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[26]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(25) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[25]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(24) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[24]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(23) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[23]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(22) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[22]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(21) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[21]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(20) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[20]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(19) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[19]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(18) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[18]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(17) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[17]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(16) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[16]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(15) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[15]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(14) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[14]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(13) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[13]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(12) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[12]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(11) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[11]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(10) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[10]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(9) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[9]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(8) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[8]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(7) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[7]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(6) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[6]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(5) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[5]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(4) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[4]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(3) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[3]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(2) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[2]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(1) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[1]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(0) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[0]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(31) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[31]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(30) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[30]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(29) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[29]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(28) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[28]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(27) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[27]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(26) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[26]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(25) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[25]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(24) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[24]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(23) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[23]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(22) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[22]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(21) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[21]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(20) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[20]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(19) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[19]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(18) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[18]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(17) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[17]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(16) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[16]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(15) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[15]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(14) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[14]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(13) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[13]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(12) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[12]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(11) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[11]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(10) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[10]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(9) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[9]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(8) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[8]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(7) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[7]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(6) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[6]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(5) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[5]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(4) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[4]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(3) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[3]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(2) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[2]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(1) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[1]\, 
        CoreAHBLite_0_AHBmslave3_HWDATA(0) => 
        \CoreAHBLite_0_AHBmslave3_HWDATA[0]\, MSS_READY => 
        MSS_READY, FAB_CCC_GL0 => FAB_CCC_GL0, N_25_i_0 => 
        N_25_i_0, N_7_i_0 => N_7_i_0, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, M0GATEDHWRITE => 
        M0GATEDHWRITE, defSlaveSMNextState_m => 
        defSlaveSMNextState_m, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, 
        un1_hready_m_xhdl342_1_i_0_o3_3 => 
        un1_hready_m_xhdl342_1_i_0_o3_3, defSlaveSMCurrentState
         => defSlaveSMCurrentState, 
        un1_hready_m_xhdl342_1_i_0_o3_2 => 
        un1_hready_m_xhdl342_1_i_0_o3_2);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem is

    port( DEVRST_N     : in    std_logic;
          MMUART_1_RXD : in    std_logic;
          SPI_0_DI     : in    std_logic;
          GPIO_0_M2F   : out   std_logic;
          MMUART_1_TXD : out   std_logic;
          SPI_0_DO     : out   std_logic;
          SPI_0_CLK    : inout std_logic := 'Z';
          SPI_0_SS0    : inout std_logic := 'Z'
        );

end CertificationSystem;

architecture DEF_ARCH of CertificationSystem is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CertificationSystem_sb
    port( DEVRST_N     : in    std_logic := 'U';
          SPI_0_SS0    : inout   std_logic;
          SPI_0_DO     : out   std_logic;
          SPI_0_DI     : in    std_logic := 'U';
          SPI_0_CLK    : inout   std_logic;
          MMUART_1_TXD : out   std_logic;
          MMUART_1_RXD : in    std_logic := 'U';
          GPIO_0_M2F_c : out   std_logic
        );
  end component;

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1, GPIO_0_M2F_c : std_logic;

    for all : CertificationSystem_sb
	Use entity work.CertificationSystem_sb(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    CertificationSystem_sb_0 : CertificationSystem_sb
      port map(DEVRST_N => DEVRST_N, SPI_0_SS0 => SPI_0_SS0, 
        SPI_0_DO => SPI_0_DO, SPI_0_DI => SPI_0_DI, SPI_0_CLK => 
        SPI_0_CLK, MMUART_1_TXD => MMUART_1_TXD, MMUART_1_RXD => 
        MMUART_1_RXD, GPIO_0_M2F_c => GPIO_0_M2F_c);
    
    GPIO_0_M2F_obuf : OUTBUF
      port map(D => GPIO_0_M2F_c, PAD => GPIO_0_M2F);
    

end DEF_ARCH; 
