-- Version: v11.7 SP1 11.7.1.14

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_controller is

    port( sha256_controller_0_read_addr_0      : out   std_logic_vector(3 downto 0);
          reg_17x32_0_last_word                : in    std_logic_vector(3 downto 0);
          di_o_0                               : in    std_logic_vector(1 to 1);
          state_1                              : out   std_logic;
          state_4                              : out   std_logic;
          state_3                              : out   std_logic;
          sha256_controller_0_di_o_5           : out   std_logic;
          sha256_controller_0_di_o_3           : out   std_logic;
          sha256_controller_0_di_o_0           : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F  : in    std_logic;
          SHA256_Module_0_waiting_data         : out   std_logic;
          bytes_sel                            : out   std_logic;
          N_484                                : out   std_logic;
          data_out_ready                       : in    std_logic;
          prev_sig                             : in    std_logic;
          prev_sig_0                           : in    std_logic;
          first_block                          : in    std_logic;
          SHA256_Module_0_di_req_o             : in    std_logic;
          SHA256_BLOCK_0_do_valid_o            : in    std_logic;
          N_1705                               : in    std_logic;
          N_1703                               : in    std_logic;
          N_1700                               : in    std_logic;
          SHA256_BLOCK_0_start_o               : out   std_logic
        );

end sha256_controller;

architecture DEF_ARCH of sha256_controller is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal un2_rst_n_i, \un2_rst_n\, \blocks_counter[0]_net_1\, 
        \blocks_counter_s[0]\, 
        \sha256_controller_0_read_addr_0[1]\, VCC_net_1, 
        N_694_i_0_i, \counter_4[1]\, GND_net_1, 
        \sha256_controller_0_read_addr_0[2]\, \counter_4[2]\, 
        \sha256_controller_0_read_addr_0[3]\, N_482_i_0, 
        \sha256_controller_0_read_addr_0[0]\, \counter_4[0]\, 
        \state_1\, N_100_i_0, \state[0]_net_1\, \state_ns[5]\, 
        \SHA256_Module_0_waiting_data\, \state_ns[0]\, \state_4\, 
        \state_ns_i_i_a2[1]_net_1\, \state_3\, \state_ns[2]\, 
        \state[2]_net_1\, N_98_i_0, \un1_state_2_0_a3_0_a2\, 
        \blocks_counter[1]_net_1\, \blocks_counter_s[1]\, 
        \blocks_counter[2]_net_1\, \blocks_counter_s[2]\, 
        \blocks_counter[3]_net_1\, \blocks_counter_s[3]\, 
        \blocks_counter[4]_net_1\, \blocks_counter_s[4]\, 
        \blocks_counter[5]_net_1\, \blocks_counter_s[5]\, 
        \blocks_counter[6]_net_1\, \blocks_counter_s[6]\, 
        \blocks_counter[7]_net_1\, \blocks_counter_s[7]\, 
        \blocks_counter[8]_net_1\, \blocks_counter_s[8]\, 
        \blocks_counter[9]_net_1\, \blocks_counter_s[9]\, 
        \blocks_counter[10]_net_1\, \blocks_counter_s[10]\, 
        \blocks_counter[11]_net_1\, \blocks_counter_s[11]\, 
        \blocks_counter[12]_net_1\, \blocks_counter_s[12]\, 
        \blocks_counter[13]_net_1\, \blocks_counter_s[13]\, 
        \blocks_counter[14]_net_1\, \blocks_counter_s[14]\, 
        \blocks_counter[15]_net_1\, \blocks_counter_s[15]\, 
        \blocks_counter[16]_net_1\, \blocks_counter_s[16]\, 
        \blocks_counter[17]_net_1\, \blocks_counter_s[17]\, 
        \blocks_counter[18]_net_1\, \blocks_counter_s[18]\, 
        \blocks_counter[19]_net_1\, \blocks_counter_s[19]\, 
        \blocks_counter[20]_net_1\, \blocks_counter_s[20]\, 
        \blocks_counter[21]_net_1\, \blocks_counter_s[21]\, 
        \blocks_counter[22]_net_1\, \blocks_counter_s[22]\, 
        \blocks_counter[23]_net_1\, \blocks_counter_s[23]\, 
        \blocks_counter[24]_net_1\, \blocks_counter_s[24]\, 
        \blocks_counter[25]_net_1\, \blocks_counter_s[25]\, 
        \blocks_counter[26]_net_1\, \blocks_counter_s[26]\, 
        \blocks_counter[27]_net_1\, \blocks_counter_s[27]\, 
        \blocks_counter[28]_net_1\, \blocks_counter_s[28]\, 
        \blocks_counter[29]_net_1\, \blocks_counter_s[29]\, 
        \blocks_counter[30]_net_1\, \blocks_counter_s[30]\, 
        \blocks_counter[31]_net_1\, \blocks_counter_s[31]_net_1\, 
        blocks_counter_s_970_FCO, \blocks_counter_cry[1]_net_1\, 
        \blocks_counter_cry[2]_net_1\, 
        \blocks_counter_cry[3]_net_1\, 
        \blocks_counter_cry[4]_net_1\, 
        \blocks_counter_cry[5]_net_1\, 
        \blocks_counter_cry[6]_net_1\, 
        \blocks_counter_cry[7]_net_1\, 
        \blocks_counter_cry[8]_net_1\, 
        \blocks_counter_cry[9]_net_1\, 
        \blocks_counter_cry[10]_net_1\, 
        \blocks_counter_cry[11]_net_1\, 
        \blocks_counter_cry[12]_net_1\, 
        \blocks_counter_cry[13]_net_1\, 
        \blocks_counter_cry[14]_net_1\, 
        \blocks_counter_cry[15]_net_1\, 
        \blocks_counter_cry[16]_net_1\, 
        \blocks_counter_cry[17]_net_1\, 
        \blocks_counter_cry[18]_net_1\, 
        \blocks_counter_cry[19]_net_1\, 
        \blocks_counter_cry[20]_net_1\, 
        \blocks_counter_cry[21]_net_1\, 
        \blocks_counter_cry[22]_net_1\, 
        \blocks_counter_cry[23]_net_1\, 
        \blocks_counter_cry[24]_net_1\, 
        \blocks_counter_cry[25]_net_1\, 
        \blocks_counter_cry[26]_net_1\, 
        \blocks_counter_cry[27]_net_1\, 
        \blocks_counter_cry[28]_net_1\, 
        \blocks_counter_cry[29]_net_1\, 
        \blocks_counter_cry[30]_net_1\, N_494, N_491, N_760, 
        \N_484\, \start_o_0_sqmuxa_0_a2_23\, 
        \start_o_0_sqmuxa_0_a2_22\, \start_o_0_sqmuxa_0_a2_21\, 
        \start_o_0_sqmuxa_0_a2_20\, \start_o_0_sqmuxa_0_a2_19\, 
        \start_o_0_sqmuxa_0_a2_18\, \start_o_0_sqmuxa_0_a2_17\, 
        \start_o_0_sqmuxa_0_a2_16\, \state_ns_0_o3_2[2]_net_1\, 
        \state_ns_i_0_o2_0[4]_net_1\, N_493, N_717, N_698, N_497, 
        N_709, \start_o_0_sqmuxa_0_a2_29\, 
        \start_o_0_sqmuxa_0_a2_28\, N_701 : std_logic;

begin 

    sha256_controller_0_read_addr_0(3) <= 
        \sha256_controller_0_read_addr_0[3]\;
    sha256_controller_0_read_addr_0(2) <= 
        \sha256_controller_0_read_addr_0[2]\;
    sha256_controller_0_read_addr_0(1) <= 
        \sha256_controller_0_read_addr_0[1]\;
    sha256_controller_0_read_addr_0(0) <= 
        \sha256_controller_0_read_addr_0[0]\;
    state_1 <= \state_1\;
    state_4 <= \state_4\;
    state_3 <= \state_3\;
    SHA256_Module_0_waiting_data <= 
        \SHA256_Module_0_waiting_data\;
    N_484 <= \N_484\;

    \state_ns_0_o3_2[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => reg_17x32_0_last_word(3), B => 
        reg_17x32_0_last_word(2), C => reg_17x32_0_last_word(1), 
        D => reg_17x32_0_last_word(0), Y => 
        \state_ns_0_o3_2[2]_net_1\);
    
    start_o_0_sqmuxa_0_a2 : CFG4
      generic map(INIT => x"8000")

      port map(A => \start_o_0_sqmuxa_0_a2_21\, B => 
        \start_o_0_sqmuxa_0_a2_22\, C => 
        \start_o_0_sqmuxa_0_a2_28\, D => 
        \start_o_0_sqmuxa_0_a2_29\, Y => SHA256_BLOCK_0_start_o);
    
    \bytes_sel\ : SLE
      port map(D => \state_1\, CLK => \un1_state_2_0_a3_0_a2\, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        bytes_sel);
    
    \blocks_counter_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[2]_net_1\, S => \blocks_counter_s[3]\, 
        Y => OPEN, FCO => \blocks_counter_cry[3]_net_1\);
    
    \blocks_counter_cry[26]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[26]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[25]_net_1\, S => 
        \blocks_counter_s[26]\, Y => OPEN, FCO => 
        \blocks_counter_cry[26]_net_1\);
    
    \blocks_counter[31]\ : SLE
      port map(D => \blocks_counter_s[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[31]_net_1\);
    
    \blocks_counter_s[31]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[31]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[30]_net_1\, S => 
        \blocks_counter_s[31]_net_1\, Y => OPEN, FCO => OPEN);
    
    \blocks_counter_cry[22]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[22]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[21]_net_1\, S => 
        \blocks_counter_s[22]\, Y => OPEN, FCO => 
        \blocks_counter_cry[22]_net_1\);
    
    \counter_4_0_o3_0[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \sha256_controller_0_read_addr_0[3]\, B => 
        \sha256_controller_0_read_addr_0[2]\, C => 
        \sha256_controller_0_read_addr_0[1]\, D => 
        \sha256_controller_0_read_addr_0[0]\, Y => N_493);
    
    \counter_4_0_a2_1[0]\ : CFG3
      generic map(INIT => x"20")

      port map(A => SHA256_Module_0_di_req_o, B => N_493, C => 
        \state[2]_net_1\, Y => N_709);
    
    \blocks_counter_cry[25]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[25]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[24]_net_1\, S => 
        \blocks_counter_s[25]\, Y => OPEN, FCO => 
        \blocks_counter_cry[25]_net_1\);
    
    blocks_counter_s_970 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => blocks_counter_s_970_FCO);
    
    \blocks_counter_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        blocks_counter_s_970_FCO, S => \blocks_counter_s[1]\, Y
         => OPEN, FCO => \blocks_counter_cry[1]_net_1\);
    
    \blocks_counter_cry[16]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[16]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[15]_net_1\, S => 
        \blocks_counter_s[16]\, Y => OPEN, FCO => 
        \blocks_counter_cry[16]_net_1\);
    
    \counter[2]\ : SLE
      port map(D => \counter_4[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => N_694_i_0_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sha256_controller_0_read_addr_0[2]\);
    
    \blocks_counter_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[11]_net_1\, S => 
        \blocks_counter_s[12]\, Y => OPEN, FCO => 
        \blocks_counter_cry[12]_net_1\);
    
    \blocks_counter[20]\ : SLE
      port map(D => \blocks_counter_s[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[20]_net_1\);
    
    \blocks_counter[13]\ : SLE
      port map(D => \blocks_counter_s[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[13]_net_1\);
    
    \state[5]\ : SLE
      port map(D => \state_ns[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_0_GPIO_9_M2F, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SHA256_Module_0_waiting_data\);
    
    start_o_0_sqmuxa_0_a2_19 : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[8]_net_1\, B => 
        \blocks_counter[7]_net_1\, C => \blocks_counter[2]_net_1\, 
        D => \blocks_counter[1]_net_1\, Y => 
        \start_o_0_sqmuxa_0_a2_19\);
    
    \blocks_counter_cry[15]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[14]_net_1\, S => 
        \blocks_counter_s[15]\, Y => OPEN, FCO => 
        \blocks_counter_cry[15]_net_1\);
    
    \blocks_counter[26]\ : SLE
      port map(D => \blocks_counter_s[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[26]_net_1\);
    
    \blocks_counter[15]\ : SLE
      port map(D => \blocks_counter_s[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[15]_net_1\);
    
    start_o_0_sqmuxa_0_a2_18 : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[14]_net_1\, B => 
        \blocks_counter[13]_net_1\, C => 
        \blocks_counter[4]_net_1\, D => \blocks_counter[3]_net_1\, 
        Y => \start_o_0_sqmuxa_0_a2_18\);
    
    \blocks_counter[30]\ : SLE
      port map(D => \blocks_counter_s[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[30]_net_1\);
    
    \state[4]\ : SLE
      port map(D => \state_ns_i_i_a2[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_0_GPIO_9_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \state_4\);
    
    \blocks_counter[0]\ : SLE
      port map(D => \blocks_counter_s[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[0]_net_1\);
    
    \blocks_counter_cry[23]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[23]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[22]_net_1\, S => 
        \blocks_counter_s[23]\, Y => OPEN, FCO => 
        \blocks_counter_cry[23]_net_1\);
    
    \state[2]\ : SLE
      port map(D => N_98_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_0_GPIO_9_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \state[2]_net_1\);
    
    start_o_0_sqmuxa_0_a2_20 : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[31]_net_1\, B => 
        \blocks_counter[30]_net_1\, C => 
        \blocks_counter[6]_net_1\, D => \blocks_counter[5]_net_1\, 
        Y => \start_o_0_sqmuxa_0_a2_20\);
    
    \state_ns_i_0_x3_2[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \sha256_controller_0_read_addr_0[0]\, B => 
        reg_17x32_0_last_word(0), Y => N_760);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \state_RNIJFAP[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => CertificationSystem_sb_0_GPIO_9_M2F, B => 
        \SHA256_Module_0_waiting_data\, Y => N_694_i_0_i);
    
    \blocks_counter[11]\ : SLE
      port map(D => \blocks_counter_s[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[11]_net_1\);
    
    \state[3]\ : SLE
      port map(D => \state_ns[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_0_GPIO_9_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \state_3\);
    
    \blocks_counter_cry[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[12]_net_1\, S => 
        \blocks_counter_s[13]\, Y => OPEN, FCO => 
        \blocks_counter_cry[13]_net_1\);
    
    \di_o[16]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1703, B => di_o_0(1), Y => 
        sha256_controller_0_di_o_3);
    
    \blocks_counter_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[1]_net_1\, S => \blocks_counter_s[2]\, 
        Y => OPEN, FCO => \blocks_counter_cry[2]_net_1\);
    
    \blocks_counter_cry[27]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[27]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[26]_net_1\, S => 
        \blocks_counter_s[27]\, Y => OPEN, FCO => 
        \blocks_counter_cry[27]_net_1\);
    
    \blocks_counter[24]\ : SLE
      port map(D => \blocks_counter_s[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[24]_net_1\);
    
    \blocks_counter_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[5]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[4]_net_1\, S => \blocks_counter_s[5]\, 
        Y => OPEN, FCO => \blocks_counter_cry[5]_net_1\);
    
    \state_ns_i_0_o2_0[4]\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => reg_17x32_0_last_word(3), B => 
        reg_17x32_0_last_word(1), C => 
        \sha256_controller_0_read_addr_0[3]\, D => 
        \sha256_controller_0_read_addr_0[1]\, Y => 
        \state_ns_i_0_o2_0[4]_net_1\);
    
    \blocks_counter_cry[28]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[28]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[27]_net_1\, S => 
        \blocks_counter_s[28]\, Y => OPEN, FCO => 
        \blocks_counter_cry[28]_net_1\);
    
    \blocks_counter[22]\ : SLE
      port map(D => \blocks_counter_s[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[22]_net_1\);
    
    \blocks_counter_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[8]_net_1\, S => \blocks_counter_s[9]\, 
        Y => OPEN, FCO => \blocks_counter_cry[9]_net_1\);
    
    un2_rst_n_RNIE1K2 : CLKINT
      port map(A => \un2_rst_n\, Y => un2_rst_n_i);
    
    \blocks_counter_cry[17]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[17]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[16]_net_1\, S => 
        \blocks_counter_s[17]\, Y => OPEN, FCO => 
        \blocks_counter_cry[17]_net_1\);
    
    \blocks_counter[5]\ : SLE
      port map(D => \blocks_counter_s[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[5]_net_1\);
    
    \blocks_counter[10]\ : SLE
      port map(D => \blocks_counter_s[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[10]_net_1\);
    
    \blocks_counter[16]\ : SLE
      port map(D => \blocks_counter_s[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[16]_net_1\);
    
    \state_ns_i_i_a2[1]\ : CFG3
      generic map(INIT => x"20")

      port map(A => data_out_ready, B => prev_sig, C => 
        \SHA256_Module_0_waiting_data\, Y => 
        \state_ns_i_i_a2[1]_net_1\);
    
    \counter_4_0[1]\ : CFG4
      generic map(INIT => x"66A2")

      port map(A => \sha256_controller_0_read_addr_0[1]\, B => 
        \sha256_controller_0_read_addr_0[0]\, C => N_491, D => 
        \N_484\, Y => \counter_4[1]\);
    
    \blocks_counter_cry[18]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[18]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[17]_net_1\, S => 
        \blocks_counter_s[18]\, Y => OPEN, FCO => 
        \blocks_counter_cry[18]_net_1\);
    
    di_wr_o_0_o3_i_o3 : CFG2
      generic map(INIT => x"E")

      port map(A => \state_1\, B => \state_3\, Y => \N_484\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \counter_4_0_o3[1]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \sha256_controller_0_read_addr_0[2]\, B => 
        \sha256_controller_0_read_addr_0[3]\, Y => N_491);
    
    \blocks_counter[1]\ : SLE
      port map(D => \blocks_counter_s[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[1]_net_1\);
    
    \blocks_counter[8]\ : SLE
      port map(D => \blocks_counter_s[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[8]_net_1\);
    
    \state[0]\ : SLE
      port map(D => \state_ns[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_0_GPIO_9_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \state[0]_net_1\);
    
    \blocks_counter[2]\ : SLE
      port map(D => \blocks_counter_s[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[2]_net_1\);
    
    \blocks_counter[27]\ : SLE
      port map(D => \blocks_counter_s[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[27]_net_1\);
    
    \blocks_counter[3]\ : SLE
      port map(D => \blocks_counter_s[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[3]_net_1\);
    
    \counter_RNO[3]\ : CFG4
      generic map(INIT => x"A6A2")

      port map(A => \sha256_controller_0_read_addr_0[3]\, B => 
        \sha256_controller_0_read_addr_0[2]\, C => N_494, D => 
        \N_484\, Y => N_482_i_0);
    
    \counter_4_0[0]\ : CFG4
      generic map(INIT => x"CFDC")

      port map(A => N_717, B => N_709, C => 
        \sha256_controller_0_read_addr_0[0]\, D => \N_484\, Y => 
        \counter_4[0]\);
    
    \blocks_counter_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[7]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[6]_net_1\, S => \blocks_counter_s[7]\, 
        Y => OPEN, FCO => \blocks_counter_cry[7]_net_1\);
    
    \blocks_counter_cry[30]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[30]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[29]_net_1\, S => 
        \blocks_counter_s[30]\, Y => OPEN, FCO => 
        \blocks_counter_cry[30]_net_1\);
    
    \blocks_counter[14]\ : SLE
      port map(D => \blocks_counter_s[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[14]_net_1\);
    
    \counter[1]\ : SLE
      port map(D => \counter_4[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => N_694_i_0_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sha256_controller_0_read_addr_0[1]\);
    
    start_o_0_sqmuxa_0_a2_17 : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[16]_net_1\, B => 
        \blocks_counter[15]_net_1\, C => 
        \blocks_counter[10]_net_1\, D => 
        \blocks_counter[9]_net_1\, Y => 
        \start_o_0_sqmuxa_0_a2_17\);
    
    \blocks_counter[12]\ : SLE
      port map(D => \blocks_counter_s[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[12]_net_1\);
    
    \counter[3]\ : SLE
      port map(D => N_482_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => N_694_i_0_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sha256_controller_0_read_addr_0[3]\);
    
    \blocks_counter_cry[21]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[21]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[20]_net_1\, S => 
        \blocks_counter_s[21]\, Y => OPEN, FCO => 
        \blocks_counter_cry[21]_net_1\);
    
    \state_ns_i_0_o2[4]\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \sha256_controller_0_read_addr_0[2]\, B => 
        reg_17x32_0_last_word(2), C => N_760, D => 
        \state_ns_i_0_o2_0[4]_net_1\, Y => N_497);
    
    \state_ns_0_a2[2]\ : CFG4
      generic map(INIT => x"A080")

      port map(A => SHA256_Module_0_di_req_o, B => N_493, C => 
        \state[2]_net_1\, D => \state_ns_0_o3_2[2]_net_1\, Y => 
        N_701);
    
    \counter_4_i_a2_0[3]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_494, B => N_491, Y => N_717);
    
    \di_o[18]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1705, B => di_o_0(1), Y => 
        sha256_controller_0_di_o_5);
    
    \blocks_counter_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \blocks_counter[0]_net_1\, Y => 
        \blocks_counter_s[0]\);
    
    start_o_0_sqmuxa_0_a2_22 : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[25]_net_1\, B => 
        \blocks_counter[22]_net_1\, C => 
        \blocks_counter[21]_net_1\, D => 
        \blocks_counter[0]_net_1\, Y => 
        \start_o_0_sqmuxa_0_a2_22\);
    
    \counter_4_0_o3[2]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \sha256_controller_0_read_addr_0[0]\, B => 
        \sha256_controller_0_read_addr_0[1]\, Y => N_494);
    
    \blocks_counter_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[4]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[3]_net_1\, S => \blocks_counter_s[4]\, 
        Y => OPEN, FCO => \blocks_counter_cry[4]_net_1\);
    
    \blocks_counter_cry[29]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[29]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[28]_net_1\, S => 
        \blocks_counter_s[29]\, Y => OPEN, FCO => 
        \blocks_counter_cry[29]_net_1\);
    
    \blocks_counter[28]\ : SLE
      port map(D => \blocks_counter_s[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[28]_net_1\);
    
    \state_ns_0_a2[0]\ : CFG3
      generic map(INIT => x"D0")

      port map(A => data_out_ready, B => prev_sig, C => 
        \SHA256_Module_0_waiting_data\, Y => N_698);
    
    \blocks_counter_cry[20]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[20]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[19]_net_1\, S => 
        \blocks_counter_s[20]\, Y => OPEN, FCO => 
        \blocks_counter_cry[20]_net_1\);
    
    \blocks_counter[29]\ : SLE
      port map(D => \blocks_counter_s[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[29]_net_1\);
    
    \state[1]\ : SLE
      port map(D => N_100_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_0_GPIO_9_M2F, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \state_1\);
    
    \blocks_counter_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[6]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[5]_net_1\, S => \blocks_counter_s[6]\, 
        Y => OPEN, FCO => \blocks_counter_cry[6]_net_1\);
    
    \blocks_counter[6]\ : SLE
      port map(D => \blocks_counter_s[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[6]_net_1\);
    
    un1_state_2_0_a3_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \state[0]_net_1\, B => \state[2]_net_1\, Y
         => \un1_state_2_0_a3_0_a2\);
    
    \blocks_counter_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[10]_net_1\, S => 
        \blocks_counter_s[11]\, Y => OPEN, FCO => 
        \blocks_counter_cry[11]_net_1\);
    
    \state_ns_0[2]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => \state_3\, B => SHA256_Module_0_di_req_o, C
         => N_497, D => N_701, Y => \state_ns[2]\);
    
    \blocks_counter_cry[19]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[19]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[18]_net_1\, S => 
        \blocks_counter_s[19]\, Y => OPEN, FCO => 
        \blocks_counter_cry[19]_net_1\);
    
    \blocks_counter[17]\ : SLE
      port map(D => \blocks_counter_s[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[17]_net_1\);
    
    \state_RNO[2]\ : CFG4
      generic map(INIT => x"F0FE")

      port map(A => \state_3\, B => \state[2]_net_1\, C => 
        \state_4\, D => SHA256_Module_0_di_req_o, Y => N_98_i_0);
    
    \blocks_counter_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[9]_net_1\, S => 
        \blocks_counter_s[10]\, Y => OPEN, FCO => 
        \blocks_counter_cry[10]_net_1\);
    
    \blocks_counter_cry[24]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[24]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[23]_net_1\, S => 
        \blocks_counter_s[24]\, Y => OPEN, FCO => 
        \blocks_counter_cry[24]_net_1\);
    
    \blocks_counter[7]\ : SLE
      port map(D => \blocks_counter_s[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[7]_net_1\);
    
    \state_ns_0[5]\ : CFG4
      generic map(INIT => x"F0F2")

      port map(A => \state[0]_net_1\, B => 
        SHA256_BLOCK_0_do_valid_o, C => \state_1\, D => 
        SHA256_Module_0_di_req_o, Y => \state_ns[5]\);
    
    start_o_0_sqmuxa_0_a2_21 : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[29]_net_1\, B => 
        \blocks_counter[28]_net_1\, C => 
        \blocks_counter[27]_net_1\, D => 
        \blocks_counter[26]_net_1\, Y => 
        \start_o_0_sqmuxa_0_a2_21\);
    
    \blocks_counter_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[7]_net_1\, S => \blocks_counter_s[8]\, 
        Y => OPEN, FCO => \blocks_counter_cry[8]_net_1\);
    
    \di_o[13]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1700, B => di_o_0(1), Y => 
        sha256_controller_0_di_o_0);
    
    \blocks_counter_cry[14]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \blocks_counter[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \blocks_counter_cry[13]_net_1\, S => 
        \blocks_counter_s[14]\, Y => OPEN, FCO => 
        \blocks_counter_cry[14]_net_1\);
    
    \blocks_counter[23]\ : SLE
      port map(D => \blocks_counter_s[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[23]_net_1\);
    
    \blocks_counter[25]\ : SLE
      port map(D => \blocks_counter_s[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[25]_net_1\);
    
    \counter_4_0[2]\ : CFG4
      generic map(INIT => x"C3C4")

      port map(A => \sha256_controller_0_read_addr_0[3]\, B => 
        \sha256_controller_0_read_addr_0[2]\, C => N_494, D => 
        \N_484\, Y => \counter_4[2]\);
    
    \blocks_counter[4]\ : SLE
      port map(D => \blocks_counter_s[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[4]_net_1\);
    
    start_o_0_sqmuxa_0_a2_29 : CFG4
      generic map(INIT => x"8000")

      port map(A => \start_o_0_sqmuxa_0_a2_20\, B => 
        \start_o_0_sqmuxa_0_a2_19\, C => 
        \start_o_0_sqmuxa_0_a2_18\, D => 
        \start_o_0_sqmuxa_0_a2_17\, Y => 
        \start_o_0_sqmuxa_0_a2_29\);
    
    \blocks_counter[18]\ : SLE
      port map(D => \blocks_counter_s[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[18]_net_1\);
    
    start_o_0_sqmuxa_0_a2_23 : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[24]_net_1\, B => 
        \blocks_counter[23]_net_1\, C => 
        \blocks_counter[18]_net_1\, D => 
        \blocks_counter[17]_net_1\, Y => 
        \start_o_0_sqmuxa_0_a2_23\);
    
    un2_rst_n : CFG3
      generic map(INIT => x"B0")

      port map(A => prev_sig_0, B => first_block, C => 
        CertificationSystem_sb_0_GPIO_9_M2F, Y => \un2_rst_n\);
    
    start_o_0_sqmuxa_0_a2_28 : CFG3
      generic map(INIT => x"80")

      port map(A => \start_o_0_sqmuxa_0_a2_16\, B => \state_4\, C
         => \start_o_0_sqmuxa_0_a2_23\, Y => 
        \start_o_0_sqmuxa_0_a2_28\);
    
    \blocks_counter[19]\ : SLE
      port map(D => \blocks_counter_s[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[19]_net_1\);
    
    \state_RNO[1]\ : CFG4
      generic map(INIT => x"0C08")

      port map(A => \state_3\, B => SHA256_Module_0_di_req_o, C
         => N_497, D => N_709, Y => N_100_i_0);
    
    \counter[0]\ : SLE
      port map(D => \counter_4[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => N_694_i_0_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sha256_controller_0_read_addr_0[0]\);
    
    \blocks_counter[9]\ : SLE
      port map(D => \blocks_counter_s[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[9]_net_1\);
    
    \blocks_counter[21]\ : SLE
      port map(D => \blocks_counter_s[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \state_4\, 
        ALn => un2_rst_n_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \blocks_counter[21]_net_1\);
    
    \state_ns_0[0]\ : CFG4
      generic map(INIT => x"FCEC")

      port map(A => SHA256_Module_0_di_req_o, B => N_698, C => 
        \state[0]_net_1\, D => SHA256_BLOCK_0_do_valid_o, Y => 
        \state_ns[0]\);
    
    start_o_0_sqmuxa_0_a2_16 : CFG4
      generic map(INIT => x"0001")

      port map(A => \blocks_counter[20]_net_1\, B => 
        \blocks_counter[19]_net_1\, C => 
        \blocks_counter[12]_net_1\, D => 
        \blocks_counter[11]_net_1\, Y => 
        \start_o_0_sqmuxa_0_a2_16\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_control is

    port( hash_control_st_reg_i                     : out   std_logic_vector(6 to 6);
          msg_bitlen                                : out   std_logic_vector(63 downto 3);
          Kt_addr                                   : out   std_logic_vector(5 downto 0);
          Kt_addr_fast                              : out   std_logic_vector(4 downto 0);
          state                                     : in    std_logic_vector(1 to 1);
          hash_control_st_reg_ns_i_0_a2_0           : out   std_logic_vector(4 to 4);
          reg_17x32_0_valid_bytes_0                 : in    std_logic_vector(1 downto 0);
          hash_control_st_reg_ns_i_0_a2_2           : in    std_logic_vector(4 to 4);
          hash_control_st_reg_2                     : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0      : in    std_logic;
          one_insert                                : out   std_logic;
          sha_last_blk_reg                          : out   std_logic;
          SHA256_Module_0_di_req_o                  : out   std_logic;
          SHA256_BLOCK_0_do_valid_o                 : out   std_logic;
          Kt_addr_1_rep1                            : out   std_logic;
          Kt_addr_1_rep2                            : out   std_logic;
          Kt_addr_2_rep1                            : out   std_logic;
          Kt_addr_2_rep2                            : out   std_logic;
          Kt_addr_0_rep1                            : out   std_logic;
          Kt_addr_0_rep2                            : out   std_logic;
          Kt_addr_4_rep1                            : out   std_logic;
          Kt_addr_4_rep2                            : out   std_logic;
          Kt_addr_3_rep1                            : out   std_logic;
          Kt_addr_3_rep2                            : out   std_logic;
          N_112                                     : out   std_logic;
          SHA256_Module_0_waiting_data              : in    std_logic;
          N_223                                     : out   std_logic;
          N_361                                     : out   std_logic;
          N_102                                     : out   std_logic;
          SHA256_Module_0_data_available_lastbank_8 : in    std_logic;
          N_168_i_0                                 : out   std_logic;
          pad_one_reg_0_0_a2_0                      : out   std_logic;
          oregs_ce_i_a2_0_a2                        : out   std_logic;
          sha_last_blk_next_0_o2_2_out_0            : out   std_logic;
          N_484                                     : in    std_logic;
          bytes_sel                                 : in    std_logic;
          sha_last_blk_next_0_a4_0                  : in    std_logic;
          N_388                                     : in    std_logic;
          N_111                                     : out   std_logic;
          core_ce_o_iv_i_0                          : out   std_logic;
          N_244_i_0                                 : out   std_logic;
          SHA256_Module_0_error_o                   : out   std_logic;
          ld_i_i_3                                  : out   std_logic;
          SHA256_BLOCK_0_start_o                    : in    std_logic
        );

end sha256_control;

architecture DEF_ARCH of sha256_control is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \padding_reg\, VCC_net_1, \padding_reg_0_0\, 
        GND_net_1, \hash_control_st_reg_i[6]_net_1\, \one_insert\, 
        \pad_one_reg_0_0\, \msg_bitlen[3]\, 
        un1_msg_bit_cnt_reg_cry_0_Y, \msg_bitlen[4]\, 
        un1_msg_bit_cnt_reg_cry_1_S, \msg_bitlen[5]\, 
        un1_msg_bit_cnt_reg_cry_2_S, \msg_bitlen[6]\, 
        un1_msg_bit_cnt_reg_cry_3_S, \msg_bitlen[7]\, 
        un1_msg_bit_cnt_reg_cry_4_S, \msg_bitlen[8]\, 
        un1_msg_bit_cnt_reg_cry_5_S, \msg_bitlen[9]\, 
        un1_msg_bit_cnt_reg_cry_6_S, \msg_bitlen[10]\, 
        un1_msg_bit_cnt_reg_cry_7_S, \msg_bitlen[11]\, 
        un1_msg_bit_cnt_reg_cry_8_S, \msg_bitlen[12]\, 
        un1_msg_bit_cnt_reg_cry_9_S, \msg_bitlen[13]\, 
        un1_msg_bit_cnt_reg_cry_10_S, \msg_bitlen[14]\, 
        un1_msg_bit_cnt_reg_cry_11_S, \msg_bitlen[15]\, 
        un1_msg_bit_cnt_reg_cry_12_S, \msg_bitlen[16]\, 
        un1_msg_bit_cnt_reg_cry_13_S, \msg_bitlen[17]\, 
        un1_msg_bit_cnt_reg_cry_14_S, \msg_bitlen[18]\, 
        un1_msg_bit_cnt_reg_cry_15_S, \msg_bitlen[19]\, 
        un1_msg_bit_cnt_reg_cry_16_S, \msg_bitlen[20]\, 
        un1_msg_bit_cnt_reg_cry_17_S, \msg_bitlen[21]\, 
        un1_msg_bit_cnt_reg_cry_18_S, \msg_bitlen[22]\, 
        un1_msg_bit_cnt_reg_cry_19_S, \msg_bitlen[23]\, 
        un1_msg_bit_cnt_reg_cry_20_S, \msg_bitlen[24]\, 
        un1_msg_bit_cnt_reg_cry_21_S, \msg_bitlen[25]\, 
        un1_msg_bit_cnt_reg_cry_22_S, \msg_bitlen[26]\, 
        un1_msg_bit_cnt_reg_cry_23_S, \msg_bitlen[27]\, 
        un1_msg_bit_cnt_reg_cry_24_S, \msg_bitlen[28]\, 
        un1_msg_bit_cnt_reg_cry_25_S, \msg_bitlen[29]\, 
        un1_msg_bit_cnt_reg_cry_26_S, \msg_bitlen[30]\, 
        un1_msg_bit_cnt_reg_cry_27_S, \msg_bitlen[31]\, 
        un1_msg_bit_cnt_reg_cry_28_S, \msg_bitlen[32]\, 
        un1_msg_bit_cnt_reg_cry_29_S, \msg_bitlen[33]\, 
        un1_msg_bit_cnt_reg_cry_30_S, \msg_bitlen[34]\, 
        un1_msg_bit_cnt_reg_cry_31_S, \msg_bitlen[35]\, 
        un1_msg_bit_cnt_reg_cry_32_S, \msg_bitlen[36]\, 
        un1_msg_bit_cnt_reg_cry_33_S, \msg_bitlen[37]\, 
        un1_msg_bit_cnt_reg_cry_34_S, \msg_bitlen[38]\, 
        un1_msg_bit_cnt_reg_cry_35_S, \msg_bitlen[39]\, 
        un1_msg_bit_cnt_reg_cry_36_S, \msg_bitlen[40]\, 
        un1_msg_bit_cnt_reg_cry_37_S, \msg_bitlen[41]\, 
        un1_msg_bit_cnt_reg_cry_38_S, \msg_bitlen[42]\, 
        un1_msg_bit_cnt_reg_cry_39_S, \msg_bitlen[43]\, 
        un1_msg_bit_cnt_reg_cry_40_S, \msg_bitlen[44]\, 
        un1_msg_bit_cnt_reg_cry_41_S, \msg_bitlen[45]\, 
        un1_msg_bit_cnt_reg_cry_42_S, \msg_bitlen[46]\, 
        un1_msg_bit_cnt_reg_cry_43_S, \msg_bitlen[47]\, 
        un1_msg_bit_cnt_reg_cry_44_S, \msg_bitlen[48]\, 
        un1_msg_bit_cnt_reg_cry_45_S, \msg_bitlen[49]\, 
        un1_msg_bit_cnt_reg_cry_46_S, \msg_bitlen[50]\, 
        un1_msg_bit_cnt_reg_cry_47_S, \msg_bitlen[51]\, 
        un1_msg_bit_cnt_reg_cry_48_S, \msg_bitlen[52]\, 
        un1_msg_bit_cnt_reg_cry_49_S, \msg_bitlen[53]\, 
        un1_msg_bit_cnt_reg_cry_50_S, \msg_bitlen[54]\, 
        un1_msg_bit_cnt_reg_cry_51_S, \msg_bitlen[55]\, 
        un1_msg_bit_cnt_reg_cry_52_S, \msg_bitlen[56]\, 
        un1_msg_bit_cnt_reg_cry_53_S, \msg_bitlen[57]\, 
        un1_msg_bit_cnt_reg_cry_54_S, \msg_bitlen[58]\, 
        un1_msg_bit_cnt_reg_cry_55_S, \msg_bitlen[59]\, 
        un1_msg_bit_cnt_reg_cry_56_S, \msg_bitlen[60]\, 
        un1_msg_bit_cnt_reg_cry_57_S, \msg_bitlen[61]\, 
        un1_msg_bit_cnt_reg_cry_58_S, \msg_bitlen[62]\, 
        un1_msg_bit_cnt_reg_cry_59_S, \msg_bitlen[63]\, 
        un1_msg_bit_cnt_reg_s_60_S, 
        \hash_control_st_reg_nsss_i_0[0]\, sha_last_blk_reg_net_1, 
        \sha_last_blk_reg_RNO\, \sha_last_blk_regce\, 
        \Kt_addr[0]\, \st_cnt_reg_s[0]\, st_cnt_rege, 
        \Kt_addr[1]\, \st_cnt_reg_s[1]\, \Kt_addr[2]\, 
        \st_cnt_reg_s[2]\, \Kt_addr[3]\, \st_cnt_reg_s[3]\, 
        \Kt_addr[4]\, \st_cnt_reg_s[4]\, \Kt_addr[5]\, 
        \st_cnt_reg_s[5]\, \st_cnt_reg[6]_net_1\, 
        \st_cnt_reg_s[6]_net_1\, \SHA256_Module_0_di_req_o\, 
        hash_control_st_reg_4, \hash_control_st_reg[0]_net_1\, 
        hash_control_st_reg_3, \SHA256_BLOCK_0_do_valid_o\, 
        hash_control_st_reg_2_0, \hash_control_st_reg_2\, 
        hash_control_st_reg_1, \hash_control_st_reg[3]_net_1\, 
        hash_control_st_reg_0, \hash_control_st_reg[4]_net_1\, 
        hash_control_st_reg, \Kt_addr_fast[1]\, \Kt_addr_1_rep1\, 
        \Kt_addr_fast[2]\, \Kt_addr_2_rep1\, \Kt_addr_0_rep2\, 
        \Kt_addr_4_rep1\, \Kt_addr_fast[3]\, st_cnt_reg_cry_cy, 
        st_cnt_clr, \st_cnt_reg_cry[0]_net_1\, 
        \st_cnt_reg_cry[1]_net_1\, \st_cnt_reg_cry[2]_net_1\, 
        \st_cnt_reg_cry[3]_net_1\, \st_cnt_reg_cry[4]_net_1\, 
        \st_cnt_reg_cry[5]_net_1\, \un1_msg_bit_cnt_reg_cry_0\, 
        \N_112\, N_115, \un1_msg_bit_cnt_reg_cry_1\, \N_223\, 
        \un1_msg_bit_cnt_reg_cry_2\, \N_361\, 
        \un1_msg_bit_cnt_reg_cry_3\, \un1_msg_bit_cnt_reg_cry_4\, 
        \un1_msg_bit_cnt_reg_cry_5\, \un1_msg_bit_cnt_reg_cry_6\, 
        \un1_msg_bit_cnt_reg_cry_7\, \un1_msg_bit_cnt_reg_cry_8\, 
        \un1_msg_bit_cnt_reg_cry_9\, \un1_msg_bit_cnt_reg_cry_10\, 
        \un1_msg_bit_cnt_reg_cry_11\, 
        \un1_msg_bit_cnt_reg_cry_12\, 
        \un1_msg_bit_cnt_reg_cry_13\, 
        \un1_msg_bit_cnt_reg_cry_14\, 
        \un1_msg_bit_cnt_reg_cry_15\, 
        \un1_msg_bit_cnt_reg_cry_16\, 
        \un1_msg_bit_cnt_reg_cry_17\, 
        \un1_msg_bit_cnt_reg_cry_18\, 
        \un1_msg_bit_cnt_reg_cry_19\, 
        \un1_msg_bit_cnt_reg_cry_20\, 
        \un1_msg_bit_cnt_reg_cry_21\, 
        \un1_msg_bit_cnt_reg_cry_22\, 
        \un1_msg_bit_cnt_reg_cry_23\, 
        \un1_msg_bit_cnt_reg_cry_24\, 
        \un1_msg_bit_cnt_reg_cry_25\, 
        \un1_msg_bit_cnt_reg_cry_26\, 
        \un1_msg_bit_cnt_reg_cry_27\, 
        \un1_msg_bit_cnt_reg_cry_28\, 
        \un1_msg_bit_cnt_reg_cry_29\, 
        \un1_msg_bit_cnt_reg_cry_30\, 
        \un1_msg_bit_cnt_reg_cry_31\, 
        \un1_msg_bit_cnt_reg_cry_32\, 
        \un1_msg_bit_cnt_reg_cry_33\, 
        \un1_msg_bit_cnt_reg_cry_34\, 
        \un1_msg_bit_cnt_reg_cry_35\, 
        \un1_msg_bit_cnt_reg_cry_36\, 
        \un1_msg_bit_cnt_reg_cry_37\, 
        \un1_msg_bit_cnt_reg_cry_38\, 
        \un1_msg_bit_cnt_reg_cry_39\, 
        \un1_msg_bit_cnt_reg_cry_40\, 
        \un1_msg_bit_cnt_reg_cry_41\, 
        \un1_msg_bit_cnt_reg_cry_42\, 
        \un1_msg_bit_cnt_reg_cry_43\, 
        \un1_msg_bit_cnt_reg_cry_44\, 
        \un1_msg_bit_cnt_reg_cry_45\, 
        \un1_msg_bit_cnt_reg_cry_46\, 
        \un1_msg_bit_cnt_reg_cry_47\, 
        \un1_msg_bit_cnt_reg_cry_48\, 
        \un1_msg_bit_cnt_reg_cry_49\, 
        \un1_msg_bit_cnt_reg_cry_50\, 
        \un1_msg_bit_cnt_reg_cry_51\, 
        \un1_msg_bit_cnt_reg_cry_52\, 
        \un1_msg_bit_cnt_reg_cry_53\, 
        \un1_msg_bit_cnt_reg_cry_54\, 
        \un1_msg_bit_cnt_reg_cry_55\, 
        \un1_msg_bit_cnt_reg_cry_56\, 
        \un1_msg_bit_cnt_reg_cry_57\, 
        \un1_msg_bit_cnt_reg_cry_58\, 
        \un1_msg_bit_cnt_reg_cry_59\, 
        \hash_control_st_reg_ns_0_0_a4_1_2[2]\, \N_102\, N_374, 
        N_114, \hash_control_st_reg_ns_i_0_a4_2_0[1]\, 
        \hash_control_st_reg_ns_0_0_a4_0[3]_net_1\, N_398, 
        oregs_ce_i_a2_0_a2_net_1, N_119, 
        \hash_control_st_reg_ns_i_0_a4_1_1[4]_net_1\, 
        \hash_control_st_reg_ns_0_0_o2_1[2]_net_1\, 
        \sha_last_blk_next_0_a4_1\, \pad_one_reg_0_0_a4_0_1\, 
        \sha_last_blk_next_0_o2_2_out_0\, N_399, N_391, N_402, 
        N_218, N_340, N_354, N_338, N_352, N_400, N_356, 
        \hash_control_st_reg_ns_i_0_0[4]_net_1\, N_355, N_369, 
        \N_111\, N_375, N_118, N_372, N_364, \pad_one_reg_0_0_0\, 
        \hash_control_st_reg_ns_i_0_1[1]_net_1\, N_220, N_373, 
        N_358, N_341 : std_logic;

begin 

    hash_control_st_reg_i(6) <= \hash_control_st_reg_i[6]_net_1\;
    msg_bitlen(63) <= \msg_bitlen[63]\;
    msg_bitlen(62) <= \msg_bitlen[62]\;
    msg_bitlen(61) <= \msg_bitlen[61]\;
    msg_bitlen(60) <= \msg_bitlen[60]\;
    msg_bitlen(59) <= \msg_bitlen[59]\;
    msg_bitlen(58) <= \msg_bitlen[58]\;
    msg_bitlen(57) <= \msg_bitlen[57]\;
    msg_bitlen(56) <= \msg_bitlen[56]\;
    msg_bitlen(55) <= \msg_bitlen[55]\;
    msg_bitlen(54) <= \msg_bitlen[54]\;
    msg_bitlen(53) <= \msg_bitlen[53]\;
    msg_bitlen(52) <= \msg_bitlen[52]\;
    msg_bitlen(51) <= \msg_bitlen[51]\;
    msg_bitlen(50) <= \msg_bitlen[50]\;
    msg_bitlen(49) <= \msg_bitlen[49]\;
    msg_bitlen(48) <= \msg_bitlen[48]\;
    msg_bitlen(47) <= \msg_bitlen[47]\;
    msg_bitlen(46) <= \msg_bitlen[46]\;
    msg_bitlen(45) <= \msg_bitlen[45]\;
    msg_bitlen(44) <= \msg_bitlen[44]\;
    msg_bitlen(43) <= \msg_bitlen[43]\;
    msg_bitlen(42) <= \msg_bitlen[42]\;
    msg_bitlen(41) <= \msg_bitlen[41]\;
    msg_bitlen(40) <= \msg_bitlen[40]\;
    msg_bitlen(39) <= \msg_bitlen[39]\;
    msg_bitlen(38) <= \msg_bitlen[38]\;
    msg_bitlen(37) <= \msg_bitlen[37]\;
    msg_bitlen(36) <= \msg_bitlen[36]\;
    msg_bitlen(35) <= \msg_bitlen[35]\;
    msg_bitlen(34) <= \msg_bitlen[34]\;
    msg_bitlen(33) <= \msg_bitlen[33]\;
    msg_bitlen(32) <= \msg_bitlen[32]\;
    msg_bitlen(31) <= \msg_bitlen[31]\;
    msg_bitlen(30) <= \msg_bitlen[30]\;
    msg_bitlen(29) <= \msg_bitlen[29]\;
    msg_bitlen(28) <= \msg_bitlen[28]\;
    msg_bitlen(27) <= \msg_bitlen[27]\;
    msg_bitlen(26) <= \msg_bitlen[26]\;
    msg_bitlen(25) <= \msg_bitlen[25]\;
    msg_bitlen(24) <= \msg_bitlen[24]\;
    msg_bitlen(23) <= \msg_bitlen[23]\;
    msg_bitlen(22) <= \msg_bitlen[22]\;
    msg_bitlen(21) <= \msg_bitlen[21]\;
    msg_bitlen(20) <= \msg_bitlen[20]\;
    msg_bitlen(19) <= \msg_bitlen[19]\;
    msg_bitlen(18) <= \msg_bitlen[18]\;
    msg_bitlen(17) <= \msg_bitlen[17]\;
    msg_bitlen(16) <= \msg_bitlen[16]\;
    msg_bitlen(15) <= \msg_bitlen[15]\;
    msg_bitlen(14) <= \msg_bitlen[14]\;
    msg_bitlen(13) <= \msg_bitlen[13]\;
    msg_bitlen(12) <= \msg_bitlen[12]\;
    msg_bitlen(11) <= \msg_bitlen[11]\;
    msg_bitlen(10) <= \msg_bitlen[10]\;
    msg_bitlen(9) <= \msg_bitlen[9]\;
    msg_bitlen(8) <= \msg_bitlen[8]\;
    msg_bitlen(7) <= \msg_bitlen[7]\;
    msg_bitlen(6) <= \msg_bitlen[6]\;
    msg_bitlen(5) <= \msg_bitlen[5]\;
    msg_bitlen(4) <= \msg_bitlen[4]\;
    msg_bitlen(3) <= \msg_bitlen[3]\;
    Kt_addr(5) <= \Kt_addr[5]\;
    Kt_addr(4) <= \Kt_addr[4]\;
    Kt_addr(3) <= \Kt_addr[3]\;
    Kt_addr(2) <= \Kt_addr[2]\;
    Kt_addr(1) <= \Kt_addr[1]\;
    Kt_addr(0) <= \Kt_addr[0]\;
    Kt_addr_fast(3) <= \Kt_addr_fast[3]\;
    Kt_addr_fast(2) <= \Kt_addr_fast[2]\;
    Kt_addr_fast(1) <= \Kt_addr_fast[1]\;
    hash_control_st_reg_2 <= \hash_control_st_reg_2\;
    one_insert <= \one_insert\;
    sha_last_blk_reg <= sha_last_blk_reg_net_1;
    SHA256_Module_0_di_req_o <= \SHA256_Module_0_di_req_o\;
    SHA256_BLOCK_0_do_valid_o <= \SHA256_BLOCK_0_do_valid_o\;
    Kt_addr_1_rep1 <= \Kt_addr_1_rep1\;
    Kt_addr_2_rep1 <= \Kt_addr_2_rep1\;
    Kt_addr_0_rep2 <= \Kt_addr_0_rep2\;
    Kt_addr_4_rep1 <= \Kt_addr_4_rep1\;
    N_112 <= \N_112\;
    N_223 <= \N_223\;
    N_361 <= \N_361\;
    N_102 <= \N_102\;
    oregs_ce_i_a2_0_a2 <= oregs_ce_i_a2_0_a2_net_1;
    sha_last_blk_next_0_o2_2_out_0 <= 
        \sha_last_blk_next_0_o2_2_out_0\;
    N_111 <= \N_111\;

    \msg_bit_cnt_reg[42]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_39_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[42]\);
    
    \hash_control_st_reg_r[3]\ : CFG4
      generic map(INIT => x"0F04")

      port map(A => N_484, B => 
        \hash_control_st_reg_ns_0_0_a4_0[3]_net_1\, C => 
        SHA256_BLOCK_0_start_o, D => N_364, Y => 
        hash_control_st_reg_0);
    
    un1_msg_bit_cnt_reg_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[17]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_13\, S => 
        un1_msg_bit_cnt_reg_cry_14_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_14\);
    
    un1_msg_bit_cnt_reg_cry_18 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[21]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_17\, S => 
        un1_msg_bit_cnt_reg_cry_18_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_18\);
    
    un1_msg_bit_cnt_reg_cry_16 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[19]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_15\, S => 
        un1_msg_bit_cnt_reg_cry_16_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_16\);
    
    un1_msg_bit_cnt_reg_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[14]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_10\, S => 
        un1_msg_bit_cnt_reg_cry_11_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_11\);
    
    \msg_bit_cnt_reg[35]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_32_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[35]\);
    
    \hash_control_st_reg_ns_i_0_o2[4]\ : CFG4
      generic map(INIT => x"C0AA")

      port map(A => N_399, B => 
        hash_control_st_reg_ns_i_0_a2_2(4), C => \Kt_addr[3]\, D
         => \Kt_addr[0]\, Y => N_118);
    
    sha_last_blk_regce : CFG4
      generic map(INIT => x"0BBB")

      port map(A => N_338, B => \N_111\, C => 
        SHA256_Module_0_waiting_data, D => 
        \hash_control_st_reg_i[6]_net_1\, Y => 
        \sha_last_blk_regce\);
    
    un1_msg_bit_cnt_reg_cry_20 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[23]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_19\, S => 
        un1_msg_bit_cnt_reg_cry_20_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_20\);
    
    \msg_bit_cnt_reg[63]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_s_60_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[63]\);
    
    \msg_bit_cnt_reg[48]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_45_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[48]\);
    
    \hash_control_st_reg_ns_i_0_a4[4]\ : CFG4
      generic map(INIT => x"4CCC")

      port map(A => \SHA256_Module_0_di_req_o\, B => N_484, C => 
        SHA256_Module_0_data_available_lastbank_8, D => state(1), 
        Y => N_356);
    
    st_cnt_reg_1_rep2 : SLE
      port map(D => \st_cnt_reg_s[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => Kt_addr_1_rep2);
    
    \msg_bit_cnt_reg[39]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_36_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[39]\);
    
    sch_ld_o_i_0_0 : CFG4
      generic map(INIT => x"DCCC")

      port map(A => \Kt_addr[0]\, B => 
        \hash_control_st_reg[4]_net_1\, C => N_399, D => N_402, Y
         => ld_i_i_3);
    
    st_cnt_reg_0_rep2 : SLE
      port map(D => \st_cnt_reg_s[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr_0_rep2\);
    
    un1_msg_bit_cnt_reg_cry_49 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[52]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_48\, S => 
        un1_msg_bit_cnt_reg_cry_49_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_49\);
    
    \st_cnt_reg_cry_cy[0]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => st_cnt_clr, C => GND_net_1, D
         => GND_net_1, FCI => VCC_net_1, S => OPEN, Y => OPEN, 
        FCO => st_cnt_reg_cry_cy);
    
    un1_msg_bit_cnt_reg_cry_57 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[60]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_56\, S => 
        un1_msg_bit_cnt_reg_cry_57_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_57\);
    
    \un1_ce_i_i_a4[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SHA256_Module_0_data_available_lastbank_8, B
         => state(1), C => N_114, Y => \N_361\);
    
    un1_msg_bit_cnt_reg_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_3\, S => 
        un1_msg_bit_cnt_reg_cry_4_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_4\);
    
    st_cnt_reg_4_rep1 : SLE
      port map(D => \st_cnt_reg_s[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr_4_rep1\);
    
    \msg_bit_cnt_reg[34]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_31_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[34]\);
    
    \hash_control_st_reg_ns_0_0_a4_0_0[6]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \SHA256_Module_0_di_req_o\, B => N_398, C => 
        \SHA256_BLOCK_0_do_valid_o\, Y => st_cnt_clr);
    
    pad_one_reg_0_0_a2 : CFG4
      generic map(INIT => x"0004")

      port map(A => \Kt_addr[1]\, B => \Kt_addr[4]\, C => 
        \Kt_addr[3]\, D => \Kt_addr[2]\, Y => N_399);
    
    \msg_bit_cnt_reg[4]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_1_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[4]\);
    
    sha_last_blk_next_0_a4_1 : CFG4
      generic map(INIT => x"0020")

      port map(A => \Kt_addr[3]\, B => \st_cnt_reg[6]_net_1\, C
         => \Kt_addr[0]\, D => \Kt_addr[4]\, Y => 
        \sha_last_blk_next_0_a4_1\);
    
    \hash_control_st_reg_ns_0_0_a4_0[2]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => N_402, B => SHA256_Module_0_waiting_data, C
         => N_118, D => N_484, Y => N_373);
    
    
        \core_error_combi_proc.core_error_combi_proc.un9_core_error_0_a2\ : 
        CFG3
      generic map(INIT => x"70")

      port map(A => SHA256_Module_0_data_available_lastbank_8, B
         => state(1), C => N_114, Y => N_400);
    
    \hash_control_st_reg[0]\ : SLE
      port map(D => hash_control_st_reg_3, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \hash_control_st_reg[0]_net_1\);
    
    \st_cnt_reg_fast[4]\ : SLE
      port map(D => \st_cnt_reg_s[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => Kt_addr_fast(4));
    
    un1_msg_bit_cnt_reg_cry_45 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[48]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_44\, S => 
        un1_msg_bit_cnt_reg_cry_45_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_45\);
    
    sch_ld_o_i_0_0_a2_0 : CFG3
      generic map(INIT => x"02")

      port map(A => \hash_control_st_reg_2\, B => \Kt_addr[5]\, C
         => \st_cnt_reg[6]_net_1\, Y => N_402);
    
    \msg_bit_cnt_reg[23]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_20_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[23]\);
    
    un1_msg_bit_cnt_reg_cry_23 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[26]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_22\, S => 
        un1_msg_bit_cnt_reg_cry_23_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_23\);
    
    \state_counter_proc.un15_ce_i_i_0_a2_RNIKNCQ\ : CFG2
      generic map(INIT => x"7")

      port map(A => N_115, B => N_398, Y => N_244_i_0);
    
    \msg_bit_cnt_reg[10]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_7_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[10]\);
    
    \hash_control_st_reg_ns_i_0_a4_1[1]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => SHA256_Module_0_waiting_data, B => 
        SHA256_Module_0_data_available_lastbank_8, C => N_391, D
         => state(1), Y => N_354);
    
    \hash_control_st_reg[3]\ : SLE
      port map(D => hash_control_st_reg_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \hash_control_st_reg[3]_net_1\);
    
    \hash_control_st_reg_nsss_i[0]\ : CFG3
      generic map(INIT => x"51")

      port map(A => SHA256_BLOCK_0_start_o, B => 
        SHA256_Module_0_waiting_data, C => 
        \hash_control_st_reg_i[6]_net_1\, Y => 
        \hash_control_st_reg_nsss_i_0[0]\);
    
    \st_cnt_reg[2]\ : SLE
      port map(D => \st_cnt_reg_s[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr[2]\);
    
    st_cnt_reg_2_rep2 : SLE
      port map(D => \st_cnt_reg_s[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => Kt_addr_2_rep2);
    
    un1_msg_bit_cnt_reg_cry_44 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[47]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_43\, S => 
        un1_msg_bit_cnt_reg_cry_44_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_44\);
    
    un1_msg_bit_cnt_reg_cry_48 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[51]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_47\, S => 
        un1_msg_bit_cnt_reg_cry_48_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_48\);
    
    un1_msg_bit_cnt_reg_cry_46 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[49]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_45\, S => 
        un1_msg_bit_cnt_reg_cry_46_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_46\);
    
    \hash_control_st_reg_ns_0_0_a4_1[2]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => \hash_control_st_reg_ns_0_0_a4_1_2[2]\, B => 
        N_115, C => \Kt_addr[4]\, D => \N_102\, Y => N_374);
    
    un1_msg_bit_cnt_reg_cry_37 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[40]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_36\, S => 
        un1_msg_bit_cnt_reg_cry_37_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_37\);
    
    un1_msg_bit_cnt_reg_cry_41 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[44]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_40\, S => 
        un1_msg_bit_cnt_reg_cry_41_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_41\);
    
    \msg_bit_cnt_reg[11]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_8_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[11]\);
    
    un1_msg_bit_cnt_reg_s_60 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[63]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_59\, S => 
        un1_msg_bit_cnt_reg_s_60_S, Y => OPEN, FCO => OPEN);
    
    \msg_bit_cnt_reg[40]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_37_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[40]\);
    
    \st_cnt_reg_fast[0]\ : SLE
      port map(D => \st_cnt_reg_s[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => Kt_addr_fast(0));
    
    \msg_bit_cnt_reg[52]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_49_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[52]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un1_msg_bit_cnt_reg_cry_29 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[32]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_28\, S => 
        un1_msg_bit_cnt_reg_cry_29_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_29\);
    
    \st_cnt_reg_cry[4]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[4]\, 
        D => GND_net_1, FCI => \st_cnt_reg_cry[3]_net_1\, S => 
        \st_cnt_reg_s[4]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[4]_net_1\);
    
    \hash_control_st_reg_ns_0_0_a4_0[3]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \N_102\, B => N_484, C => 
        \hash_control_st_reg[4]_net_1\, D => 
        \hash_control_st_reg_ns_0_0_o2_1[2]_net_1\, Y => N_364);
    
    un1_msg_bit_cnt_reg_cry_2 : ARI1
      generic map(INIT => x"5FE01")

      port map(A => \msg_bitlen[5]\, B => N_115, C => \N_361\, D
         => SHA256_Module_0_waiting_data, FCI => 
        \un1_msg_bit_cnt_reg_cry_1\, S => 
        un1_msg_bit_cnt_reg_cry_2_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_2\);
    
    \hash_control_st_reg_ns_i_0_a2_0[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \Kt_addr_fast[1]\, B => \Kt_addr_fast[2]\, Y
         => hash_control_st_reg_ns_i_0_a2_0(4));
    
    \msg_bit_cnt_reg[41]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_38_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[41]\);
    
    \msg_bit_cnt_reg[58]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_55_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[58]\);
    
    \hash_control_st_reg_ns_0_0_a4_0_0[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => SHA256_Module_0_waiting_data, B => 
        \hash_control_st_reg[3]_net_1\, Y => 
        \hash_control_st_reg_ns_0_0_a4_0[3]_net_1\);
    
    \st_cnt_reg[3]\ : SLE
      port map(D => \st_cnt_reg_s[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr[3]\);
    
    \st_cnt_reg_fast[3]\ : SLE
      port map(D => \st_cnt_reg_s[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr_fast[3]\);
    
    \msg_bit_cnt_reg[27]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_24_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[27]\);
    
    un1_msg_bit_cnt_reg_cry_25 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[28]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_24\, S => 
        un1_msg_bit_cnt_reg_cry_25_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_25\);
    
    \msg_bit_cnt_reg[26]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_23_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[26]\);
    
    \msg_bit_cnt_reg[3]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_0_Y, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[3]\);
    
    un1_msg_bit_cnt_reg_cry_24 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[27]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_23\, S => 
        un1_msg_bit_cnt_reg_cry_24_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_24\);
    
    un1_msg_bit_cnt_reg_cry_28 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[31]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_27\, S => 
        un1_msg_bit_cnt_reg_cry_28_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_28\);
    
    un1_msg_bit_cnt_reg_cry_26 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[29]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_25\, S => 
        un1_msg_bit_cnt_reg_cry_26_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_26\);
    
    \state_counter_proc.un15_ce_i_i_0_o2\ : CFG2
      generic map(INIT => x"7")

      port map(A => N_484, B => \SHA256_Module_0_di_req_o\, Y => 
        N_115);
    
    un1_msg_bit_cnt_reg_cry_21 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[24]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_20\, S => 
        un1_msg_bit_cnt_reg_cry_21_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_21\);
    
    \un1_ce_i_i_o2[0]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => bytes_sel, B => reg_17x32_0_valid_bytes_0(1), 
        C => reg_17x32_0_valid_bytes_0(0), Y => N_114);
    
    \msg_bit_cnt_reg[6]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_3_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[6]\);
    
    un1_msg_bit_cnt_reg_cry_17 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[20]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_16\, S => 
        un1_msg_bit_cnt_reg_cry_17_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_17\);
    
    \st_cnt_reg_s[6]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => 
        \st_cnt_reg[6]_net_1\, D => GND_net_1, FCI => 
        \st_cnt_reg_cry[5]_net_1\, S => \st_cnt_reg_s[6]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \hash_control_st_reg_ns_0_0_a4_1_0[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \Kt_addr[5]\, B => 
        SHA256_Module_0_waiting_data, C => \Kt_addr[0]\, Y => 
        \hash_control_st_reg_ns_i_0_a4_2_0[1]\);
    
    un1_msg_bit_cnt_reg_cry_52 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[55]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_51\, S => 
        un1_msg_bit_cnt_reg_cry_52_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_52\);
    
    \msg_bit_cnt_reg[32]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_29_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[32]\);
    
    \msg_bit_cnt_reg[25]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_22_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[25]\);
    
    \hash_control_st_reg_ns_i_0_o2_1[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \hash_control_st_reg[3]_net_1\, B => 
        sha_last_blk_reg_net_1, Y => N_119);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    st_cnt_reg_3_rep2 : SLE
      port map(D => \st_cnt_reg_s[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => Kt_addr_3_rep2);
    
    un1_msg_bit_cnt_reg_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_5\, S => 
        un1_msg_bit_cnt_reg_cry_6_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_6\);
    
    un1_msg_bit_cnt_reg_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_7\, S => 
        un1_msg_bit_cnt_reg_cry_8_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_8\);
    
    \st_cnt_reg_fast[1]\ : SLE
      port map(D => \st_cnt_reg_s[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr_fast[1]\);
    
    \msg_bit_cnt_reg[50]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_47_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[50]\);
    
    \msg_bit_cnt_reg[29]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_26_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[29]\);
    
    \st_cnt_reg_cry[2]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[2]\, 
        D => GND_net_1, FCI => \st_cnt_reg_cry[1]_net_1\, S => 
        \st_cnt_reg_s[2]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[2]_net_1\);
    
    \st_cnt_reg[5]\ : SLE
      port map(D => \st_cnt_reg_s[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr[5]\);
    
    \msg_bit_cnt_reg[38]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_35_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[38]\);
    
    \hash_control_st_reg_ns_i_0_a4_1[4]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \hash_control_st_reg_ns_i_0_a4_1_1[4]_net_1\, 
        B => SHA256_Module_0_waiting_data, C => N_118, D => N_484, 
        Y => N_358);
    
    \msg_bit_cnt_reg[13]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_10_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[13]\);
    
    \st_cnt_reg[6]\ : SLE
      port map(D => \st_cnt_reg_s[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \st_cnt_reg[6]_net_1\);
    
    \hash_control_st_reg_ns_i_0_a4_1_1[4]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \hash_control_st_reg[3]_net_1\, B => 
        \Kt_addr[5]\, C => \st_cnt_reg[6]_net_1\, Y => 
        \hash_control_st_reg_ns_i_0_a4_1_1[4]_net_1\);
    
    \msg_bit_cnt_reg[51]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_48_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[51]\);
    
    \msg_bit_cnt_reg[24]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_21_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[24]\);
    
    pad_one_reg_0_0 : CFG4
      generic map(INIT => x"ECCC")

      port map(A => N_220, B => \pad_one_reg_0_0_0\, C => 
        \one_insert\, D => \hash_control_st_reg_i[6]_net_1\, Y
         => \pad_one_reg_0_0\);
    
    \hash_control_st_reg[4]\ : SLE
      port map(D => hash_control_st_reg, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \hash_control_st_reg[4]_net_1\);
    
    \hash_control_st_reg_ns_0_0_o2_0[2]\ : CFG4
      generic map(INIT => x"F7FF")

      port map(A => \Kt_addr_2_rep1\, B => \Kt_addr_1_rep1\, C
         => \st_cnt_reg[6]_net_1\, D => \Kt_addr_fast[3]\, Y => 
        \N_102\);
    
    un1_msg_bit_cnt_reg_cry_32 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[35]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_31\, S => 
        un1_msg_bit_cnt_reg_cry_32_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_32\);
    
    \hash_control_st_reg_ns_i_0_0[4]\ : CFG4
      generic map(INIT => x"2322")

      port map(A => SHA256_Module_0_waiting_data, B => 
        \hash_control_st_reg_2\, C => N_484, D => N_218, Y => 
        \hash_control_st_reg_ns_i_0_0[4]_net_1\);
    
    \st_cnt_reg_cry[0]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[0]\, 
        D => GND_net_1, FCI => st_cnt_reg_cry_cy, S => 
        \st_cnt_reg_s[0]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[0]_net_1\);
    
    \msg_bit_cnt_reg[43]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_40_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[43]\);
    
    \hash_control_st_reg[2]\ : SLE
      port map(D => hash_control_st_reg_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \hash_control_st_reg_2\);
    
    \hash_control_st_reg_ns_i_0_1[1]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \SHA256_Module_0_di_req_o\, B => 
        SHA256_Module_0_waiting_data, C => N_354, D => N_352, Y
         => \hash_control_st_reg_ns_i_0_1[1]_net_1\);
    
    pad_one_reg_0_0_a4_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_388, B => N_402, C => 
        \hash_control_st_reg_i[6]_net_1\, D => N_399, Y => N_369);
    
    un1_msg_bit_cnt_reg_cry_47 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[50]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_46\, S => 
        un1_msg_bit_cnt_reg_cry_47_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_47\);
    
    un1_msg_bit_cnt_reg_cry_0 : ARI1
      generic map(INIT => x"5FE01")

      port map(A => \msg_bitlen[3]\, B => \N_112\, C => N_115, D
         => SHA256_Module_0_waiting_data, FCI => GND_net_1, S => 
        OPEN, Y => un1_msg_bit_cnt_reg_cry_0_Y, FCO => 
        \un1_msg_bit_cnt_reg_cry_0\);
    
    \st_cnt_reg[1]\ : SLE
      port map(D => \st_cnt_reg_s[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr[1]\);
    
    sha_last_blk_reg_RNO : CFG2
      generic map(INIT => x"B")

      port map(A => \sha_last_blk_regce\, B => 
        \hash_control_st_reg_i[6]_net_1\, Y => 
        \sha_last_blk_reg_RNO\);
    
    un1_msg_bit_cnt_reg_cry_50 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[53]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_49\, S => 
        un1_msg_bit_cnt_reg_cry_50_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_50\);
    
    sha_last_blk_next_0_o2_2_s_0 : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \Kt_addr_0_rep2\, B => \Kt_addr[5]\, C => 
        \hash_control_st_reg_2\, D => \Kt_addr_4_rep1\, Y => 
        \sha_last_blk_next_0_o2_2_out_0\);
    
    pad_one_reg : SLE
      port map(D => \pad_one_reg_0_0\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => VCC_net_1, LAT
         => GND_net_1, Q => \one_insert\);
    
    \hash_control_st_reg_ns_0_0_a4[6]\ : CFG3
      generic map(INIT => x"D0")

      port map(A => \SHA256_Module_0_di_req_o\, B => N_400, C => 
        N_391, Y => N_341);
    
    \hash_control_st_reg_ns_0_0_a4_0[5]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => SHA256_Module_0_waiting_data, B => N_484, C
         => sha_last_blk_reg_net_1, D => 
        \hash_control_st_reg[3]_net_1\, Y => N_340);
    
    \msg_bit_cnt_reg[17]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_14_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[17]\);
    
    \msg_bit_cnt_reg[16]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_13_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[16]\);
    
    un1_msg_bit_cnt_reg_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_8\, S => 
        un1_msg_bit_cnt_reg_cry_9_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_9\);
    
    \msg_bit_cnt_reg[30]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_27_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[30]\);
    
    sha_last_blk_next_0_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \one_insert\, B => \N_102\, C => 
        \sha_last_blk_next_0_o2_2_out_0\, Y => \N_111\);
    
    \hash_control_st_reg_ns_0_0_a4_1_3[2]\ : CFG4
      generic map(INIT => x"0700")

      port map(A => SHA256_Module_0_data_available_lastbank_8, B
         => state(1), C => N_114, D => 
        \hash_control_st_reg_ns_i_0_a4_2_0[1]\, Y => 
        \hash_control_st_reg_ns_0_0_a4_1_2[2]\);
    
    st_cnt_reg_4_rep2 : SLE
      port map(D => \st_cnt_reg_s[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => Kt_addr_4_rep2);
    
    oregs_ce_i_a2_0_a2_i : CFG2
      generic map(INIT => x"D")

      port map(A => \hash_control_st_reg_i[6]_net_1\, B => 
        \hash_control_st_reg[3]_net_1\, Y => N_168_i_0);
    
    \hash_control_st_reg[1]\ : SLE
      port map(D => hash_control_st_reg_2_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_do_valid_o\);
    
    \hash_control_st_reg_r[0]\ : CFG4
      generic map(INIT => x"0F08")

      port map(A => st_cnt_clr, B => oregs_ce_i_a2_0_a2_net_1, C
         => SHA256_BLOCK_0_start_o, D => N_341, Y => 
        hash_control_st_reg_3);
    
    \msg_bit_cnt_reg[31]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_28_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[31]\);
    
    st_cnt_reg_1_rep1 : SLE
      port map(D => \st_cnt_reg_s[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr_1_rep1\);
    
    \msg_bit_cnt_reg[47]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_44_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[47]\);
    
    \st_cnt_reg[4]\ : SLE
      port map(D => \st_cnt_reg_s[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr[4]\);
    
    \sha_last_blk_reg\ : SLE
      port map(D => VCC_net_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \sha_last_blk_reg_RNO\, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => \hash_control_st_reg_i[6]_net_1\, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        sha_last_blk_reg_net_1);
    
    \st_cnt_reg_cry[1]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[1]\, 
        D => GND_net_1, FCI => \st_cnt_reg_cry[0]_net_1\, S => 
        \st_cnt_reg_s[1]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[1]_net_1\);
    
    un1_msg_bit_cnt_reg_cry_30 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[33]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_29\, S => 
        un1_msg_bit_cnt_reg_cry_30_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_30\);
    
    \msg_bit_cnt_reg[46]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_43_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[46]\);
    
    st_cnt_reg_0_rep1 : SLE
      port map(D => \st_cnt_reg_s[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => Kt_addr_0_rep1);
    
    \msg_bit_cnt_reg[62]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_59_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[62]\);
    
    un1_msg_bit_cnt_reg_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[15]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_11\, S => 
        un1_msg_bit_cnt_reg_cry_12_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_12\);
    
    un1_msg_bit_cnt_reg_cry_53 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[56]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_52\, S => 
        un1_msg_bit_cnt_reg_cry_53_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_53\);
    
    padding_reg : SLE
      port map(D => \padding_reg_0_0\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \padding_reg\);
    
    sha_last_blk_next_0_a4 : CFG4
      generic map(INIT => x"0080")

      port map(A => sha_last_blk_next_0_a4_0, B => 
        \sha_last_blk_next_0_a4_1\, C => \hash_control_st_reg_2\, 
        D => \Kt_addr[5]\, Y => N_338);
    
    un1_msg_bit_cnt_reg_cry_27 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[30]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_26\, S => 
        un1_msg_bit_cnt_reg_cry_27_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_27\);
    
    \msg_bit_cnt_reg[15]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_12_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[15]\);
    
    \hash_control_st_reg_ns_i_0_a4_2[1]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \hash_control_st_reg_ns_i_0_a4_2_0[1]\, B => 
        \Kt_addr[4]\, C => N_391, D => \N_102\, Y => N_355);
    
    \st_cnt_reg_cry[3]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[3]\, 
        D => GND_net_1, FCI => \st_cnt_reg_cry[2]_net_1\, S => 
        \st_cnt_reg_s[3]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[3]_net_1\);
    
    \msg_bit_cnt_reg[53]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_50_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[53]\);
    
    \msg_bit_cnt_reg[19]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_16_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[19]\);
    
    \hash_control_st_reg_r[1]\ : CFG4
      generic map(INIT => x"0F04")

      port map(A => N_484, B => \SHA256_BLOCK_0_do_valid_o\, C
         => SHA256_BLOCK_0_start_o, D => N_340, Y => 
        hash_control_st_reg_2_0);
    
    \st_cnt_reg_fast[2]\ : SLE
      port map(D => \st_cnt_reg_s[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr_fast[2]\);
    
    un1_msg_bit_cnt_reg_cry_59 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[62]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_58\, S => 
        un1_msg_bit_cnt_reg_cry_59_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_59\);
    
    \msg_bit_cnt_reg[45]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_42_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[45]\);
    
    \msg_bit_cnt_reg[22]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_19_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[22]\);
    
    \hash_control_st_reg_r[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => N_356, B => 
        \hash_control_st_reg_ns_i_0_0[4]_net_1\, C => 
        SHA256_BLOCK_0_start_o, D => N_358, Y => 
        hash_control_st_reg_1);
    
    st_cnt_reg_2_rep1 : SLE
      port map(D => \st_cnt_reg_s[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr_2_rep1\);
    
    un1_msg_bit_cnt_reg_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_4\, S => 
        un1_msg_bit_cnt_reg_cry_5_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_5\);
    
    un1_msg_bit_cnt_reg_cry_33 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[36]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_32\, S => 
        un1_msg_bit_cnt_reg_cry_33_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_33\);
    
    \msg_bit_cnt_reg[14]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_11_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[14]\);
    
    \state_counter_proc.un15_ce_i_i_0_a2\ : CFG2
      generic map(INIT => x"1")

      port map(A => \hash_control_st_reg_2\, B => 
        \hash_control_st_reg[4]_net_1\, Y => N_398);
    
    \hash_control_st_reg_RNIM1OU[0]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => \SHA256_Module_0_di_req_o\, B => N_484, C => 
        \hash_control_st_reg[0]_net_1\, D => 
        \SHA256_BLOCK_0_do_valid_o\, Y => core_ce_o_iv_i_0);
    
    pad_one_reg_0_0_a4_0_1 : CFG3
      generic map(INIT => x"20")

      port map(A => \hash_control_st_reg_i[6]_net_1\, B => 
        \hash_control_st_reg_2\, C => \one_insert\, Y => 
        \pad_one_reg_0_0_a4_0_1\);
    
    \msg_bit_cnt_reg[49]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_46_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[49]\);
    
    \hash_control_st_reg_i[6]\ : SLE
      port map(D => \hash_control_st_reg_nsss_i_0[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \hash_control_st_reg_i[6]_net_1\);
    
    \st_cnt_reg_cry[5]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => st_cnt_clr, C => \Kt_addr[5]\, 
        D => GND_net_1, FCI => \st_cnt_reg_cry[4]_net_1\, S => 
        \st_cnt_reg_s[5]\, Y => OPEN, FCO => 
        \st_cnt_reg_cry[5]_net_1\);
    
    \oregs_ce_i_a2_0_a2\ : CFG2
      generic map(INIT => x"2")

      port map(A => \hash_control_st_reg_i[6]_net_1\, B => 
        \hash_control_st_reg[3]_net_1\, Y => 
        oregs_ce_i_a2_0_a2_net_1);
    
    un1_msg_bit_cnt_reg_cry_55 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[58]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_54\, S => 
        un1_msg_bit_cnt_reg_cry_55_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_55\);
    
    \msg_bit_cnt_reg[28]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_25_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[28]\);
    
    \hash_control_st_reg_ns_i_0_a4[1]\ : CFG4
      generic map(INIT => x"5040")

      port map(A => \SHA256_Module_0_di_req_o\, B => 
        \padding_reg\, C => \hash_control_st_reg_i[6]_net_1\, D
         => N_119, Y => N_352);
    
    un1_msg_bit_cnt_reg_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_6\, S => 
        un1_msg_bit_cnt_reg_cry_7_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_7\);
    
    un1_msg_bit_cnt_reg_cry_42 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[45]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_41\, S => 
        un1_msg_bit_cnt_reg_cry_42_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_42\);
    
    \msg_bit_cnt_reg[44]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_41_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[44]\);
    
    \hash_control_st_reg_r[5]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => SHA256_BLOCK_0_start_o, B => N_355, C => 
        N_341, D => \hash_control_st_reg_ns_i_0_1[1]_net_1\, Y
         => hash_control_st_reg_4);
    
    \hash_control_st_reg_ns_0_0_a2[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_484, B => \hash_control_st_reg_i[6]_net_1\, 
        Y => N_391);
    
    un1_msg_bit_cnt_reg_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[13]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_9\, S => 
        un1_msg_bit_cnt_reg_cry_10_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_10\);
    
    \state_counter_proc.un15_ce_i_i_0_a2_RNICG0A1\ : CFG4
      generic map(INIT => x"FF13")

      port map(A => N_398, B => SHA256_Module_0_waiting_data, C
         => N_115, D => st_cnt_clr, Y => st_cnt_rege);
    
    un1_msg_bit_cnt_reg_cry_54 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[57]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_53\, S => 
        un1_msg_bit_cnt_reg_cry_54_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_54\);
    
    \msg_bit_cnt_reg[57]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_54_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[57]\);
    
    un1_msg_bit_cnt_reg_cry_58 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[61]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_57\, S => 
        un1_msg_bit_cnt_reg_cry_58_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_58\);
    
    un1_msg_bit_cnt_reg_cry_56 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[59]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_55\, S => 
        un1_msg_bit_cnt_reg_cry_56_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_56\);
    
    un1_msg_bit_cnt_reg_cry_39 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[42]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_38\, S => 
        un1_msg_bit_cnt_reg_cry_39_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_39\);
    
    un1_msg_bit_cnt_reg_cry_51 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[54]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_50\, S => 
        un1_msg_bit_cnt_reg_cry_51_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_51\);
    
    \msg_bit_cnt_reg[60]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_57_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[60]\);
    
    un1_msg_bit_cnt_reg_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_2\, S => 
        un1_msg_bit_cnt_reg_cry_3_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_3\);
    
    \msg_bit_cnt_reg[56]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_53_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[56]\);
    
    \msg_bit_cnt_reg[5]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_2_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[5]\);
    
    \msg_bit_cnt_reg[33]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_30_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[33]\);
    
    \msg_bit_cnt_reg[61]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_58_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[61]\);
    
    un1_msg_bit_cnt_reg_cry_35 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[38]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_34\, S => 
        un1_msg_bit_cnt_reg_cry_35_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_35\);
    
    \hash_control_st_reg[5]\ : SLE
      port map(D => hash_control_st_reg_4, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_Module_0_di_req_o\);
    
    \msg_bit_cnt_reg[8]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_5_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[8]\);
    
    \hash_control_st_reg_ns_0_0_o2_1[2]\ : CFG4
      generic map(INIT => x"DFFF")

      port map(A => \Kt_addr[4]\, B => 
        SHA256_Module_0_waiting_data, C => \Kt_addr[5]\, D => 
        \Kt_addr[0]\, Y => 
        \hash_control_st_reg_ns_0_0_o2_1[2]_net_1\);
    
    \st_cnt_reg[0]\ : SLE
      port map(D => \st_cnt_reg_s[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \Kt_addr[0]\);
    
    un1_msg_bit_cnt_reg_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[16]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_12\, S => 
        un1_msg_bit_cnt_reg_cry_13_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_13\);
    
    un1_msg_bit_cnt_reg_cry_34 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[37]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_33\, S => 
        un1_msg_bit_cnt_reg_cry_34_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_34\);
    
    un1_msg_bit_cnt_reg_cry_38 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[41]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_37\, S => 
        un1_msg_bit_cnt_reg_cry_38_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_38\);
    
    un1_msg_bit_cnt_reg_cry_36 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[39]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_35\, S => 
        un1_msg_bit_cnt_reg_cry_36_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_36\);
    
    un1_msg_bit_cnt_reg_cry_31 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[34]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_30\, S => 
        un1_msg_bit_cnt_reg_cry_31_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_31\);
    
    padding_reg_0_0 : CFG4
      generic map(INIT => x"AEFF")

      port map(A => \padding_reg\, B => \hash_control_st_reg_2\, 
        C => SHA256_Module_0_waiting_data, D => 
        \hash_control_st_reg_i[6]_net_1\, Y => \padding_reg_0_0\);
    
    \msg_bit_cnt_reg[20]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_17_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[20]\);
    
    \msg_bit_cnt_reg[55]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_52_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[55]\);
    
    un1_msg_bit_cnt_reg_cry_22 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[25]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_21\, S => 
        un1_msg_bit_cnt_reg_cry_22_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_22\);
    
    
        \core_error_combi_proc.core_error_combi_proc.un9_core_error_0_a4\ : 
        CFG2
      generic map(INIT => x"4")

      port map(A => N_115, B => N_400, Y => N_375);
    
    \msg_bit_cnt_reg[7]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_4_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[7]\);
    
    un1_msg_bit_cnt_reg_cry_40 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[43]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_39\, S => 
        un1_msg_bit_cnt_reg_cry_40_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_40\);
    
    st_cnt_reg_3_rep1 : SLE
      port map(D => \st_cnt_reg_s[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => st_cnt_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => Kt_addr_3_rep1);
    
    \msg_bit_cnt_reg[59]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_56_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[59]\);
    
    \msg_bit_cnt_reg[21]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_18_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[21]\);
    
    \msg_bit_cnt_reg[9]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_6_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[9]\);
    
    \hash_control_st_reg_ns_i_0_o2_0[4]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_119, B => \padding_reg\, Y => N_218);
    
    \msg_bit_cnt_reg[37]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_34_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[37]\);
    
    un1_msg_bit_cnt_reg_cry_19 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[22]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_18\, S => 
        un1_msg_bit_cnt_reg_cry_19_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_19\);
    
    \msg_bit_cnt_reg[54]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_51_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[54]\);
    
    \msg_bit_cnt_reg[36]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_33_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[36]\);
    
    un1_msg_bit_cnt_reg_cry_1 : ARI1
      generic map(INIT => x"5FE01")

      port map(A => \msg_bitlen[4]\, B => N_115, C => \N_223\, D
         => SHA256_Module_0_waiting_data, FCI => 
        \un1_msg_bit_cnt_reg_cry_0\, S => 
        un1_msg_bit_cnt_reg_cry_1_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_1\);
    
    pad_one_reg_0_0_o2 : CFG4
      generic map(INIT => x"FFF2")

      port map(A => \SHA256_Module_0_di_req_o\, B => \N_361\, C
         => \hash_control_st_reg[4]_net_1\, D => 
        SHA256_Module_0_waiting_data, Y => N_220);
    
    pad_one_reg_0_0_0 : CFG3
      generic map(INIT => x"F8")

      port map(A => N_115, B => \pad_one_reg_0_0_a4_0_1\, C => 
        N_369, Y => \pad_one_reg_0_0_0\);
    
    \msg_bit_cnt_reg[12]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_9_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[12]\);
    
    un1_msg_bit_cnt_reg_cry_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[18]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_14\, S => 
        un1_msg_bit_cnt_reg_cry_15_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_15\);
    
    \hash_control_st_reg_ns_0_0_a4[2]\ : CFG4
      generic map(INIT => x"3020")

      port map(A => \N_102\, B => N_484, C => 
        \hash_control_st_reg[4]_net_1\, D => 
        \hash_control_st_reg_ns_0_0_o2_1[2]_net_1\, Y => N_372);
    
    \un1_ce_i_i_o4[2]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => bytes_sel, B => reg_17x32_0_valid_bytes_0(0), 
        C => SHA256_Module_0_data_available_lastbank_8, D => 
        state(1), Y => \N_112\);
    
    \hash_control_st_reg_r[4]\ : CFG4
      generic map(INIT => x"00FE")

      port map(A => N_374, B => N_373, C => N_372, D => 
        SHA256_BLOCK_0_start_o, Y => hash_control_st_reg);
    
    \un1_ce_i_i_o4[1]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => bytes_sel, B => reg_17x32_0_valid_bytes_0(1), 
        C => SHA256_Module_0_data_available_lastbank_8, D => 
        state(1), Y => \N_223\);
    
    un1_msg_bit_cnt_reg_cry_43 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \msg_bitlen[46]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un1_msg_bit_cnt_reg_cry_42\, S => 
        un1_msg_bit_cnt_reg_cry_43_S, Y => OPEN, FCO => 
        \un1_msg_bit_cnt_reg_cry_43\);
    
    \msg_bit_cnt_reg[18]\ : SLE
      port map(D => un1_msg_bit_cnt_reg_cry_15_S, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        \hash_control_st_reg_i[6]_net_1\, SD => GND_net_1, LAT
         => GND_net_1, Q => \msg_bitlen[18]\);
    
    pad_one_reg_0_0_a2_0_0 : CFG2
      generic map(INIT => x"1")

      port map(A => \Kt_addr_1_rep1\, B => \Kt_addr_2_rep1\, Y
         => pad_one_reg_0_0_a2_0);
    
    
        \core_error_combi_proc.core_error_combi_proc.un9_core_error_0\ : 
        CFG4
      generic map(INIT => x"FCFE")

      port map(A => N_391, B => N_375, C => 
        \hash_control_st_reg[0]_net_1\, D => 
        \SHA256_Module_0_di_req_o\, Y => SHA256_Module_0_error_o);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_hash_core is

    port( R1_data                              : out   std_logic_vector(31 downto 0);
          R2_data                              : out   std_logic_vector(31 downto 0);
          R3_data                              : out   std_logic_vector(31 downto 0);
          R5_data                              : out   std_logic_vector(31 downto 0);
          R6_data                              : out   std_logic_vector(31 downto 0);
          R7_data                              : out   std_logic_vector(31 downto 0);
          R0_data                              : out   std_logic_vector(31 downto 0);
          R4_data                              : out   std_logic_vector(31 downto 0);
          N4_data                              : in    std_logic_vector(31 downto 1);
          N0_data                              : in    std_logic_vector(31 downto 1);
          W_out_i_1                            : in    std_logic_vector(0 to 0);
          Kt_addr                              : in    std_logic_vector(5 to 5);
          N3_data                              : in    std_logic_vector(31 downto 1);
          N2_data                              : in    std_logic_vector(31 downto 1);
          N1_data                              : in    std_logic_vector(31 downto 1);
          N7_data                              : in    std_logic_vector(31 downto 1);
          N6_data                              : in    std_logic_vector(31 downto 1);
          N5_data                              : in    std_logic_vector(31 downto 1);
          Wt_data                              : in    std_logic_vector(31 downto 0);
          Kt_data_0                            : in    std_logic;
          Kt_data_9                            : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          core_ce_o_iv_i_0                     : in    std_logic;
          oregs_ce_i_a2_0_a2                   : in    std_logic;
          next_reg_H4_cry_0_0_Y                : in    std_logic;
          next_reg_H0_cry_0_0_Y                : in    std_logic;
          next_r0_0_cry_0_Y                    : in    std_logic;
          ld_i_i_3                             : in    std_logic;
          N_98                                 : in    std_logic;
          m34                                  : in    std_logic;
          m49_am                               : in    std_logic;
          m49_bm                               : in    std_logic;
          m62_am                               : in    std_logic;
          m62_bm                               : in    std_logic;
          m67_ns                               : in    std_logic;
          m73                                  : in    std_logic;
          m78                                  : in    std_logic;
          m83_ns                               : in    std_logic;
          m95_1_0                              : in    std_logic;
          m95_1_1                              : in    std_logic;
          m104_am                              : in    std_logic;
          m104_bm                              : in    std_logic;
          m110_ns                              : in    std_logic;
          m114                                 : in    std_logic;
          m119_ns                              : in    std_logic;
          m124                                 : in    std_logic;
          m137_am                              : in    std_logic;
          m137_bm                              : in    std_logic;
          m141                                 : in    std_logic;
          m144_ns                              : in    std_logic;
          m157                                 : in    std_logic;
          m168_1_0                             : in    std_logic;
          m168_1_1                             : in    std_logic;
          m172_ns                              : in    std_logic;
          m177                                 : in    std_logic;
          m197_1_0                             : in    std_logic;
          m197_1_1                             : in    std_logic;
          m207_1_0                             : in    std_logic;
          m207_1_1                             : in    std_logic;
          m215_am                              : in    std_logic;
          m215_bm                              : in    std_logic;
          m219                                 : in    std_logic;
          m222_ns                              : in    std_logic;
          m226_ns                              : in    std_logic;
          m230                                 : in    std_logic;
          m235_ns                              : in    std_logic;
          m239                                 : in    std_logic;
          m250_am                              : in    std_logic;
          m250_bm                              : in    std_logic;
          m254                                 : in    std_logic;
          m258_ns                              : in    std_logic;
          m273                                 : in    std_logic;
          m276_ns                              : in    std_logic;
          m281_ns                              : in    std_logic;
          m285                                 : in    std_logic;
          m289                                 : in    std_logic;
          m292_ns                              : in    std_logic;
          m296                                 : in    std_logic;
          m300_ns                              : in    std_logic;
          m304                                 : in    std_logic;
          i3_mux_1                             : in    std_logic;
          m325                                 : in    std_logic;
          m316                                 : in    std_logic;
          next_reg_H3_cry_0_0_Y                : in    std_logic;
          next_reg_H2_cry_0_0_Y                : in    std_logic;
          next_reg_H1_cry_0_0_Y                : in    std_logic;
          next_reg_H7_cry_0_0_Y                : in    std_logic;
          next_reg_H6_cry_0_0_Y                : in    std_logic;
          next_reg_H5_cry_0_0_Y                : in    std_logic;
          m10_ns                               : in    std_logic;
          m19                                  : in    std_logic
        );

end sha256_hash_core;

architecture DEF_ARCH of sha256_hash_core is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \R1_data[31]\, VCC_net_1, \next_reg_b[31]_net_1\, 
        GND_net_1, \R1_data[16]\, \next_reg_b[16]_net_1\, 
        \R1_data[17]\, \next_reg_b[17]_net_1\, \R1_data[18]\, 
        \next_reg_b[18]_net_1\, \R1_data[19]\, 
        \next_reg_b[19]_net_1\, \R1_data[20]\, 
        \next_reg_b[20]_net_1\, \R1_data[21]\, 
        \next_reg_b[21]_net_1\, \R1_data[22]\, 
        \next_reg_b[22]_net_1\, \R1_data[23]\, 
        \next_reg_b[23]_net_1\, \R1_data[24]\, 
        \next_reg_b[24]_net_1\, \R1_data[25]\, 
        \next_reg_b[25]_net_1\, \R1_data[26]\, 
        \next_reg_b[26]_net_1\, \R1_data[27]\, 
        \next_reg_b[27]_net_1\, \R1_data[28]\, 
        \next_reg_b[28]_net_1\, \R1_data[29]\, 
        \next_reg_b[29]_net_1\, \R1_data[30]\, 
        \next_reg_b[30]_net_1\, \R1_data[1]\, 
        \next_reg_b[1]_net_1\, \R1_data[2]\, 
        \next_reg_b[2]_net_1\, \R1_data[3]\, 
        \next_reg_b[3]_net_1\, \R1_data[4]\, 
        \next_reg_b[4]_net_1\, \R1_data[5]\, 
        \next_reg_b[5]_net_1\, \R1_data[6]\, 
        \next_reg_b[6]_net_1\, \R1_data[7]\, 
        \next_reg_b[7]_net_1\, \R1_data[8]\, 
        \next_reg_b[8]_net_1\, \R1_data[9]\, 
        \next_reg_b[9]_net_1\, \R1_data[10]\, 
        \next_reg_b[10]_net_1\, \R1_data[11]\, 
        \next_reg_b[11]_net_1\, \R1_data[12]\, 
        \next_reg_b[12]_net_1\, \R1_data[13]\, 
        \next_reg_b[13]_net_1\, \R1_data[14]\, 
        \next_reg_b[14]_net_1\, \R1_data[15]\, 
        \next_reg_b[15]_net_1\, \R2_data[18]\, 
        \next_reg_c[18]_net_1\, \R2_data[19]\, 
        \next_reg_c[19]_net_1\, \R2_data[20]\, 
        \next_reg_c[20]_net_1\, \R2_data[21]\, 
        \next_reg_c[21]_net_1\, \R2_data[22]\, 
        \next_reg_c[22]_net_1\, \R2_data[23]\, 
        \next_reg_c[23]_net_1\, \R2_data[24]\, 
        \next_reg_c[24]_net_1\, \R2_data[25]\, 
        \next_reg_c[25]_net_1\, \R2_data[26]\, 
        \next_reg_c[26]_net_1\, \R2_data[27]\, 
        \next_reg_c[27]_net_1\, \R2_data[28]\, 
        \next_reg_c[28]_net_1\, \R2_data[29]\, 
        \next_reg_c[29]_net_1\, \R2_data[30]\, 
        \next_reg_c[30]_net_1\, \R2_data[31]\, 
        \next_reg_c[31]_net_1\, \R1_data[0]\, 
        \next_reg_b[0]_net_1\, \R2_data[3]\, 
        \next_reg_c[3]_net_1\, \R2_data[4]\, 
        \next_reg_c[4]_net_1\, \R2_data[5]\, 
        \next_reg_c[5]_net_1\, \R2_data[6]\, 
        \next_reg_c[6]_net_1\, \R2_data[7]\, 
        \next_reg_c[7]_net_1\, \R2_data[8]\, 
        \next_reg_c[8]_net_1\, \R2_data[9]\, 
        \next_reg_c[9]_net_1\, \R2_data[10]\, 
        \next_reg_c[10]_net_1\, \R2_data[11]\, 
        \next_reg_c[11]_net_1\, \R2_data[12]\, 
        \next_reg_c[12]_net_1\, \R2_data[13]\, 
        \next_reg_c[13]_net_1\, \R2_data[14]\, 
        \next_reg_c[14]_net_1\, \R2_data[15]\, 
        \next_reg_c[15]_net_1\, \R2_data[16]\, 
        \next_reg_c[16]_net_1\, \R2_data[17]\, 
        \next_reg_c[17]_net_1\, \R3_data[20]\, 
        \next_reg_d[20]_net_1\, \R3_data[21]\, 
        \next_reg_d[21]_net_1\, \R3_data[22]\, 
        \next_reg_d[22]_net_1\, \R3_data[23]\, 
        \next_reg_d[23]_net_1\, \R3_data[24]\, 
        \next_reg_d[24]_net_1\, \R3_data[25]\, 
        \next_reg_d[25]_net_1\, \R3_data[26]\, 
        \next_reg_d[26]_net_1\, \R3_data[27]\, 
        \next_reg_d[27]_net_1\, \R3_data[28]\, 
        \next_reg_d[28]_net_1\, \R3_data[29]\, 
        \next_reg_d[29]_net_1\, \R3_data[30]\, 
        \next_reg_d[30]_net_1\, \R3_data[31]\, 
        \next_reg_d[31]_net_1\, \R2_data[0]\, 
        \next_reg_c[0]_net_1\, \R2_data[1]\, 
        \next_reg_c[1]_net_1\, \R2_data[2]\, 
        \next_reg_c[2]_net_1\, \R3_data[5]\, 
        \next_reg_d[5]_net_1\, \R3_data[6]\, 
        \next_reg_d[6]_net_1\, \R3_data[7]\, 
        \next_reg_d[7]_net_1\, \R3_data[8]\, 
        \next_reg_d[8]_net_1\, \R3_data[9]\, 
        \next_reg_d[9]_net_1\, \R3_data[10]\, 
        \next_reg_d[10]_net_1\, \R3_data[11]\, 
        \next_reg_d[11]_net_1\, \R3_data[12]\, 
        \next_reg_d[12]_net_1\, \R3_data[13]\, 
        \next_reg_d[13]_net_1\, \R3_data[14]\, 
        \next_reg_d[14]_net_1\, \R3_data[15]\, 
        \next_reg_d[15]_net_1\, \R3_data[16]\, 
        \next_reg_d[16]_net_1\, \R3_data[17]\, 
        \next_reg_d[17]_net_1\, \R3_data[18]\, 
        \next_reg_d[18]_net_1\, \R3_data[19]\, 
        \next_reg_d[19]_net_1\, \R5_data[22]\, 
        \next_reg_f[22]_net_1\, \R5_data[23]\, 
        \next_reg_f[23]_net_1\, \R5_data[24]\, 
        \next_reg_f[24]_net_1\, \R5_data[25]\, 
        \next_reg_f[25]_net_1\, \R5_data[26]\, 
        \next_reg_f[26]_net_1\, \R5_data[27]\, 
        \next_reg_f[27]_net_1\, \R5_data[28]\, 
        \next_reg_f[28]_net_1\, \R5_data[29]\, 
        \next_reg_f[29]_net_1\, \R5_data[30]\, 
        \next_reg_f[30]_net_1\, \R5_data[31]\, 
        \next_reg_f[31]_net_1\, \R3_data[0]\, 
        \next_reg_d[0]_net_1\, \R3_data[1]\, 
        \next_reg_d[1]_net_1\, \R3_data[2]\, 
        \next_reg_d[2]_net_1\, \R3_data[3]\, 
        \next_reg_d[3]_net_1\, \R3_data[4]\, 
        \next_reg_d[4]_net_1\, \R5_data[7]\, 
        \next_reg_f[7]_net_1\, \R5_data[8]\, 
        \next_reg_f[8]_net_1\, \R5_data[9]\, 
        \next_reg_f[9]_net_1\, \R5_data[10]\, 
        \next_reg_f[10]_net_1\, \R5_data[11]\, 
        \next_reg_f[11]_net_1\, \R5_data[12]\, 
        \next_reg_f[12]_net_1\, \R5_data[13]\, 
        \next_reg_f[13]_net_1\, \R5_data[14]\, 
        \next_reg_f[14]_net_1\, \R5_data[15]\, 
        \next_reg_f[15]_net_1\, \R5_data[16]\, 
        \next_reg_f[16]_net_1\, \R5_data[17]\, 
        \next_reg_f[17]_net_1\, \R5_data[18]\, 
        \next_reg_f[18]_net_1\, \R5_data[19]\, 
        \next_reg_f[19]_net_1\, \R5_data[20]\, 
        \next_reg_f[20]_net_1\, \R5_data[21]\, 
        \next_reg_f[21]_net_1\, \R6_data[24]\, 
        \next_reg_g[24]_net_1\, \R6_data[25]\, 
        \next_reg_g[25]_net_1\, \R6_data[26]\, 
        \next_reg_g[26]_net_1\, \R6_data[27]\, 
        \next_reg_g[27]_net_1\, \R6_data[28]\, 
        \next_reg_g[28]_net_1\, \R6_data[29]\, 
        \next_reg_g[29]_net_1\, \R6_data[30]\, 
        \next_reg_g[30]_net_1\, \R6_data[31]\, 
        \next_reg_g[31]_net_1\, \R5_data[0]\, 
        \next_reg_f[0]_net_1\, \R5_data[1]\, 
        \next_reg_f[1]_net_1\, \R5_data[2]\, 
        \next_reg_f[2]_net_1\, \R5_data[3]\, 
        \next_reg_f[3]_net_1\, \R5_data[4]\, 
        \next_reg_f[4]_net_1\, \R5_data[5]\, 
        \next_reg_f[5]_net_1\, \R5_data[6]\, 
        \next_reg_f[6]_net_1\, \R6_data[9]\, 
        \next_reg_g[9]_net_1\, \R6_data[10]\, 
        \next_reg_g[10]_net_1\, \R6_data[11]\, 
        \next_reg_g[11]_net_1\, \R6_data[12]\, 
        \next_reg_g[12]_net_1\, \R6_data[13]\, 
        \next_reg_g[13]_net_1\, \R6_data[14]\, 
        \next_reg_g[14]_net_1\, \R6_data[15]\, 
        \next_reg_g[15]_net_1\, \R6_data[16]\, 
        \next_reg_g[16]_net_1\, \R6_data[17]\, 
        \next_reg_g[17]_net_1\, \R6_data[18]\, 
        \next_reg_g[18]_net_1\, \R6_data[19]\, 
        \next_reg_g[19]_net_1\, \R6_data[20]\, 
        \next_reg_g[20]_net_1\, \R6_data[21]\, 
        \next_reg_g[21]_net_1\, \R6_data[22]\, 
        \next_reg_g[22]_net_1\, \R6_data[23]\, 
        \next_reg_g[23]_net_1\, \R7_data[26]\, 
        \next_reg_h[26]_net_1\, \R7_data[27]\, 
        \next_reg_h[27]_net_1\, \R7_data[28]\, 
        \next_reg_h[28]_net_1\, \R7_data[29]\, 
        \next_reg_h[29]_net_1\, \R7_data[30]\, 
        \next_reg_h[30]_net_1\, \R7_data[31]\, 
        \next_reg_h[31]_net_1\, \R6_data[0]\, 
        \next_reg_g[0]_net_1\, \R6_data[1]\, 
        \next_reg_g[1]_net_1\, \R6_data[2]\, 
        \next_reg_g[2]_net_1\, \R6_data[3]\, 
        \next_reg_g[3]_net_1\, \R6_data[4]\, 
        \next_reg_g[4]_net_1\, \R6_data[5]\, 
        \next_reg_g[5]_net_1\, \R6_data[6]\, 
        \next_reg_g[6]_net_1\, \R6_data[7]\, 
        \next_reg_g[7]_net_1\, \R6_data[8]\, 
        \next_reg_g[8]_net_1\, \R7_data[11]\, 
        \next_reg_h[11]_net_1\, \R7_data[12]\, 
        \next_reg_h[12]_net_1\, \R7_data[13]\, 
        \next_reg_h[13]_net_1\, \R7_data[14]\, 
        \next_reg_h[14]_net_1\, \R7_data[15]\, 
        \next_reg_h[15]_net_1\, \R7_data[16]\, 
        \next_reg_h[16]_net_1\, \R7_data[17]\, 
        \next_reg_h[17]_net_1\, \R7_data[18]\, 
        \next_reg_h[18]_net_1\, \R7_data[19]\, 
        \next_reg_h[19]_net_1\, \R7_data[20]\, 
        \next_reg_h[20]_net_1\, \R7_data[21]\, 
        \next_reg_h[21]_net_1\, \R7_data[22]\, 
        \next_reg_h[22]_net_1\, \R7_data[23]\, 
        \next_reg_h[23]_net_1\, \R7_data[24]\, 
        \next_reg_h[24]_net_1\, \R7_data[25]\, 
        \next_reg_h[25]_net_1\, \R0_data[28]\, \next_reg_a[28]\, 
        \R0_data[29]\, \next_reg_a[29]\, \R0_data[30]\, 
        \next_reg_a[30]\, \R0_data[31]\, \next_reg_a[31]\, 
        \R7_data[0]\, \next_reg_h[0]_net_1\, \R7_data[1]\, 
        \next_reg_h[1]_net_1\, \R7_data[2]\, 
        \next_reg_h[2]_net_1\, \R7_data[3]\, 
        \next_reg_h[3]_net_1\, \R7_data[4]\, 
        \next_reg_h[4]_net_1\, \R7_data[5]\, 
        \next_reg_h[5]_net_1\, \R7_data[6]\, 
        \next_reg_h[6]_net_1\, \R7_data[7]\, 
        \next_reg_h[7]_net_1\, \R7_data[8]\, 
        \next_reg_h[8]_net_1\, \R7_data[9]\, 
        \next_reg_h[9]_net_1\, \R7_data[10]\, 
        \next_reg_h[10]_net_1\, \R0_data[13]\, \next_reg_a[13]\, 
        \R0_data[14]\, \next_reg_a[14]\, \R0_data[15]\, 
        \next_reg_a[15]\, \R0_data[16]\, \next_reg_a[16]\, 
        \R0_data[17]\, \next_reg_a[17]\, \R0_data[18]\, 
        \next_reg_a[18]\, \R0_data[19]\, \next_reg_a[19]\, 
        \R0_data[20]\, \next_reg_a[20]\, \R0_data[21]\, 
        \next_reg_a[21]\, \R0_data[22]\, \next_reg_a[22]\, 
        \R0_data[23]\, \next_reg_a[23]\, \R0_data[24]\, 
        \next_reg_a[24]\, \R0_data[25]\, \next_reg_a[25]\, 
        \R0_data[26]\, \next_reg_a[26]\, \R0_data[27]\, 
        \next_reg_a[27]\, \R4_data[30]\, \next_reg_e[30]\, 
        \R4_data[31]\, \next_reg_e[31]\, \R0_data[0]\, 
        next_reg_a_cry_0_0_Y, \R0_data[1]\, \next_reg_a[1]\, 
        \R0_data[2]\, \next_reg_a[2]\, \R0_data[3]\, 
        \next_reg_a[3]\, \R0_data[4]\, \next_reg_a[4]\, 
        \R0_data[5]\, \next_reg_a[5]\, \R0_data[6]\, 
        \next_reg_a[6]\, \R0_data[7]\, \next_reg_a[7]\, 
        \R0_data[8]\, \next_reg_a[8]\, \R0_data[9]\, 
        \next_reg_a[9]\, \R0_data[10]\, \next_reg_a[10]\, 
        \R0_data[11]\, \next_reg_a[11]\, \R0_data[12]\, 
        \next_reg_a[12]\, \R4_data[15]\, \next_reg_e[15]\, 
        \R4_data[16]\, \next_reg_e[16]\, \R4_data[17]\, 
        \next_reg_e[17]\, \R4_data[18]\, \next_reg_e[18]\, 
        \R4_data[19]\, \next_reg_e[19]\, \R4_data[20]\, 
        \next_reg_e[20]\, \R4_data[21]\, \next_reg_e[21]\, 
        \R4_data[22]\, \next_reg_e[22]\, \R4_data[23]\, 
        \next_reg_e[23]\, \R4_data[24]\, \next_reg_e[24]\, 
        \R4_data[25]\, \next_reg_e[25]\, \R4_data[26]\, 
        \next_reg_e[26]\, \R4_data[27]\, \next_reg_e[27]\, 
        \R4_data[28]\, \next_reg_e[28]\, \R4_data[29]\, 
        \next_reg_e[29]\, \R4_data[0]\, next_reg_e_cry_0_0_Y, 
        \R4_data[1]\, \next_reg_e[1]\, \R4_data[2]\, 
        \next_reg_e[2]\, \R4_data[3]\, \next_reg_e[3]\, 
        \R4_data[4]\, \next_reg_e[4]\, \R4_data[5]\, 
        \next_reg_e[5]\, \R4_data[6]\, \next_reg_e[6]\, 
        \R4_data[7]\, \next_reg_e[7]\, \R4_data[8]\, 
        \next_reg_e[8]\, \R4_data[9]\, \next_reg_e[9]\, 
        \R4_data[10]\, \next_reg_e[10]\, \R4_data[11]\, 
        \next_reg_e[11]\, \R4_data[12]\, \next_reg_e[12]\, 
        \R4_data[13]\, \next_reg_e[13]\, \R4_data[14]\, 
        \next_reg_e[14]\, next_reg_e_cry_0, sum3_cry_0_Y, 
        next_reg_e_cry_1, \sum3[1]\, next_reg_e_cry_2, \sum3[2]\, 
        next_reg_e_cry_3, \sum3[3]\, next_reg_e_cry_4, \sum3[4]\, 
        next_reg_e_cry_5, \sum3[5]\, next_reg_e_cry_6, \sum3[6]\, 
        next_reg_e_cry_7, \sum3[7]\, next_reg_e_cry_8, \sum3[8]\, 
        next_reg_e_cry_9, \sum3[9]\, next_reg_e_cry_10, 
        \sum3[10]\, next_reg_e_cry_11, \sum3[11]\, 
        next_reg_e_cry_12, \sum3[12]\, next_reg_e_cry_13, 
        \sum3[13]\, next_reg_e_cry_14, \sum3[14]\, 
        next_reg_e_cry_15, \sum3[15]\, next_reg_e_cry_16, 
        \sum3[16]\, next_reg_e_cry_17, \sum3[17]\, 
        next_reg_e_cry_18, \sum3[18]\, next_reg_e_cry_19, 
        \sum3[19]\, next_reg_e_cry_20, \sum3[20]\, 
        next_reg_e_cry_21, \sum3[21]\, next_reg_e_cry_22, 
        \sum3[22]\, next_reg_e_cry_23, \sum3[23]\, 
        next_reg_e_cry_24, \sum3[24]\, next_reg_e_cry_25, 
        \sum3[25]\, next_reg_e_cry_26, \sum3[26]\, 
        next_reg_e_cry_27, \sum3[27]\, next_reg_e_cry_28, 
        \sum3[28]\, next_reg_e_cry_29, \sum3[29]\, \sum3[31]\, 
        next_reg_e_cry_30, \sum3[30]\, next_reg_a_cry_0, 
        sum0_4_cry_0_Y_0, next_reg_a_cry_1, \sum0_4[1]\, 
        next_reg_a_cry_2, \sum0_4[2]\, next_reg_a_cry_3, 
        \sum0_4[3]\, next_reg_a_cry_4, \sum0_4[4]\, 
        next_reg_a_cry_5, \sum0_4[5]\, next_reg_a_cry_6, 
        \sum0_4[6]\, next_reg_a_cry_7, \sum0_4[7]\, 
        next_reg_a_cry_8, \sum0_4[8]\, next_reg_a_cry_9, 
        \sum0_4[9]\, next_reg_a_cry_10, \sum0_4[10]\, 
        next_reg_a_cry_11, \sum0_4[11]\, next_reg_a_cry_12, 
        \sum0_4[12]\, next_reg_a_cry_13, \sum0_4[13]\, 
        next_reg_a_cry_14, \sum0_4[14]\, next_reg_a_cry_15, 
        \sum0_4[15]\, next_reg_a_cry_16, \sum0_4[16]\, 
        next_reg_a_cry_17, \sum0_4[17]\, next_reg_a_cry_18, 
        \sum0_4[18]\, next_reg_a_cry_19, \sum0_4[19]\, 
        next_reg_a_cry_20, \sum0_4[20]\, next_reg_a_cry_21, 
        \sum0_4[21]\, next_reg_a_cry_22, \sum0_4[22]\, 
        next_reg_a_cry_23, \sum0_4[23]\, next_reg_a_cry_24, 
        \sum0_4[24]\, next_reg_a_cry_25, \sum0_4[25]\, 
        next_reg_a_cry_26, \sum0_4[26]\, next_reg_a_cry_27, 
        \sum0_4[27]\, next_reg_a_cry_28, \sum0_4[28]\, 
        next_reg_a_cry_29, \sum0_4[29]\, \sum0_4[31]\, 
        next_reg_a_cry_30, \sum0_4[30]\, \sum0_4_cry_0\, sum0_4_0, 
        \sum0_4[0]\, \sum0_4_cry_1\, \SIG0_0[1]\, \sum0_4_axb_1\, 
        \sum0_4_cry_2\, \SIG0_0[2]\, \sum0_4_axb_2\, 
        \sum0_4_cry_3\, \SIG0_0[3]\, \sum0_4_axb_3\, 
        \sum0_4_cry_4\, \SIG0_0[4]\, \sum0_4_axb_4\, 
        \sum0_4_cry_5\, \SIG0_0[5]\, \sum0_4_axb_5\, 
        \sum0_4_cry_6\, \SIG0_0[6]\, \sum0_4_axb_6\, 
        \sum0_4_cry_7\, \SIG0_0[7]\, \sum0_4_axb_7\, 
        \sum0_4_cry_8\, \SIG0_0[8]\, \sum0_4_axb_8\, 
        \sum0_4_cry_9\, \SIG0_0[9]\, \sum0_4_axb_9\, 
        \sum0_4_cry_10\, \SIG0_0[10]\, \sum0_4_axb_10\, 
        \sum0_4_cry_11\, \SIG0_0[11]\, \sum0_4_axb_11\, 
        \sum0_4_cry_12\, \SIG0_0[12]\, \sum0_4_axb_12\, 
        \sum0_4_cry_13\, \SIG0_0[13]\, \sum0_4_axb_13\, 
        \sum0_4_cry_14\, \SIG0_0[14]\, \sum0_4_axb_14\, 
        \sum0_4_cry_15\, \SIG0_0[15]\, \sum0_4_axb_15\, 
        \sum0_4_cry_16\, \SIG0_0[16]\, \sum0_4_axb_16\, 
        \sum0_4_cry_17\, \SIG0_0[17]\, \sum0_4_axb_17\, 
        \sum0_4_cry_18\, \SIG0_0[18]\, \sum0_4_axb_18\, 
        \sum0_4_cry_19\, \SIG0_0[19]\, \sum0_4_axb_19\, 
        \sum0_4_cry_20\, \SIG0_0[20]\, \sum0_4_axb_20\, 
        \sum0_4_cry_21\, \SIG0_0[21]\, \sum0_4_axb_21\, 
        \sum0_4_cry_22\, \SIG0_0[22]\, \sum0_4_axb_22\, 
        \sum0_4_cry_23\, \SIG0_0[23]\, \sum0_4_axb_23\, 
        \sum0_4_cry_24\, \SIG0_0[24]\, \sum0_4_axb_24\, 
        \sum0_4_cry_25\, \SIG0_0[25]\, \sum0_4_axb_25\, 
        \sum0_4_cry_26\, \SIG0_0[26]\, \sum0_4_axb_26\, 
        \sum0_4_cry_27\, \SIG0_0[27]\, \sum0_4_axb_27\, 
        \sum0_4_cry_28\, \SIG0_0[28]\, \sum0_4_axb_28\, 
        \sum0_4_cry_29\, \SIG0_0[29]\, \sum0_4_axb_29\, 
        \Maj[31]_net_1\, \sum0_4_cry_30\, \SIG0_0[30]\, 
        \sum0_4_axb_30\, \sum3_6_cry_0\, sum3_6_cry_0_Y, 
        sum3_6_0_cry_0_Y, \sum3_6_cry_1\, \sum3_6[1]\, 
        \sum3_6_0[1]\, \sum3_6_cry_2\, \sum3_6[2]\, \sum3_6_0[2]\, 
        \sum3_6_cry_3\, \sum3_6[3]\, \sum3_6_0[3]\, 
        \sum3_6_cry_4\, \sum3_6[4]\, \sum3_6_0[4]\, 
        \sum3_6_cry_5\, \sum3_6[5]\, \sum3_6_0[5]\, 
        \sum3_6_cry_6\, \sum3_6[6]\, \sum3_6_0[6]\, 
        \sum3_6_cry_7\, \sum3_6[7]\, \sum3_6_0[7]\, 
        \sum3_6_cry_8\, \sum3_6[8]\, \sum3_6_0[8]\, 
        \sum3_6_cry_9\, \sum3_6[9]\, \sum3_6_0[9]\, 
        \sum3_6_cry_10\, \sum3_6[10]\, \sum3_6_0[10]\, 
        \sum3_6_cry_11\, \sum3_6[11]\, \sum3_6_0[11]\, 
        \sum3_6_cry_12\, \sum3_6[12]\, \sum3_6_0[12]\, 
        \sum3_6_cry_13\, \sum3_6[13]\, \sum3_6_0[13]\, 
        \sum3_6_cry_14\, \sum3_6[14]\, \sum3_6_0[14]\, 
        \sum3_6_cry_15\, \sum3_6[15]\, \sum3_6_0[15]\, 
        \sum3_6_cry_16\, \sum3_6[16]\, \sum3_6_0[16]\, 
        \sum3_6_cry_17\, \sum3_6[17]\, \sum3_6_0[17]\, 
        \sum3_6_cry_18\, \sum3_6[18]\, \sum3_6_0[18]\, 
        \sum3_6_cry_19\, \sum3_6[19]\, \sum3_6_0[19]\, 
        \sum3_6_cry_20\, \sum3_6[20]\, \sum3_6_0[20]\, 
        \sum3_6_cry_21\, \sum3_6[21]\, \sum3_6_0[21]\, 
        \sum3_6_cry_22\, \sum3_6[22]\, \sum3_6_0[22]\, 
        \sum3_6_cry_23\, \sum3_6[23]\, \sum3_6_0[23]\, 
        \sum3_6_cry_24\, \sum3_6[24]\, \sum3_6_0[24]\, 
        \sum3_6_cry_25\, \sum3_6[25]\, \sum3_6_0[25]\, 
        \sum3_6_cry_26\, \sum3_6[26]\, \sum3_6_0[26]\, 
        \sum3_6_cry_27\, \sum3_6[27]\, \sum3_6_0[27]\, 
        \sum3_6_cry_28\, \sum3_6[28]\, \sum3_6_0[28]\, 
        \sum3_6_cry_29\, \sum3_6[29]\, \sum3_6_0[29]\, 
        \sum3_6[31]\, \sum3_6_0[31]\, \sum3_6_cry_30\, 
        \sum3_6[30]\, \sum3_6_0[30]\, \sum3_6_0_cry_0\, 
        \sum3_6_0_cry_1\, \sum3_6_0_cry_2\, \sum3_6_0_cry_3\, 
        \sum3_6_0_cry_4\, \sum3_6_0_cry_5\, \sum3_6_0_cry_6\, 
        \sum3_6_0_cry_7\, \sum3_6_0_cry_8\, \sum3_6_0_cry_9\, 
        \sum3_6_0_cry_10\, \sum3_6_0_cry_11\, \sum3_6_0_cry_12\, 
        \sum3_6_0_cry_13\, \sum3_6_0_cry_14\, \sum3_6_0_cry_15\, 
        \sum3_6_0_cry_16\, \sum3_6_0_cry_17\, \sum3_6_0_cry_18\, 
        \sum3_6_0_cry_19\, \sum3_6_0_cry_20\, \sum3_6_0_cry_21\, 
        \sum3_6_0_cry_22\, \sum3_6_0_cry_23\, \sum3_6_0_cry_24\, 
        \sum3_6_0_cry_25\, \sum3_6_0_cry_26\, \sum3_6_0_cry_27\, 
        \sum3_6_0_cry_28\, \sum3_6_0_cry_29\, \sum3_6_0_cry_30\, 
        \sum3_cry_0\, \Wt_data_0[0]\, \sum3[0]\, \sum3_cry_1\, 
        \sum3_4[1]\, \sum3_cry_2\, \sum3_4[2]\, \sum3_cry_3\, 
        \sum3_4[3]\, \sum3_cry_4\, \sum3_4[4]\, \sum3_cry_5\, 
        \sum3_4[5]\, \sum3_cry_6\, \sum3_4[6]\, \sum3_cry_7\, 
        \sum3_4[7]\, \sum3_cry_8\, \sum3_4[8]\, \sum3_cry_9\, 
        \sum3_4[9]\, \sum3_cry_10\, \sum3_4[10]\, \sum3_cry_11\, 
        \sum3_4[11]\, \sum3_cry_12\, \sum3_4[12]\, \sum3_cry_13\, 
        \sum3_4[13]\, \sum3_cry_14\, \sum3_4[14]\, \sum3_cry_15\, 
        \sum3_4[15]\, \sum3_cry_16\, \sum3_4[16]\, \sum3_cry_17\, 
        \sum3_4[17]\, \sum3_cry_18\, \sum3_4[18]\, \sum3_cry_19\, 
        \sum3_4[19]\, \sum3_cry_20\, \sum3_4[20]\, \sum3_cry_21\, 
        \sum3_4[21]\, \sum3_cry_22\, \sum3_4[22]\, \sum3_cry_23\, 
        \sum3_4[23]\, \sum3_cry_24\, \sum3_4[24]\, \sum3_cry_25\, 
        \sum3_4[25]\, \sum3_cry_26\, \sum3_4[26]\, \sum3_cry_27\, 
        \sum3_4[27]\, \sum3_cry_28\, \sum3_4[28]\, \sum3_cry_29\, 
        \sum3_4[29]\, \sum3_4[31]\, \sum3_cry_30\, \sum3_4[30]\, 
        \sum3_4_cry_0\, sum3_4_cry_0_Y, sum3_4_0, \sum3_4[0]\, 
        \sum3_4_cry_1\, \sum3_4_cry_2\, \sum3_4_cry_3\, 
        \sum3_4_cry_4\, \sum3_4_cry_5\, \sum3_4_cry_6\, 
        \sum3_4_cry_7\, \sum3_4_cry_8\, \sum3_4_cry_9\, 
        \sum3_4_cry_10\, \sum3_4_cry_11\, \sum3_4_cry_12\, 
        \sum3_4_cry_13\, \sum3_4_cry_14\, \sum3_4_cry_15\, 
        \sum3_4_cry_16\, \sum3_4_cry_17\, \sum3_4_cry_18\, 
        \sum3_4_cry_19\, \sum3_4_cry_20\, \sum3_4_cry_21\, 
        \sum3_4_cry_22\, \sum3_4_cry_23\, \sum3_4_cry_24\, 
        \sum3_4_cry_25\, \sum3_4_cry_26\, \sum3_4_cry_27\, 
        \sum3_4_cry_28\, \sum3_4_cry_29\, \sum3_4_cry_30\, 
        \SIG0[13]_net_1\, \SIG0[3]_net_1\, \SIG0[1]_net_1\, 
        \SIG0[24]_net_1\, \SIG0[22]_net_1\, sum0_4, 
        \SIG0[11]_net_1\, \SIG0[10]_net_1\, \SIG0[9]_net_1\, 
        \SIG0[21]_net_1\, \SIG0[8]_net_1\, \SIG0[5]_net_1\, 
        \SIG0[26]_net_1\, \SIG0[20]_net_1\, \SIG0[17]_net_1\, 
        \SIG0[7]_net_1\, \SIG0[6]_net_1\, \SIG0[4]_net_1\, 
        \SIG0[29]_net_1\, \SIG0[28]_net_1\, \SIG0[27]_net_1\, 
        \SIG0[18]_net_1\, \SIG0[16]_net_1\, \SIG0[19]_net_1\, 
        \SIG0[23]_net_1\, \SIG0[25]_net_1\, \SIG0[30]_net_1\, 
        \SIG0[2]_net_1\, \SIG0[12]_net_1\, \SIG0[14]_net_1\, 
        \SIG0[15]_net_1\ : std_logic;

begin 

    R1_data(31) <= \R1_data[31]\;
    R1_data(30) <= \R1_data[30]\;
    R1_data(29) <= \R1_data[29]\;
    R1_data(28) <= \R1_data[28]\;
    R1_data(27) <= \R1_data[27]\;
    R1_data(26) <= \R1_data[26]\;
    R1_data(25) <= \R1_data[25]\;
    R1_data(24) <= \R1_data[24]\;
    R1_data(23) <= \R1_data[23]\;
    R1_data(22) <= \R1_data[22]\;
    R1_data(21) <= \R1_data[21]\;
    R1_data(20) <= \R1_data[20]\;
    R1_data(19) <= \R1_data[19]\;
    R1_data(18) <= \R1_data[18]\;
    R1_data(17) <= \R1_data[17]\;
    R1_data(16) <= \R1_data[16]\;
    R1_data(15) <= \R1_data[15]\;
    R1_data(14) <= \R1_data[14]\;
    R1_data(13) <= \R1_data[13]\;
    R1_data(12) <= \R1_data[12]\;
    R1_data(11) <= \R1_data[11]\;
    R1_data(10) <= \R1_data[10]\;
    R1_data(9) <= \R1_data[9]\;
    R1_data(8) <= \R1_data[8]\;
    R1_data(7) <= \R1_data[7]\;
    R1_data(6) <= \R1_data[6]\;
    R1_data(5) <= \R1_data[5]\;
    R1_data(4) <= \R1_data[4]\;
    R1_data(3) <= \R1_data[3]\;
    R1_data(2) <= \R1_data[2]\;
    R1_data(1) <= \R1_data[1]\;
    R1_data(0) <= \R1_data[0]\;
    R2_data(31) <= \R2_data[31]\;
    R2_data(30) <= \R2_data[30]\;
    R2_data(29) <= \R2_data[29]\;
    R2_data(28) <= \R2_data[28]\;
    R2_data(27) <= \R2_data[27]\;
    R2_data(26) <= \R2_data[26]\;
    R2_data(25) <= \R2_data[25]\;
    R2_data(24) <= \R2_data[24]\;
    R2_data(23) <= \R2_data[23]\;
    R2_data(22) <= \R2_data[22]\;
    R2_data(21) <= \R2_data[21]\;
    R2_data(20) <= \R2_data[20]\;
    R2_data(19) <= \R2_data[19]\;
    R2_data(18) <= \R2_data[18]\;
    R2_data(17) <= \R2_data[17]\;
    R2_data(16) <= \R2_data[16]\;
    R2_data(15) <= \R2_data[15]\;
    R2_data(14) <= \R2_data[14]\;
    R2_data(13) <= \R2_data[13]\;
    R2_data(12) <= \R2_data[12]\;
    R2_data(11) <= \R2_data[11]\;
    R2_data(10) <= \R2_data[10]\;
    R2_data(9) <= \R2_data[9]\;
    R2_data(8) <= \R2_data[8]\;
    R2_data(7) <= \R2_data[7]\;
    R2_data(6) <= \R2_data[6]\;
    R2_data(5) <= \R2_data[5]\;
    R2_data(4) <= \R2_data[4]\;
    R2_data(3) <= \R2_data[3]\;
    R2_data(2) <= \R2_data[2]\;
    R2_data(1) <= \R2_data[1]\;
    R2_data(0) <= \R2_data[0]\;
    R3_data(31) <= \R3_data[31]\;
    R3_data(30) <= \R3_data[30]\;
    R3_data(29) <= \R3_data[29]\;
    R3_data(28) <= \R3_data[28]\;
    R3_data(27) <= \R3_data[27]\;
    R3_data(26) <= \R3_data[26]\;
    R3_data(25) <= \R3_data[25]\;
    R3_data(24) <= \R3_data[24]\;
    R3_data(23) <= \R3_data[23]\;
    R3_data(22) <= \R3_data[22]\;
    R3_data(21) <= \R3_data[21]\;
    R3_data(20) <= \R3_data[20]\;
    R3_data(19) <= \R3_data[19]\;
    R3_data(18) <= \R3_data[18]\;
    R3_data(17) <= \R3_data[17]\;
    R3_data(16) <= \R3_data[16]\;
    R3_data(15) <= \R3_data[15]\;
    R3_data(14) <= \R3_data[14]\;
    R3_data(13) <= \R3_data[13]\;
    R3_data(12) <= \R3_data[12]\;
    R3_data(11) <= \R3_data[11]\;
    R3_data(10) <= \R3_data[10]\;
    R3_data(9) <= \R3_data[9]\;
    R3_data(8) <= \R3_data[8]\;
    R3_data(7) <= \R3_data[7]\;
    R3_data(6) <= \R3_data[6]\;
    R3_data(5) <= \R3_data[5]\;
    R3_data(4) <= \R3_data[4]\;
    R3_data(3) <= \R3_data[3]\;
    R3_data(2) <= \R3_data[2]\;
    R3_data(1) <= \R3_data[1]\;
    R3_data(0) <= \R3_data[0]\;
    R5_data(31) <= \R5_data[31]\;
    R5_data(30) <= \R5_data[30]\;
    R5_data(29) <= \R5_data[29]\;
    R5_data(28) <= \R5_data[28]\;
    R5_data(27) <= \R5_data[27]\;
    R5_data(26) <= \R5_data[26]\;
    R5_data(25) <= \R5_data[25]\;
    R5_data(24) <= \R5_data[24]\;
    R5_data(23) <= \R5_data[23]\;
    R5_data(22) <= \R5_data[22]\;
    R5_data(21) <= \R5_data[21]\;
    R5_data(20) <= \R5_data[20]\;
    R5_data(19) <= \R5_data[19]\;
    R5_data(18) <= \R5_data[18]\;
    R5_data(17) <= \R5_data[17]\;
    R5_data(16) <= \R5_data[16]\;
    R5_data(15) <= \R5_data[15]\;
    R5_data(14) <= \R5_data[14]\;
    R5_data(13) <= \R5_data[13]\;
    R5_data(12) <= \R5_data[12]\;
    R5_data(11) <= \R5_data[11]\;
    R5_data(10) <= \R5_data[10]\;
    R5_data(9) <= \R5_data[9]\;
    R5_data(8) <= \R5_data[8]\;
    R5_data(7) <= \R5_data[7]\;
    R5_data(6) <= \R5_data[6]\;
    R5_data(5) <= \R5_data[5]\;
    R5_data(4) <= \R5_data[4]\;
    R5_data(3) <= \R5_data[3]\;
    R5_data(2) <= \R5_data[2]\;
    R5_data(1) <= \R5_data[1]\;
    R5_data(0) <= \R5_data[0]\;
    R6_data(31) <= \R6_data[31]\;
    R6_data(30) <= \R6_data[30]\;
    R6_data(29) <= \R6_data[29]\;
    R6_data(28) <= \R6_data[28]\;
    R6_data(27) <= \R6_data[27]\;
    R6_data(26) <= \R6_data[26]\;
    R6_data(25) <= \R6_data[25]\;
    R6_data(24) <= \R6_data[24]\;
    R6_data(23) <= \R6_data[23]\;
    R6_data(22) <= \R6_data[22]\;
    R6_data(21) <= \R6_data[21]\;
    R6_data(20) <= \R6_data[20]\;
    R6_data(19) <= \R6_data[19]\;
    R6_data(18) <= \R6_data[18]\;
    R6_data(17) <= \R6_data[17]\;
    R6_data(16) <= \R6_data[16]\;
    R6_data(15) <= \R6_data[15]\;
    R6_data(14) <= \R6_data[14]\;
    R6_data(13) <= \R6_data[13]\;
    R6_data(12) <= \R6_data[12]\;
    R6_data(11) <= \R6_data[11]\;
    R6_data(10) <= \R6_data[10]\;
    R6_data(9) <= \R6_data[9]\;
    R6_data(8) <= \R6_data[8]\;
    R6_data(7) <= \R6_data[7]\;
    R6_data(6) <= \R6_data[6]\;
    R6_data(5) <= \R6_data[5]\;
    R6_data(4) <= \R6_data[4]\;
    R6_data(3) <= \R6_data[3]\;
    R6_data(2) <= \R6_data[2]\;
    R6_data(1) <= \R6_data[1]\;
    R6_data(0) <= \R6_data[0]\;
    R7_data(31) <= \R7_data[31]\;
    R7_data(30) <= \R7_data[30]\;
    R7_data(29) <= \R7_data[29]\;
    R7_data(28) <= \R7_data[28]\;
    R7_data(27) <= \R7_data[27]\;
    R7_data(26) <= \R7_data[26]\;
    R7_data(25) <= \R7_data[25]\;
    R7_data(24) <= \R7_data[24]\;
    R7_data(23) <= \R7_data[23]\;
    R7_data(22) <= \R7_data[22]\;
    R7_data(21) <= \R7_data[21]\;
    R7_data(20) <= \R7_data[20]\;
    R7_data(19) <= \R7_data[19]\;
    R7_data(18) <= \R7_data[18]\;
    R7_data(17) <= \R7_data[17]\;
    R7_data(16) <= \R7_data[16]\;
    R7_data(15) <= \R7_data[15]\;
    R7_data(14) <= \R7_data[14]\;
    R7_data(13) <= \R7_data[13]\;
    R7_data(12) <= \R7_data[12]\;
    R7_data(11) <= \R7_data[11]\;
    R7_data(10) <= \R7_data[10]\;
    R7_data(9) <= \R7_data[9]\;
    R7_data(8) <= \R7_data[8]\;
    R7_data(7) <= \R7_data[7]\;
    R7_data(6) <= \R7_data[6]\;
    R7_data(5) <= \R7_data[5]\;
    R7_data(4) <= \R7_data[4]\;
    R7_data(3) <= \R7_data[3]\;
    R7_data(2) <= \R7_data[2]\;
    R7_data(1) <= \R7_data[1]\;
    R7_data(0) <= \R7_data[0]\;
    R0_data(31) <= \R0_data[31]\;
    R0_data(30) <= \R0_data[30]\;
    R0_data(29) <= \R0_data[29]\;
    R0_data(28) <= \R0_data[28]\;
    R0_data(27) <= \R0_data[27]\;
    R0_data(26) <= \R0_data[26]\;
    R0_data(25) <= \R0_data[25]\;
    R0_data(24) <= \R0_data[24]\;
    R0_data(23) <= \R0_data[23]\;
    R0_data(22) <= \R0_data[22]\;
    R0_data(21) <= \R0_data[21]\;
    R0_data(20) <= \R0_data[20]\;
    R0_data(19) <= \R0_data[19]\;
    R0_data(18) <= \R0_data[18]\;
    R0_data(17) <= \R0_data[17]\;
    R0_data(16) <= \R0_data[16]\;
    R0_data(15) <= \R0_data[15]\;
    R0_data(14) <= \R0_data[14]\;
    R0_data(13) <= \R0_data[13]\;
    R0_data(12) <= \R0_data[12]\;
    R0_data(11) <= \R0_data[11]\;
    R0_data(10) <= \R0_data[10]\;
    R0_data(9) <= \R0_data[9]\;
    R0_data(8) <= \R0_data[8]\;
    R0_data(7) <= \R0_data[7]\;
    R0_data(6) <= \R0_data[6]\;
    R0_data(5) <= \R0_data[5]\;
    R0_data(4) <= \R0_data[4]\;
    R0_data(3) <= \R0_data[3]\;
    R0_data(2) <= \R0_data[2]\;
    R0_data(1) <= \R0_data[1]\;
    R0_data(0) <= \R0_data[0]\;
    R4_data(31) <= \R4_data[31]\;
    R4_data(30) <= \R4_data[30]\;
    R4_data(29) <= \R4_data[29]\;
    R4_data(28) <= \R4_data[28]\;
    R4_data(27) <= \R4_data[27]\;
    R4_data(26) <= \R4_data[26]\;
    R4_data(25) <= \R4_data[25]\;
    R4_data(24) <= \R4_data[24]\;
    R4_data(23) <= \R4_data[23]\;
    R4_data(22) <= \R4_data[22]\;
    R4_data(21) <= \R4_data[21]\;
    R4_data(20) <= \R4_data[20]\;
    R4_data(19) <= \R4_data[19]\;
    R4_data(18) <= \R4_data[18]\;
    R4_data(17) <= \R4_data[17]\;
    R4_data(16) <= \R4_data[16]\;
    R4_data(15) <= \R4_data[15]\;
    R4_data(14) <= \R4_data[14]\;
    R4_data(13) <= \R4_data[13]\;
    R4_data(12) <= \R4_data[12]\;
    R4_data(11) <= \R4_data[11]\;
    R4_data(10) <= \R4_data[10]\;
    R4_data(9) <= \R4_data[9]\;
    R4_data(8) <= \R4_data[8]\;
    R4_data(7) <= \R4_data[7]\;
    R4_data(6) <= \R4_data[6]\;
    R4_data(5) <= \R4_data[5]\;
    R4_data(4) <= \R4_data[4]\;
    R4_data(3) <= \R4_data[3]\;
    R4_data(2) <= \R4_data[2]\;
    R4_data(1) <= \R4_data[1]\;
    R4_data(0) <= \R4_data[0]\;

    sum3_6_0_cry_24 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[24]\, B => \R4_data[24]\, C => 
        \R5_data[24]\, D => \R6_data[24]\, FCI => 
        \sum3_6_0_cry_23\, S => \sum3_6_0[24]\, Y => OPEN, FCO
         => \sum3_6_0_cry_24\);
    
    \next_reg_h[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(11), B => \R6_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[11]_net_1\);
    
    sum3_cry_24 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[24]\, B => Wt_data(24), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_23\, S => 
        \sum3[24]\, Y => OPEN, FCO => \sum3_cry_24\);
    
    \reg_f[12]\ : SLE
      port map(D => \next_reg_f[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[12]\);
    
    sum3_cry_30 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[30]\, B => Wt_data(30), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_29\, S => 
        \sum3[30]\, Y => OPEN, FCO => \sum3_cry_30\);
    
    \next_reg_c[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(14), B => \R1_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[14]_net_1\);
    
    \reg_f[11]\ : SLE
      port map(D => \next_reg_f[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[11]\);
    
    sum3_6_0_cry_21 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[21]\, B => \R4_data[21]\, C => 
        \R5_data[21]\, D => \R6_data[21]\, FCI => 
        \sum3_6_0_cry_20\, S => \sum3_6_0[21]\, Y => OPEN, FCO
         => \sum3_6_0_cry_21\);
    
    \reg_h[22]\ : SLE
      port map(D => \next_reg_h[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[22]\);
    
    sum0_4_cry_0 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => sum0_4_0, C => \sum0_4[0]\, D
         => GND_net_1, FCI => GND_net_1, S => OPEN, Y => 
        sum0_4_cry_0_Y_0, FCO => \sum0_4_cry_0\);
    
    \reg_e[14]\ : SLE
      port map(D => \next_reg_e[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[14]\);
    
    \reg_h[21]\ : SLE
      port map(D => \next_reg_h[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[21]\);
    
    sum3_6_cry_11 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[11]\, B => \R4_data[4]\, C => 
        \R4_data[17]\, D => \R4_data[22]\, FCI => \sum3_6_cry_10\, 
        S => \sum3_6[11]\, Y => OPEN, FCO => \sum3_6_cry_11\);
    
    \SIG0[26]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[16]\, C => 
        \R0_data[7]\, Y => \SIG0[26]_net_1\);
    
    \next_reg_f[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(9), B => \R4_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[9]_net_1\);
    
    next_reg_a_cry_23_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[23]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[23]\, D => N0_data(23), FCI => next_reg_a_cry_22, S
         => \next_reg_a[23]\, Y => OPEN, FCO => next_reg_a_cry_23);
    
    \next_reg_g[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[0]\, B => next_reg_H6_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_g[0]_net_1\);
    
    sum3_cry_0_972 : CFG4
      generic map(INIT => x"A3A0")

      port map(A => next_r0_0_cry_0_Y, B => W_out_i_1(0), C => 
        ld_i_i_3, D => N_98, Y => \Wt_data_0[0]\);
    
    \next_reg_g[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(10), B => \R5_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[10]_net_1\);
    
    \next_reg_b[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(27), B => \R0_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[27]_net_1\);
    
    \next_reg_b[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(25), B => \R0_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[25]_net_1\);
    
    sum3_cry_26 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[26]\, B => Wt_data(26), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_25\, S => 
        \sum3[26]\, Y => OPEN, FCO => \sum3_cry_26\);
    
    \reg_d[17]\ : SLE
      port map(D => \next_reg_d[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[17]\);
    
    sum3_4_cry_5 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[5]\, B => m78, C => m83_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_4\, S => \sum3_4[5]\, Y
         => OPEN, FCO => \sum3_4_cry_5\);
    
    \reg_f[3]\ : SLE
      port map(D => \next_reg_f[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[3]\);
    
    \next_reg_f[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(27), B => \R4_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[27]_net_1\);
    
    sum0_4_cry_20 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[20]\, C => 
        \sum0_4_axb_20\, D => GND_net_1, FCI => \sum0_4_cry_19\, 
        S => \sum0_4[20]\, Y => OPEN, FCO => \sum0_4_cry_20\);
    
    sum3_6_cry_29 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[29]\, B => \R4_data[3]\, C => 
        \R4_data[8]\, D => \R4_data[22]\, FCI => \sum3_6_cry_28\, 
        S => \sum3_6[29]\, Y => OPEN, FCO => \sum3_6_cry_29\);
    
    \reg_g[13]\ : SLE
      port map(D => \next_reg_g[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[13]\);
    
    \next_reg_f[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(25), B => \R4_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[25]_net_1\);
    
    \reg_c[23]\ : SLE
      port map(D => \next_reg_c[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[23]\);
    
    sum0_4_cry_0_993 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[0]\, C => 
        \R0_data[12]\, Y => \SIG0_0[10]\);
    
    next_reg_e_cry_11_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[11]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(11), D => \R3_data[11]\, FCI => next_reg_e_cry_10, 
        S => \next_reg_e[11]\, Y => OPEN, FCO => 
        next_reg_e_cry_11);
    
    \reg_f[16]\ : SLE
      port map(D => \next_reg_f[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[16]\);
    
    \next_reg_d[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(13), B => \R2_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[13]_net_1\);
    
    \reg_b[29]\ : SLE
      port map(D => \next_reg_b[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[29]\);
    
    \reg_h[26]\ : SLE
      port map(D => \next_reg_h[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[26]\);
    
    sum3_6_cry_26 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[26]\, B => \R4_data[0]\, C => 
        \R4_data[5]\, D => \R4_data[19]\, FCI => \sum3_6_cry_25\, 
        S => \sum3_6[26]\, Y => OPEN, FCO => \sum3_6_cry_26\);
    
    \reg_a[15]\ : SLE
      port map(D => \next_reg_a[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[15]\);
    
    \reg_e[22]\ : SLE
      port map(D => \next_reg_e[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[22]\);
    
    \next_reg_h[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(20), B => \R6_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[20]_net_1\);
    
    \next_reg_g[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(12), B => \R5_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[12]_net_1\);
    
    \reg_e[21]\ : SLE
      port map(D => \next_reg_e[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[21]\);
    
    \next_reg_g[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(21), B => \R5_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[21]_net_1\);
    
    next_reg_a_cry_13_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[13]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[13]\, D => N0_data(13), FCI => next_reg_a_cry_12, S
         => \next_reg_a[13]\, Y => OPEN, FCO => next_reg_a_cry_13);
    
    \reg_d[8]\ : SLE
      port map(D => \next_reg_d[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[8]\);
    
    next_reg_e_cry_18_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[18]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(18), D => \R3_data[18]\, FCI => next_reg_e_cry_17, 
        S => \next_reg_e[18]\, Y => OPEN, FCO => 
        next_reg_e_cry_18);
    
    \next_reg_c[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(8), B => \R1_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[8]_net_1\);
    
    \reg_a[25]\ : SLE
      port map(D => \next_reg_a[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[25]\);
    
    \next_reg_g[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(31), B => \R5_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[31]_net_1\);
    
    \next_reg_c[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[2]\, B => N2_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[2]_net_1\);
    
    sum3_6_0_cry_2 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[2]\, B => \R4_data[2]\, C => 
        \R5_data[2]\, D => \R6_data[2]\, FCI => \sum3_6_0_cry_1\, 
        S => \sum3_6_0[2]\, Y => OPEN, FCO => \sum3_6_0_cry_2\);
    
    \next_reg_b[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(14), B => \R0_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[14]_net_1\);
    
    \next_reg_b[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(7), B => \R0_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[7]_net_1\);
    
    sum0_4_cry_23 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[23]\, C => 
        \sum0_4_axb_23\, D => GND_net_1, FCI => \sum0_4_cry_22\, 
        S => \sum0_4[23]\, Y => OPEN, FCO => \sum0_4_cry_23\);
    
    \reg_f[18]\ : SLE
      port map(D => \next_reg_f[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[18]\);
    
    \reg_b[4]\ : SLE
      port map(D => \next_reg_b[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[4]\);
    
    \next_reg_f[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(31), B => \R4_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[31]_net_1\);
    
    sum0_4_cry_0_1003 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[22]\, B => \R0_data[13]\, C => 
        \R0_data[2]\, Y => sum0_4_0);
    
    \SIG0[14]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[16]\, C => 
        \R0_data[4]\, Y => \SIG0[14]_net_1\);
    
    \reg_h[28]\ : SLE
      port map(D => \next_reg_h[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[28]\);
    
    \reg_b[7]\ : SLE
      port map(D => \next_reg_b[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[7]\);
    
    sum0_4_cry_17 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[17]\, C => 
        \sum0_4_axb_17\, D => GND_net_1, FCI => \sum0_4_cry_16\, 
        S => \sum0_4[17]\, Y => OPEN, FCO => \sum0_4_cry_17\);
    
    \reg_g[14]\ : SLE
      port map(D => \next_reg_g[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[14]\);
    
    \reg_c[24]\ : SLE
      port map(D => \next_reg_c[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[24]\);
    
    \next_reg_b[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(9), B => \R0_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[9]_net_1\);
    
    sum0_4_cry_0_996 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[20]\, C => 
        \R0_data[9]\, Y => \SIG0_0[7]\);
    
    \reg_h[15]\ : SLE
      port map(D => \next_reg_h[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[15]\);
    
    next_reg_e_cry_3_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[3]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(3), D => \R3_data[3]\, FCI => next_reg_e_cry_2, S
         => \next_reg_e[3]\, Y => OPEN, FCO => next_reg_e_cry_3);
    
    \next_reg_h[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(22), B => \R6_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[22]_net_1\);
    
    sum0_4_cry_28 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[28]\, C => 
        \sum0_4_axb_28\, D => GND_net_1, FCI => \sum0_4_cry_27\, 
        S => \sum0_4[28]\, Y => OPEN, FCO => \sum0_4_cry_28\);
    
    \reg_f[23]\ : SLE
      port map(D => \next_reg_f[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[23]\);
    
    \reg_e[26]\ : SLE
      port map(D => \next_reg_e[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[26]\);
    
    sum3_6_cry_8 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[8]\, B => \R4_data[1]\, C => 
        \R4_data[14]\, D => \R4_data[19]\, FCI => \sum3_6_cry_7\, 
        S => \sum3_6[8]\, Y => OPEN, FCO => \sum3_6_cry_8\);
    
    sum3_6_cry_22 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[22]\, B => \R4_data[1]\, C => 
        \R4_data[15]\, D => \R4_data[28]\, FCI => \sum3_6_cry_21\, 
        S => \sum3_6[22]\, Y => OPEN, FCO => \sum3_6_cry_22\);
    
    \reg_e[9]\ : SLE
      port map(D => \next_reg_e[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[9]\);
    
    \reg_g[9]\ : SLE
      port map(D => \next_reg_g[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[9]\);
    
    \reg_d[22]\ : SLE
      port map(D => \next_reg_d[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[22]\);
    
    \next_reg_d[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(7), B => \R2_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[7]_net_1\);
    
    \next_reg_c[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(7), B => \R1_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[7]_net_1\);
    
    \reg_d[21]\ : SLE
      port map(D => \next_reg_d[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[21]\);
    
    sum3_4_cry_11 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[11]\, B => m141, C => m144_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_10\, S => \sum3_4[11]\, Y
         => OPEN, FCO => \sum3_4_cry_11\);
    
    \next_reg_c[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(17), B => \R1_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[17]_net_1\);
    
    \next_reg_h[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(31), B => \R6_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[31]_net_1\);
    
    \next_reg_c[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(15), B => \R1_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[15]_net_1\);
    
    \next_reg_b[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(20), B => \R0_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[20]_net_1\);
    
    \reg_e[19]\ : SLE
      port map(D => \next_reg_e[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[19]\);
    
    sum3_cry_10 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[10]\, B => Wt_data(10), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_9\, S => 
        \sum3[10]\, Y => OPEN, FCO => \sum3_cry_10\);
    
    sum3_cry_2 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[2]\, B => Wt_data(2), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_1\, S => \sum3[2]\, Y
         => OPEN, FCO => \sum3_cry_2\);
    
    \next_reg_d[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(18), B => \R2_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[18]_net_1\);
    
    \reg_e[28]\ : SLE
      port map(D => \next_reg_e[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[28]\);
    
    sum3_cry_27 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[27]\, B => Wt_data(27), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_26\, S => 
        \sum3[27]\, Y => OPEN, FCO => \sum3_cry_27\);
    
    \reg_e[8]\ : SLE
      port map(D => \next_reg_e[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[8]\);
    
    sum0_4_cry_0_1002 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[14]\, C => 
        \R0_data[3]\, Y => \SIG0_0[1]\);
    
    \next_reg_d[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[0]\, B => next_reg_H3_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_d[0]_net_1\);
    
    \next_reg_f[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(20), B => \R4_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[20]_net_1\);
    
    \reg_b[27]\ : SLE
      port map(D => \next_reg_b[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[27]\);
    
    \next_reg_h[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(9), B => \R6_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[9]_net_1\);
    
    \next_reg_b[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[0]\, B => next_reg_H1_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_b[0]_net_1\);
    
    sum0_4_cry_0_980 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[13]\, C => 
        \R0_data[4]\, Y => \SIG0_0[23]\);
    
    \reg_b[13]\ : SLE
      port map(D => \next_reg_b[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[13]\);
    
    \reg_e[31]\ : SLE
      port map(D => \next_reg_e[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[31]\);
    
    sum3_6_0_cry_30 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[30]\, B => \R4_data[30]\, C => 
        \R5_data[30]\, D => \R6_data[30]\, FCI => 
        \sum3_6_0_cry_29\, S => \sum3_6_0[30]\, Y => OPEN, FCO
         => \sum3_6_0_cry_30\);
    
    sum3_6_0_cry_13 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[13]\, B => \R4_data[13]\, C => 
        \R5_data[13]\, D => \R6_data[13]\, FCI => 
        \sum3_6_0_cry_12\, S => \sum3_6_0[13]\, Y => OPEN, FCO
         => \sum3_6_0_cry_13\);
    
    \reg_f[24]\ : SLE
      port map(D => \next_reg_f[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[24]\);
    
    \next_reg_d[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(29), B => \R2_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[29]_net_1\);
    
    \next_reg_f[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(11), B => \R4_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[11]_net_1\);
    
    \SIG0[15]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[17]\, C => 
        \R0_data[5]\, Y => \SIG0[15]_net_1\);
    
    \reg_a[10]\ : SLE
      port map(D => \next_reg_a[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[10]\);
    
    \next_reg_f[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[6]\, B => N5_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[6]_net_1\);
    
    \reg_d[9]\ : SLE
      port map(D => \next_reg_d[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[9]\);
    
    \reg_d[26]\ : SLE
      port map(D => \next_reg_d[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[26]\);
    
    \reg_a[20]\ : SLE
      port map(D => \next_reg_a[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[20]\);
    
    \next_reg_b[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(22), B => \R0_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[22]_net_1\);
    
    \next_reg_c[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(24), B => \R1_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[24]_net_1\);
    
    \reg_f[1]\ : SLE
      port map(D => \next_reg_f[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[1]\);
    
    sum3_6_0_cry_25 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[25]\, B => \R4_data[25]\, C => 
        \R5_data[25]\, D => \R6_data[25]\, FCI => 
        \sum3_6_0_cry_24\, S => \sum3_6_0[25]\, Y => OPEN, FCO
         => \sum3_6_0_cry_25\);
    
    sum3_4_cry_4 : ARI1
      generic map(INIT => x"5C53A")

      port map(A => \sum3_6[4]\, B => m67_ns, C => m73, D => 
        Kt_addr(5), FCI => \sum3_4_cry_3\, S => \sum3_4[4]\, Y
         => OPEN, FCO => \sum3_4_cry_4\);
    
    \next_reg_f[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(22), B => \R4_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[22]_net_1\);
    
    sum0_4_axb_28 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[28]\, B => \R1_data[28]\, C => 
        \R0_data[28]\, D => \SIG0[28]_net_1\, Y => 
        \sum0_4_axb_28\);
    
    sum0_4_cry_14 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[14]\, C => 
        \sum0_4_axb_14\, D => GND_net_1, FCI => \sum0_4_cry_13\, 
        S => \sum0_4[14]\, Y => OPEN, FCO => \sum0_4_cry_14\);
    
    sum3_6_cry_30 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[30]\, B => \R4_data[4]\, C => 
        \R4_data[9]\, D => \R4_data[23]\, FCI => \sum3_6_cry_29\, 
        S => \sum3_6[30]\, Y => OPEN, FCO => \sum3_6_cry_30\);
    
    \next_reg_b[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(17), B => \R0_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[17]_net_1\);
    
    \reg_a[0]\ : SLE
      port map(D => next_reg_a_cry_0_0_Y, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[0]\);
    
    \reg_h[10]\ : SLE
      port map(D => \next_reg_h[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[10]\);
    
    \reg_b[14]\ : SLE
      port map(D => \next_reg_b[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[14]\);
    
    \next_reg_b[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(15), B => \R0_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[15]_net_1\);
    
    sum3_6_cry_10 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[10]\, B => \R4_data[3]\, C => 
        \R4_data[16]\, D => \R4_data[21]\, FCI => \sum3_6_cry_9\, 
        S => \sum3_6[10]\, Y => OPEN, FCO => \sum3_6_cry_10\);
    
    \reg_d[28]\ : SLE
      port map(D => \next_reg_d[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[28]\);
    
    \reg_d[2]\ : SLE
      port map(D => \next_reg_d[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[2]\);
    
    next_reg_e_cry_26_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[26]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(26), D => \R3_data[26]\, FCI => next_reg_e_cry_25, 
        S => \next_reg_e[26]\, Y => OPEN, FCO => 
        next_reg_e_cry_26);
    
    \reg_f[4]\ : SLE
      port map(D => \next_reg_f[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[4]\);
    
    \next_reg_c[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[5]\, B => N2_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[5]_net_1\);
    
    \reg_f[9]\ : SLE
      port map(D => \next_reg_f[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[9]\);
    
    sum3_4_cry_27 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[27]\, B => m289, C => m292_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_26\, S => \sum3_4[27]\, Y
         => OPEN, FCO => \sum3_4_cry_27\);
    
    sum3_6_0_cry_6 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[6]\, B => \R4_data[6]\, C => 
        \R5_data[6]\, D => \R6_data[6]\, FCI => \sum3_6_0_cry_5\, 
        S => \sum3_6_0[6]\, Y => OPEN, FCO => \sum3_6_0_cry_6\);
    
    \reg_g[19]\ : SLE
      port map(D => \next_reg_g[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[19]\);
    
    \next_reg_d[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(16), B => \R2_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[16]_net_1\);
    
    \next_reg_c[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[4]\, B => N2_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[4]_net_1\);
    
    \reg_c[29]\ : SLE
      port map(D => \next_reg_c[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[29]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \next_reg_g[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(8), B => \R5_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[8]_net_1\);
    
    sum0_4_cry_29 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[29]\, C => 
        \sum0_4_axb_29\, D => GND_net_1, FCI => \sum0_4_cry_28\, 
        S => \sum0_4[29]\, Y => OPEN, FCO => \sum0_4_cry_29\);
    
    \next_reg_g[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(11), B => \R5_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[11]_net_1\);
    
    \reg_e[17]\ : SLE
      port map(D => \next_reg_e[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[17]\);
    
    \reg_g[1]\ : SLE
      port map(D => \next_reg_g[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[1]\);
    
    \next_reg_b[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[3]\, B => N1_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[3]_net_1\);
    
    sum3_cry_19 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[19]\, B => Wt_data(19), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_18\, S => 
        \sum3[19]\, Y => OPEN, FCO => \sum3_cry_19\);
    
    sum0_4_cry_26 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[26]\, C => 
        \sum0_4_axb_26\, D => GND_net_1, FCI => \sum0_4_cry_25\, 
        S => \sum0_4[26]\, Y => OPEN, FCO => \sum0_4_cry_26\);
    
    \next_reg_c[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(10), B => \R1_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[10]_net_1\);
    
    sum3_cry_18 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[18]\, B => Wt_data(18), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_17\, S => 
        \sum3[18]\, Y => OPEN, FCO => \sum3_cry_18\);
    
    \reg_a[31]\ : SLE
      port map(D => \next_reg_a[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[31]\);
    
    \next_reg_h[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(13), B => \R6_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[13]_net_1\);
    
    sum3_6_cry_13 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[13]\, B => \R4_data[6]\, C => 
        \R4_data[19]\, D => \R4_data[24]\, FCI => \sum3_6_cry_12\, 
        S => \sum3_6[13]\, Y => OPEN, FCO => \sum3_6_cry_13\);
    
    sum0_4_axb_6 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[6]\, B => \R1_data[6]\, C => 
        \R0_data[6]\, D => \SIG0[6]_net_1\, Y => \sum0_4_axb_6\);
    
    \reg_g[25]\ : SLE
      port map(D => \next_reg_g[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[25]\);
    
    sum0_4_cry_0_979 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[14]\, C => 
        \R0_data[5]\, Y => \SIG0_0[24]\);
    
    \next_reg_h[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(21), B => \R6_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[21]_net_1\);
    
    sum3_6_cry_18 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[18]\, B => \R4_data[11]\, C => 
        \R4_data[24]\, D => \R4_data[29]\, FCI => \sum3_6_cry_17\, 
        S => \sum3_6[18]\, Y => OPEN, FCO => \sum3_6_cry_18\);
    
    \reg_h[0]\ : SLE
      port map(D => \next_reg_h[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[0]\);
    
    sum3_4_cry_6 : ARI1
      generic map(INIT => x"53AC5")

      port map(A => \sum3_6[6]\, B => m95_1_0, C => m95_1_1, D
         => Kt_addr(5), FCI => \sum3_4_cry_5\, S => \sum3_4[6]\, 
        Y => OPEN, FCO => \sum3_4_cry_6\);
    
    \reg_c[31]\ : SLE
      port map(D => \next_reg_c[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[31]\);
    
    \next_reg_c[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(12), B => \R1_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[12]_net_1\);
    
    \reg_f[29]\ : SLE
      port map(D => \next_reg_f[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[29]\);
    
    next_reg_e_cry_21_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[21]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(21), D => \R3_data[21]\, FCI => next_reg_e_cry_20, 
        S => \next_reg_e[21]\, Y => OPEN, FCO => 
        next_reg_e_cry_21);
    
    sum3_6_cry_4 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[4]\, B => \R4_data[10]\, C => 
        \R4_data[15]\, D => \R4_data[29]\, FCI => \sum3_6_cry_3\, 
        S => \sum3_6[4]\, Y => OPEN, FCO => \sum3_6_cry_4\);
    
    sum0_4_cry_22 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[22]\, C => 
        \sum0_4_axb_22\, D => GND_net_1, FCI => \sum0_4_cry_21\, 
        S => \sum0_4[22]\, Y => OPEN, FCO => \sum0_4_cry_22\);
    
    \next_reg_c[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(27), B => \R1_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[27]_net_1\);
    
    sum3_cry_7 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[7]\, B => Wt_data(7), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_6\, S => \sum3[7]\, Y
         => OPEN, FCO => \sum3_cry_7\);
    
    \reg_g[6]\ : SLE
      port map(D => \next_reg_g[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[6]\);
    
    \next_reg_c[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(25), B => \R1_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[25]_net_1\);
    
    next_reg_e_cry_28_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[28]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(28), D => \R3_data[28]\, FCI => next_reg_e_cry_27, 
        S => \next_reg_e[28]\, Y => OPEN, FCO => 
        next_reg_e_cry_28);
    
    \next_reg_g[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(23), B => \R5_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[23]_net_1\);
    
    \next_reg_b[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(10), B => \R0_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[10]_net_1\);
    
    \SIG0[12]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[14]\, C => 
        \R0_data[2]\, Y => \SIG0[12]_net_1\);
    
    \reg_g[17]\ : SLE
      port map(D => \next_reg_g[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[17]\);
    
    \reg_c[27]\ : SLE
      port map(D => \next_reg_c[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[27]\);
    
    sum3_4_cry_24 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_6[24]\, B => Kt_data_9, C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_4_cry_23\, S => \sum3_4[24]\, 
        Y => OPEN, FCO => \sum3_4_cry_24\);
    
    \reg_d[0]\ : SLE
      port map(D => \next_reg_d[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[0]\);
    
    sum3_4_cry_10 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[10]\, B => m137_am, C => m137_bm, D
         => Kt_addr(5), FCI => \sum3_4_cry_9\, S => \sum3_4[10]\, 
        Y => OPEN, FCO => \sum3_4_cry_10\);
    
    \next_reg_d[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[2]\, B => N3_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[2]_net_1\);
    
    \reg_a[13]\ : SLE
      port map(D => \next_reg_a[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[13]\);
    
    \reg_h[4]\ : SLE
      port map(D => \next_reg_h[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[4]\);
    
    \reg_b[19]\ : SLE
      port map(D => \next_reg_b[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[19]\);
    
    \next_reg_h[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[6]\, B => N7_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[6]_net_1\);
    
    \next_reg_h[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(18), B => \R6_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[18]_net_1\);
    
    \reg_a[23]\ : SLE
      port map(D => \next_reg_a[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[23]\);
    
    sum3_cry_15 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[15]\, B => Wt_data(15), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_14\, S => 
        \sum3[15]\, Y => OPEN, FCO => \sum3_cry_15\);
    
    \next_reg_b[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(21), B => \R0_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[21]_net_1\);
    
    sum3_6_0_cry_28 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[28]\, B => \R4_data[28]\, C => 
        \R5_data[28]\, D => \R6_data[28]\, FCI => 
        \sum3_6_0_cry_27\, S => \sum3_6_0[28]\, Y => OPEN, FCO
         => \sum3_6_0_cry_28\);
    
    \reg_b[5]\ : SLE
      port map(D => \next_reg_b[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[5]\);
    
    \reg_b[3]\ : SLE
      port map(D => \next_reg_b[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[3]\);
    
    next_reg_a_cry_26_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[26]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[26]\, D => N0_data(26), FCI => next_reg_a_cry_25, S
         => \next_reg_a[26]\, Y => OPEN, FCO => next_reg_a_cry_26);
    
    sum3_6_cry_5 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[5]\, B => \R4_data[11]\, C => 
        \R4_data[16]\, D => \R4_data[30]\, FCI => \sum3_6_cry_4\, 
        S => \sum3_6[5]\, Y => OPEN, FCO => \sum3_6_cry_5\);
    
    \SIG0[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[22]\, B => \R0_data[13]\, C => 
        \R0_data[2]\, Y => sum0_4);
    
    \next_reg_b[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(12), B => \R0_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[12]_net_1\);
    
    \next_reg_f[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(21), B => \R4_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[21]_net_1\);
    
    sum3_6_cry_27 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[27]\, B => \R4_data[1]\, C => 
        \R4_data[6]\, D => \R4_data[20]\, FCI => \sum3_6_cry_26\, 
        S => \sum3_6[27]\, Y => OPEN, FCO => \sum3_6_cry_27\);
    
    \next_reg_d[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(24), B => \R2_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[24]_net_1\);
    
    sum3_4_cry_13 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[13]\, B => m168_1_0, C => m168_1_1, D
         => Kt_addr(5), FCI => \sum3_4_cry_12\, S => \sum3_4[13]\, 
        Y => OPEN, FCO => \sum3_4_cry_13\);
    
    sum3_6_0_cry_10 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[10]\, B => \R4_data[10]\, C => 
        \R5_data[10]\, D => \R6_data[10]\, FCI => 
        \sum3_6_0_cry_9\, S => \sum3_6_0[10]\, Y => OPEN, FCO => 
        \sum3_6_0_cry_10\);
    
    \reg_h[13]\ : SLE
      port map(D => \next_reg_h[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[13]\);
    
    \reg_g[20]\ : SLE
      port map(D => \next_reg_g[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[20]\);
    
    sum3_6_0_cry_16 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[16]\, B => \R4_data[16]\, C => 
        \R5_data[16]\, D => \R6_data[16]\, FCI => 
        \sum3_6_0_cry_15\, S => \sum3_6_0[16]\, Y => OPEN, FCO
         => \sum3_6_0_cry_16\);
    
    \SIG0[30]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[20]\, B => \R0_data[11]\, C => 
        \R0_data[0]\, Y => \SIG0[30]_net_1\);
    
    sum3_6_0_cry_3 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[3]\, B => \R4_data[3]\, C => 
        \R5_data[3]\, D => \R6_data[3]\, FCI => \sum3_6_0_cry_2\, 
        S => \sum3_6_0[3]\, Y => OPEN, FCO => \sum3_6_0_cry_3\);
    
    \reg_a[14]\ : SLE
      port map(D => \next_reg_a[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[14]\);
    
    \reg_e[5]\ : SLE
      port map(D => \next_reg_e[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[5]\);
    
    \reg_f[27]\ : SLE
      port map(D => \next_reg_f[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[27]\);
    
    \reg_c[12]\ : SLE
      port map(D => \next_reg_c[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[12]\);
    
    \reg_f[15]\ : SLE
      port map(D => \next_reg_f[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[15]\);
    
    \reg_c[11]\ : SLE
      port map(D => \next_reg_c[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[11]\);
    
    sum3_4_cry_18 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[18]\, B => m215_am, C => m215_bm, D
         => Kt_addr(5), FCI => \sum3_4_cry_17\, S => \sum3_4[18]\, 
        Y => OPEN, FCO => \sum3_4_cry_18\);
    
    \SIG0[16]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[18]\, C => 
        \R0_data[6]\, Y => \SIG0[16]_net_1\);
    
    \reg_h[25]\ : SLE
      port map(D => \next_reg_h[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[25]\);
    
    sum3_6_cry_19 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[19]\, B => \R4_data[12]\, C => 
        \R4_data[25]\, D => \R4_data[30]\, FCI => \sum3_6_cry_18\, 
        S => \sum3_6[19]\, Y => OPEN, FCO => \sum3_6_cry_19\);
    
    \reg_b[2]\ : SLE
      port map(D => \next_reg_b[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[2]\);
    
    \reg_a[24]\ : SLE
      port map(D => \next_reg_a[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[24]\);
    
    sum3_cry_22 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[22]\, B => Wt_data(22), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_21\, S => 
        \sum3[22]\, Y => OPEN, FCO => \sum3_cry_22\);
    
    next_reg_e_cry_12_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[12]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(12), D => \R3_data[12]\, FCI => next_reg_e_cry_11, 
        S => \next_reg_e[12]\, Y => OPEN, FCO => 
        next_reg_e_cry_12);
    
    \next_reg_f[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[0]\, B => next_reg_H5_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_f[0]_net_1\);
    
    next_reg_a_cry_16_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[16]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[16]\, D => N0_data(16), FCI => next_reg_a_cry_15, S
         => \next_reg_a[16]\, Y => OPEN, FCO => next_reg_a_cry_16);
    
    \next_reg_g[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(28), B => \R5_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[28]_net_1\);
    
    sum3_6_cry_16 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[16]\, B => \R4_data[9]\, C => 
        \R4_data[22]\, D => \R4_data[27]\, FCI => \sum3_6_cry_15\, 
        S => \sum3_6[16]\, Y => OPEN, FCO => \sum3_6_cry_16\);
    
    \next_reg_d[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[1]\, B => N3_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[1]_net_1\);
    
    \next_reg_f[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(13), B => \R4_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[13]_net_1\);
    
    next_reg_e_cry_4_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[4]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(4), D => \R3_data[4]\, FCI => next_reg_e_cry_3, S
         => \next_reg_e[4]\, Y => OPEN, FCO => next_reg_e_cry_4);
    
    \reg_f[2]\ : SLE
      port map(D => \next_reg_f[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[2]\);
    
    \next_reg_h[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(16), B => \R6_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[16]_net_1\);
    
    sum0_4_cry_1 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[1]\, C => 
        \sum0_4_axb_1\, D => GND_net_1, FCI => \sum0_4_cry_0\, S
         => \sum0_4[1]\, Y => OPEN, FCO => \sum0_4_cry_1\);
    
    \next_reg_c[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(20), B => \R1_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[20]_net_1\);
    
    sum0_4_cry_15 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[15]\, C => 
        \sum0_4_axb_15\, D => GND_net_1, FCI => \sum0_4_cry_14\, 
        S => \sum0_4[15]\, Y => OPEN, FCO => \sum0_4_cry_15\);
    
    \next_reg_b[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[5]\, B => N1_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[5]_net_1\);
    
    \reg_h[14]\ : SLE
      port map(D => \next_reg_h[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[14]\);
    
    next_reg_e_cry_9_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[9]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(9), D => \R3_data[9]\, FCI => next_reg_e_cry_8, S
         => \next_reg_e[9]\, Y => OPEN, FCO => next_reg_e_cry_9);
    
    \reg_b[17]\ : SLE
      port map(D => \next_reg_b[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[17]\);
    
    \SIG0[29]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[19]\, C => 
        \R0_data[10]\, Y => \SIG0[29]_net_1\);
    
    next_reg_a_cry_21_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[21]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[21]\, D => N0_data(21), FCI => next_reg_a_cry_20, S
         => \next_reg_a[21]\, Y => OPEN, FCO => next_reg_a_cry_21);
    
    \reg_c[16]\ : SLE
      port map(D => \next_reg_c[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[16]\);
    
    sum0_4_cry_7 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[7]\, C => 
        \sum0_4_axb_7\, D => GND_net_1, FCI => \sum0_4_cry_6\, S
         => \sum0_4[7]\, Y => OPEN, FCO => \sum0_4_cry_7\);
    
    \reg_h[8]\ : SLE
      port map(D => \next_reg_h[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[8]\);
    
    next_reg_a_cry_4_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[4]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[4]\, D => N0_data(4), FCI => next_reg_a_cry_3, S
         => \next_reg_a[4]\, Y => OPEN, FCO => next_reg_a_cry_4);
    
    \reg_e[25]\ : SLE
      port map(D => \next_reg_e[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[25]\);
    
    \reg_a[8]\ : SLE
      port map(D => \next_reg_a[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[8]\);
    
    sum3_cry_14 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[14]\, B => Wt_data(14), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_13\, S => 
        \sum3[14]\, Y => OPEN, FCO => \sum3_cry_14\);
    
    \next_reg_c[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(11), B => \R1_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[11]_net_1\);
    
    sum3_cry_3 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[3]\, B => Wt_data(3), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_2\, S => \sum3[3]\, Y
         => OPEN, FCO => \sum3_cry_3\);
    
    next_reg_a_cry_28_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[28]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[28]\, D => N0_data(28), FCI => next_reg_a_cry_27, S
         => \next_reg_a[28]\, Y => OPEN, FCO => next_reg_a_cry_28);
    
    \next_reg_c[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(22), B => \R1_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[22]_net_1\);
    
    sum0_4_axb_18 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[18]\, B => \R1_data[18]\, C => 
        \R0_data[18]\, D => \SIG0[18]_net_1\, Y => 
        \sum0_4_axb_18\);
    
    \next_reg_h[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(8), B => \R6_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[8]_net_1\);
    
    sum0_4_cry_0_989 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[16]\, C => 
        \R0_data[4]\, Y => \SIG0_0[14]\);
    
    \reg_f[30]\ : SLE
      port map(D => \next_reg_f[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[30]\);
    
    sum3_6_cry_24 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[24]\, B => \R4_data[3]\, C => 
        \R4_data[17]\, D => \R4_data[30]\, FCI => \sum3_6_cry_23\, 
        S => \sum3_6[24]\, Y => OPEN, FCO => \sum3_6_cry_24\);
    
    sum3_6_cry_12 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[12]\, B => \R4_data[5]\, C => 
        \R4_data[18]\, D => \R4_data[23]\, FCI => \sum3_6_cry_11\, 
        S => \sum3_6[12]\, Y => OPEN, FCO => \sum3_6_cry_12\);
    
    \reg_c[18]\ : SLE
      port map(D => \next_reg_c[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[18]\);
    
    next_reg_e_cry_5_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[5]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(5), D => \R3_data[5]\, FCI => next_reg_e_cry_4, S
         => \next_reg_e[5]\, Y => OPEN, FCO => next_reg_e_cry_5);
    
    sum3_6_0_s_31 : ARI1
      generic map(INIT => x"427D8")

      port map(A => \R7_data[31]\, B => \R4_data[31]\, C => 
        \R5_data[31]\, D => \R6_data[31]\, FCI => 
        \sum3_6_0_cry_30\, S => \sum3_6_0[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_e_cry_8_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[8]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(8), D => \R3_data[8]\, FCI => next_reg_e_cry_7, S
         => \next_reg_e[8]\, Y => OPEN, FCO => next_reg_e_cry_8);
    
    \next_reg_g[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[1]\, B => N6_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[1]_net_1\);
    
    \next_reg_g[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(13), B => \R5_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[13]_net_1\);
    
    \next_reg_g[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(26), B => \R5_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[26]_net_1\);
    
    \reg_b[6]\ : SLE
      port map(D => \next_reg_b[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[6]\);
    
    sum3_cry_16 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[16]\, B => Wt_data(16), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_15\, S => 
        \sum3[16]\, Y => OPEN, FCO => \sum3_cry_16\);
    
    \next_reg_d[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(27), B => \R2_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[27]_net_1\);
    
    sum3_6_cry_6 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[6]\, B => \R4_data[12]\, C => 
        \R4_data[17]\, D => \R4_data[31]\, FCI => \sum3_6_cry_5\, 
        S => \sum3_6[6]\, Y => OPEN, FCO => \sum3_6_cry_6\);
    
    next_reg_a_cry_11_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[11]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[11]\, D => N0_data(11), FCI => next_reg_a_cry_10, S
         => \next_reg_a[11]\, Y => OPEN, FCO => next_reg_a_cry_11);
    
    sum0_4_cry_0_975 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[18]\, C => 
        \R0_data[9]\, Y => \SIG0_0[28]\);
    
    sum0_4_s_31 : ARI1
      generic map(INIT => x"46996")

      port map(A => \R0_data[21]\, B => \Maj[31]_net_1\, C => 
        \R0_data[1]\, D => \R0_data[12]\, FCI => \sum0_4_cry_30\, 
        S => \sum0_4[31]\, Y => OPEN, FCO => OPEN);
    
    \next_reg_d[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(25), B => \R2_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[25]_net_1\);
    
    \reg_f[10]\ : SLE
      port map(D => \next_reg_f[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[10]\);
    
    sum0_4_cry_0_990 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[15]\, C => 
        \R0_data[3]\, Y => \SIG0_0[13]\);
    
    \reg_h[20]\ : SLE
      port map(D => \next_reg_h[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[20]\);
    
    \reg_d[12]\ : SLE
      port map(D => \next_reg_d[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[12]\);
    
    \next_reg_h[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[5]\, B => N7_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[5]_net_1\);
    
    sum0_4_cry_6 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[6]\, C => 
        \sum0_4_axb_6\, D => GND_net_1, FCI => \sum0_4_cry_5\, S
         => \sum0_4[6]\, Y => OPEN, FCO => \sum0_4_cry_6\);
    
    \reg_d[11]\ : SLE
      port map(D => \next_reg_d[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[11]\);
    
    \reg_c[2]\ : SLE
      port map(D => \next_reg_c[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[2]\);
    
    \next_reg_f[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(18), B => \R4_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[18]_net_1\);
    
    next_reg_a_cry_7_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[7]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[7]\, D => N0_data(7), FCI => next_reg_a_cry_6, S
         => \next_reg_a[7]\, Y => OPEN, FCO => next_reg_a_cry_7);
    
    \reg_d[25]\ : SLE
      port map(D => \next_reg_d[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[25]\);
    
    sum3_6_0_cry_22 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[22]\, B => \R4_data[22]\, C => 
        \R5_data[22]\, D => \R6_data[22]\, FCI => 
        \sum3_6_0_cry_21\, S => \sum3_6_0[22]\, Y => OPEN, FCO
         => \sum3_6_0_cry_22\);
    
    \reg_a[19]\ : SLE
      port map(D => \next_reg_a[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[19]\);
    
    sum3_4_cry_19 : ARI1
      generic map(INIT => x"53AC5")

      port map(A => \sum3_6[19]\, B => m219, C => m222_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_18\, S => \sum3_4[19]\, Y
         => OPEN, FCO => \sum3_4_cry_19\);
    
    next_reg_a_cry_18_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[18]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[18]\, D => N0_data(18), FCI => next_reg_a_cry_17, S
         => \next_reg_a[18]\, Y => OPEN, FCO => next_reg_a_cry_18);
    
    next_reg_e_cry_15_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[15]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(15), D => \R3_data[15]\, FCI => next_reg_e_cry_14, 
        S => \next_reg_e[15]\, Y => OPEN, FCO => 
        next_reg_e_cry_15);
    
    sum3_6_0_cry_14 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[14]\, B => \R4_data[14]\, C => 
        \R5_data[14]\, D => \R6_data[14]\, FCI => 
        \sum3_6_0_cry_13\, S => \sum3_6_0[14]\, Y => OPEN, FCO
         => \sum3_6_0_cry_14\);
    
    \next_reg_h[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(23), B => \R6_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[23]_net_1\);
    
    \reg_f[7]\ : SLE
      port map(D => \next_reg_f[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[7]\);
    
    \reg_a[29]\ : SLE
      port map(D => \next_reg_a[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[29]\);
    
    \next_reg_b[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(11), B => \R0_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[11]_net_1\);
    
    \reg_e[0]\ : SLE
      port map(D => next_reg_e_cry_0_0_Y, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[0]\);
    
    \SIG0[7]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[20]\, C => 
        \R0_data[9]\, Y => \SIG0[7]_net_1\);
    
    sum3_4_cry_16 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[16]\, B => m197_1_0, C => m197_1_1, D
         => Kt_addr(5), FCI => \sum3_4_cry_15\, S => \sum3_4[16]\, 
        Y => OPEN, FCO => \sum3_4_cry_16\);
    
    sum3_6_0_cry_11 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[11]\, B => \R4_data[11]\, C => 
        \R5_data[11]\, D => \R6_data[11]\, FCI => 
        \sum3_6_0_cry_10\, S => \sum3_6_0[11]\, Y => OPEN, FCO
         => \sum3_6_0_cry_11\);
    
    \next_reg_g[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[6]\, B => N6_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[6]_net_1\);
    
    sum0_4_cry_0_977 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[16]\, C => 
        \R0_data[7]\, Y => \SIG0_0[26]\);
    
    \reg_e[1]\ : SLE
      port map(D => \next_reg_e[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[1]\);
    
    \SIG0[23]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[13]\, C => 
        \R0_data[4]\, Y => \SIG0[23]_net_1\);
    
    \reg_g[23]\ : SLE
      port map(D => \next_reg_g[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[23]\);
    
    sum3_6_0_cry_5 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[5]\, B => \R4_data[5]\, C => 
        \R5_data[5]\, D => \R6_data[5]\, FCI => \sum3_6_0_cry_4\, 
        S => \sum3_6_0[5]\, Y => OPEN, FCO => \sum3_6_0_cry_5\);
    
    sum3_4_cry_2 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[2]\, B => m49_am, C => m49_bm, D => 
        Kt_addr(5), FCI => \sum3_4_cry_1\, S => \sum3_4[2]\, Y
         => OPEN, FCO => \sum3_4_cry_2\);
    
    sum3_4_cry_25 : ARI1
      generic map(INIT => x"5C53A")

      port map(A => \sum3_6[25]\, B => m273, C => m276_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_24\, S => \sum3_4[25]\, Y
         => OPEN, FCO => \sum3_4_cry_25\);
    
    \next_reg_d[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(19), B => \R2_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[19]_net_1\);
    
    \reg_d[16]\ : SLE
      port map(D => \next_reg_d[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[16]\);
    
    sum0_4_cry_27 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[27]\, C => 
        \sum0_4_axb_27\, D => GND_net_1, FCI => \sum0_4_cry_26\, 
        S => \sum0_4[27]\, Y => OPEN, FCO => \sum0_4_cry_27\);
    
    sum3_4_cry_30 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \sum3_6[30]\, B => m316, C => GND_net_1, D
         => GND_net_1, FCI => \sum3_4_cry_29\, S => \sum3_4[30]\, 
        Y => OPEN, FCO => \sum3_4_cry_30\);
    
    \reg_h[19]\ : SLE
      port map(D => \next_reg_h[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[19]\);
    
    \reg_e[20]\ : SLE
      port map(D => \next_reg_e[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[20]\);
    
    \reg_c[4]\ : SLE
      port map(D => \next_reg_c[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[4]\);
    
    sum0_4_axb_26 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[26]\, B => \R1_data[26]\, C => 
        \R0_data[26]\, D => \SIG0[26]_net_1\, Y => 
        \sum0_4_axb_26\);
    
    \reg_a[2]\ : SLE
      port map(D => \next_reg_a[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[2]\);
    
    sum0_4_cry_4 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[4]\, C => 
        \sum0_4_axb_4\, D => GND_net_1, FCI => \sum0_4_cry_3\, S
         => \sum0_4[4]\, Y => OPEN, FCO => \sum0_4_cry_4\);
    
    \next_reg_b[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[1]\, B => N1_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[1]_net_1\);
    
    sum3_cry_4 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[4]\, B => Wt_data(4), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_3\, S => \sum3[4]\, Y
         => OPEN, FCO => \sum3_cry_4\);
    
    sum0_4_axb_29 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[29]\, B => \R1_data[29]\, C => 
        \R0_data[29]\, D => \SIG0[29]_net_1\, Y => 
        \sum0_4_axb_29\);
    
    next_reg_e_cry_17_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[17]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(17), D => \R3_data[17]\, FCI => next_reg_e_cry_16, 
        S => \next_reg_e[17]\, Y => OPEN, FCO => 
        next_reg_e_cry_17);
    
    \next_reg_g[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(18), B => \R5_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[18]_net_1\);
    
    \next_reg_b[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(30), B => \R0_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[30]_net_1\);
    
    sum3_6_0_cry_27 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[27]\, B => \R4_data[27]\, C => 
        \R5_data[27]\, D => \R6_data[27]\, FCI => 
        \sum3_6_0_cry_26\, S => \sum3_6_0[27]\, Y => OPEN, FCO
         => \sum3_6_0_cry_27\);
    
    sum0_4_cry_8 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[8]\, C => 
        \sum0_4_axb_8\, D => GND_net_1, FCI => \sum0_4_cry_7\, S
         => \sum0_4[8]\, Y => OPEN, FCO => \sum0_4_cry_8\);
    
    \SIG0[4]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[17]\, C => 
        \R0_data[6]\, Y => \SIG0[4]_net_1\);
    
    \reg_d[18]\ : SLE
      port map(D => \next_reg_d[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[18]\);
    
    \next_reg_f[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(16), B => \R4_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[16]_net_1\);
    
    sum0_4_cry_3 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[3]\, C => 
        \sum0_4_axb_3\, D => GND_net_1, FCI => \sum0_4_cry_2\, S
         => \sum0_4[3]\, Y => OPEN, FCO => \sum0_4_cry_3\);
    
    \reg_g[5]\ : SLE
      port map(D => \next_reg_g[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[5]\);
    
    sum3_4_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \sum3_6[12]\, B => m157, C => GND_net_1, D
         => GND_net_1, FCI => \sum3_4_cry_11\, S => \sum3_4[12]\, 
        Y => OPEN, FCO => \sum3_4_cry_12\);
    
    \reg_g[24]\ : SLE
      port map(D => \next_reg_g[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[24]\);
    
    next_reg_a_cry_5_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[5]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[5]\, D => N0_data(5), FCI => next_reg_a_cry_4, S
         => \next_reg_a[5]\, Y => OPEN, FCO => next_reg_a_cry_5);
    
    sum3_cry_1 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[1]\, B => Wt_data(1), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_0\, S => \sum3[1]\, Y
         => OPEN, FCO => \sum3_cry_1\);
    
    \next_reg_b[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(23), B => \R0_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[23]_net_1\);
    
    sum3_6_0_cry_1 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[1]\, B => \R4_data[1]\, C => 
        \R5_data[1]\, D => \R6_data[1]\, FCI => \sum3_6_0_cry_0\, 
        S => \sum3_6_0[1]\, Y => OPEN, FCO => \sum3_6_0_cry_1\);
    
    sum3_cry_17 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[17]\, B => Wt_data(17), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_16\, S => 
        \sum3[17]\, Y => OPEN, FCO => \sum3_cry_17\);
    
    \SIG0[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[14]\, C => 
        \R0_data[3]\, Y => \SIG0[1]_net_1\);
    
    \next_reg_d[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(20), B => \R2_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[20]_net_1\);
    
    sum0_4_axb_21 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[21]\, B => \R1_data[21]\, C => 
        \R0_data[21]\, D => \SIG0[21]_net_1\, Y => 
        \sum0_4_axb_21\);
    
    \reg_a[17]\ : SLE
      port map(D => \next_reg_a[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[17]\);
    
    \SIG0[6]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[19]\, C => 
        \R0_data[8]\, Y => \SIG0[6]_net_1\);
    
    \next_reg_f[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(23), B => \R4_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[23]_net_1\);
    
    \reg_b[22]\ : SLE
      port map(D => \next_reg_b[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[22]\);
    
    \next_reg_h[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(28), B => \R6_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[28]_net_1\);
    
    \reg_d[20]\ : SLE
      port map(D => \next_reg_d[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[20]\);
    
    \reg_b[21]\ : SLE
      port map(D => \next_reg_b[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[21]\);
    
    \reg_f[0]\ : SLE
      port map(D => \next_reg_f[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[0]\);
    
    \reg_c[9]\ : SLE
      port map(D => \next_reg_c[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[9]\);
    
    \reg_a[27]\ : SLE
      port map(D => \next_reg_a[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[27]\);
    
    sum0_4_cry_0_974 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[19]\, C => 
        \R0_data[10]\, Y => \SIG0_0[29]\);
    
    next_reg_a_cry_0_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => sum0_4_cry_0_Y_0, B => oregs_ce_i_a2_0_a2, C
         => sum3_cry_0_Y, D => next_reg_H0_cry_0_0_Y, FCI => 
        GND_net_1, S => OPEN, Y => next_reg_a_cry_0_0_Y, FCO => 
        next_reg_a_cry_0);
    
    \next_reg_c[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(21), B => \R1_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[21]_net_1\);
    
    sum3_cry_21 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[21]\, B => Wt_data(21), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_20\, S => 
        \sum3[21]\, Y => OPEN, FCO => \sum3_cry_21\);
    
    sum0_4_axb_30 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[30]\, B => \R1_data[30]\, C => 
        \R0_data[30]\, D => \SIG0[30]_net_1\, Y => 
        \sum0_4_axb_30\);
    
    \SIG0[8]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[10]\, C => 
        \R0_data[21]\, Y => \SIG0[8]_net_1\);
    
    \reg_g[31]\ : SLE
      port map(D => \next_reg_g[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[31]\);
    
    \reg_d[3]\ : SLE
      port map(D => \next_reg_d[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[3]\);
    
    \SIG0[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[22]\, C => 
        \R0_data[11]\, Y => \SIG0[9]_net_1\);
    
    \reg_e[30]\ : SLE
      port map(D => \next_reg_e[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[30]\);
    
    sum3_6_0_cry_9 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[9]\, B => \R4_data[9]\, C => 
        \R5_data[9]\, D => \R6_data[9]\, FCI => \sum3_6_0_cry_8\, 
        S => \sum3_6_0[9]\, Y => OPEN, FCO => \sum3_6_0_cry_9\);
    
    \reg_e[4]\ : SLE
      port map(D => \next_reg_e[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[4]\);
    
    next_reg_e_cry_22_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[22]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(22), D => \R3_data[22]\, FCI => next_reg_e_cry_21, 
        S => \next_reg_e[22]\, Y => OPEN, FCO => 
        next_reg_e_cry_22);
    
    \next_reg_d[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(22), B => \R2_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[22]_net_1\);
    
    \reg_h[17]\ : SLE
      port map(D => \next_reg_h[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[17]\);
    
    \next_reg_g[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(16), B => \R5_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[16]_net_1\);
    
    sum0_4_cry_24 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[24]\, C => 
        \sum0_4_axb_24\, D => GND_net_1, FCI => \sum0_4_cry_23\, 
        S => \sum0_4[24]\, Y => OPEN, FCO => \sum0_4_cry_24\);
    
    \SIG0[27]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[17]\, C => 
        \R0_data[8]\, Y => \SIG0[27]_net_1\);
    
    sum0_4_axb_22 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[22]\, B => \R1_data[22]\, C => 
        \R0_data[22]\, D => \SIG0[22]_net_1\, Y => 
        \sum0_4_axb_22\);
    
    sum3_cry_5 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[5]\, B => Wt_data(5), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_4\, S => \sum3[5]\, Y
         => OPEN, FCO => \sum3_cry_5\);
    
    \next_reg_c[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(9), B => \R1_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[9]_net_1\);
    
    \reg_f[13]\ : SLE
      port map(D => \next_reg_f[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[13]\);
    
    \reg_c[5]\ : SLE
      port map(D => \next_reg_c[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[5]\);
    
    \reg_b[26]\ : SLE
      port map(D => \next_reg_b[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[26]\);
    
    \reg_h[23]\ : SLE
      port map(D => \next_reg_h[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[23]\);
    
    \next_reg_f[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[1]\, B => N5_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[1]_net_1\);
    
    \reg_d[6]\ : SLE
      port map(D => \next_reg_d[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[6]\);
    
    sum0_4_axb_25 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[25]\, B => \R1_data[25]\, C => 
        \R0_data[25]\, D => \SIG0[25]_net_1\, Y => 
        \sum0_4_axb_25\);
    
    \next_reg_h[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[1]\, B => N7_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[1]_net_1\);
    
    sum0_4_cry_0_1000 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[16]\, C => 
        \R0_data[5]\, Y => \SIG0_0[3]\);
    
    sum3_6_cry_7 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[7]\, B => \R4_data[0]\, C => 
        \R4_data[13]\, D => \R4_data[18]\, FCI => \sum3_6_cry_6\, 
        S => \sum3_6[7]\, Y => OPEN, FCO => \sum3_6_cry_7\);
    
    sum0_4_cry_0_985 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[20]\, C => 
        \R0_data[8]\, Y => \SIG0_0[18]\);
    
    \next_reg_b[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(28), B => \R0_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[28]_net_1\);
    
    sum3_6_cry_2 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[2]\, B => \R4_data[8]\, C => 
        \R4_data[13]\, D => \R4_data[27]\, FCI => \sum3_6_cry_1\, 
        S => \sum3_6[2]\, Y => OPEN, FCO => \sum3_6_cry_2\);
    
    \next_reg_h[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(26), B => \R6_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[26]_net_1\);
    
    sum3_6_cry_25 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[25]\, B => \R4_data[4]\, C => 
        \R4_data[18]\, D => \R4_data[31]\, FCI => \sum3_6_cry_24\, 
        S => \sum3_6[25]\, Y => OPEN, FCO => \sum3_6_cry_25\);
    
    \reg_d[4]\ : SLE
      port map(D => \next_reg_d[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[4]\);
    
    \reg_e[12]\ : SLE
      port map(D => \next_reg_e[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[12]\);
    
    \next_reg_c[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[6]\, B => N2_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[6]_net_1\);
    
    \reg_b[28]\ : SLE
      port map(D => \next_reg_b[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[28]\);
    
    \reg_e[11]\ : SLE
      port map(D => \next_reg_e[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[11]\);
    
    \next_reg_d[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(8), B => \R2_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[8]_net_1\);
    
    \next_reg_f[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(28), B => \R4_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[28]_net_1\);
    
    \next_reg_c[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(13), B => \R1_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[13]_net_1\);
    
    sum3_6_0_cry_29 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[29]\, B => \R4_data[29]\, C => 
        \R5_data[29]\, D => \R6_data[29]\, FCI => 
        \sum3_6_0_cry_28\, S => \sum3_6_0[29]\, Y => OPEN, FCO
         => \sum3_6_0_cry_29\);
    
    \reg_h[9]\ : SLE
      port map(D => \next_reg_h[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[9]\);
    
    \reg_f[14]\ : SLE
      port map(D => \next_reg_f[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[14]\);
    
    sum3_6_0_cry_15 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[15]\, B => \R4_data[15]\, C => 
        \R5_data[15]\, D => \R6_data[15]\, FCI => 
        \sum3_6_0_cry_14\, S => \sum3_6_0[15]\, Y => OPEN, FCO
         => \sum3_6_0_cry_15\);
    
    sum3_6_cry_17 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[17]\, B => \R4_data[10]\, C => 
        \R4_data[23]\, D => \R4_data[28]\, FCI => \sum3_6_cry_16\, 
        S => \sum3_6[17]\, Y => OPEN, FCO => \sum3_6_cry_17\);
    
    \reg_h[24]\ : SLE
      port map(D => \next_reg_h[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[24]\);
    
    \SIG0[20]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[10]\, B => \R0_data[1]\, C => 
        \R0_data[22]\, Y => \SIG0[20]_net_1\);
    
    \reg_g[29]\ : SLE
      port map(D => \next_reg_g[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[29]\);
    
    \reg_e[23]\ : SLE
      port map(D => \next_reg_e[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[23]\);
    
    sum0_4_cry_0_987 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[18]\, C => 
        \R0_data[6]\, Y => \SIG0_0[16]\);
    
    \next_reg_g[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[5]\, B => N6_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[5]_net_1\);
    
    \reg_a[30]\ : SLE
      port map(D => \next_reg_a[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[30]\);
    
    \next_reg_f[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(8), B => \R4_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[8]_net_1\);
    
    \reg_b[31]\ : SLE
      port map(D => \next_reg_b[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[31]\);
    
    \next_reg_f[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(7), B => \R4_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[7]_net_1\);
    
    \next_reg_h[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(19), B => \R6_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[19]_net_1\);
    
    \next_reg_g[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[2]\, B => N6_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[2]_net_1\);
    
    \reg_d[31]\ : SLE
      port map(D => \next_reg_d[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[31]\);
    
    \reg_e[16]\ : SLE
      port map(D => \next_reg_e[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[16]\);
    
    \reg_c[7]\ : SLE
      port map(D => \next_reg_c[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[7]\);
    
    next_reg_a_cry_1_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[1]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[1]\, D => N0_data(1), FCI => next_reg_a_cry_0, S
         => \next_reg_a[1]\, Y => OPEN, FCO => next_reg_a_cry_1);
    
    next_reg_e_cry_0_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => sum3_cry_0_Y, B => oregs_ce_i_a2_0_a2, C => 
        next_reg_H4_cry_0_0_Y, D => \R3_data[0]\, FCI => 
        GND_net_1, S => OPEN, Y => next_reg_e_cry_0_0_Y, FCO => 
        next_reg_e_cry_0);
    
    \next_reg_d[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(14), B => \R2_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[14]_net_1\);
    
    \reg_f[5]\ : SLE
      port map(D => \next_reg_f[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[5]\);
    
    sum0_4_cry_0_978 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[15]\, C => 
        \R0_data[6]\, Y => \SIG0_0[25]\);
    
    sum3_4_s_31 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \sum3_6[31]\, C => m325, D
         => GND_net_1, FCI => \sum3_4_cry_30\, S => \sum3_4[31]\, 
        Y => OPEN, FCO => OPEN);
    
    \next_reg_g[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(7), B => \R5_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[7]_net_1\);
    
    next_reg_e_cry_25_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[25]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(25), D => \R3_data[25]\, FCI => next_reg_e_cry_24, 
        S => \next_reg_e[25]\, Y => OPEN, FCO => 
        next_reg_e_cry_25);
    
    \next_reg_b[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(26), B => \R0_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[26]_net_1\);
    
    sum3_cry_9 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[9]\, B => Wt_data(9), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_8\, S => \sum3[9]\, Y
         => OPEN, FCO => \sum3_cry_9\);
    
    next_reg_e_cry_14_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[14]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(14), D => \R3_data[14]\, FCI => next_reg_e_cry_13, 
        S => \next_reg_e[14]\, Y => OPEN, FCO => 
        next_reg_e_cry_14);
    
    \reg_c[30]\ : SLE
      port map(D => \next_reg_c[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[30]\);
    
    sum0_4_cry_0_1001 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[24]\, B => \R0_data[15]\, C => 
        \R0_data[4]\, Y => \SIG0_0[2]\);
    
    \SIG0[28]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[18]\, C => 
        \R0_data[9]\, Y => \SIG0[28]_net_1\);
    
    \reg_e[24]\ : SLE
      port map(D => \next_reg_e[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[24]\);
    
    \reg_c[15]\ : SLE
      port map(D => \next_reg_c[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[15]\);
    
    \reg_h[31]\ : SLE
      port map(D => \next_reg_h[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[31]\);
    
    \next_reg_b[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(13), B => \R0_data[13]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[13]_net_1\);
    
    \reg_g[12]\ : SLE
      port map(D => \next_reg_g[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[12]\);
    
    \reg_e[18]\ : SLE
      port map(D => \next_reg_e[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[18]\);
    
    \reg_c[22]\ : SLE
      port map(D => \next_reg_c[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[22]\);
    
    \next_reg_f[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(26), B => \R4_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[26]_net_1\);
    
    \reg_g[11]\ : SLE
      port map(D => \next_reg_g[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[11]\);
    
    sum0_4_cry_11 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[11]\, C => 
        \sum0_4_axb_11\, D => GND_net_1, FCI => \sum0_4_cry_10\, 
        S => \sum0_4[11]\, Y => OPEN, FCO => \sum0_4_cry_11\);
    
    \reg_d[23]\ : SLE
      port map(D => \next_reg_d[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[23]\);
    
    \next_reg_b[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(31), B => \R0_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[31]_net_1\);
    
    \reg_c[21]\ : SLE
      port map(D => \next_reg_c[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[21]\);
    
    sum0_4_axb_3 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[3]\, B => \R1_data[3]\, C => 
        \R0_data[3]\, D => \SIG0[3]_net_1\, Y => \sum0_4_axb_3\);
    
    next_reg_a_cry_22_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[22]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[22]\, D => N0_data(22), FCI => next_reg_a_cry_21, S
         => \next_reg_a[22]\, Y => OPEN, FCO => next_reg_a_cry_22);
    
    \reg_b[0]\ : SLE
      port map(D => \next_reg_b[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[0]\);
    
    \next_reg_c[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(18), B => \R1_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[18]_net_1\);
    
    sum3_4_cry_0_971 : CFG4
      generic map(INIT => x"6996")

      port map(A => \R4_data[25]\, B => \R4_data[11]\, C => 
        \R4_data[6]\, D => sum3_6_0_cry_0_Y, Y => sum3_4_0);
    
    \next_reg_g[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(9), B => \R5_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[9]_net_1\);
    
    \reg_f[8]\ : SLE
      port map(D => \next_reg_f[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[8]\);
    
    next_reg_e_cry_19_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[19]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(19), D => \R3_data[19]\, FCI => next_reg_e_cry_18, 
        S => \next_reg_e[19]\, Y => OPEN, FCO => 
        next_reg_e_cry_19);
    
    sum0_4_cry_0_999 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[17]\, C => 
        \R0_data[6]\, Y => \SIG0_0[4]\);
    
    \next_reg_g[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(29), B => \R5_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[29]_net_1\);
    
    next_reg_e_cry_27_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[27]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(27), D => \R3_data[27]\, FCI => next_reg_e_cry_26, 
        S => \next_reg_e[27]\, Y => OPEN, FCO => 
        next_reg_e_cry_27);
    
    \next_reg_d[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(21), B => \R2_data[21]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[21]_net_1\);
    
    \SIG0[19]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[21]\, B => \R0_data[9]\, C => 
        \R0_data[0]\, Y => \SIG0[19]_net_1\);
    
    next_reg_e_cry_2_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[2]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(2), D => \R3_data[2]\, FCI => next_reg_e_cry_1, S
         => \next_reg_e[2]\, Y => OPEN, FCO => next_reg_e_cry_2);
    
    sum3_4_cry_8 : ARI1
      generic map(INIT => x"53AC5")

      port map(A => \sum3_6[8]\, B => m110_ns, C => m114, D => 
        Kt_addr(5), FCI => \sum3_4_cry_7\, S => \sum3_4[8]\, Y
         => OPEN, FCO => \sum3_4_cry_8\);
    
    sum0_4_cry_0_984 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[21]\, B => \R0_data[9]\, C => 
        \R0_data[0]\, Y => \SIG0_0[19]\);
    
    \reg_g[27]\ : SLE
      port map(D => \next_reg_g[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[27]\);
    
    sum3_6_cry_14 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[14]\, B => \R4_data[7]\, C => 
        \R4_data[20]\, D => \R4_data[25]\, FCI => \sum3_6_cry_13\, 
        S => \sum3_6[14]\, Y => OPEN, FCO => \sum3_6_cry_14\);
    
    sum0_4_axb_16 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[16]\, B => \R1_data[16]\, C => 
        \R0_data[16]\, D => \SIG0[16]_net_1\, Y => 
        \sum0_4_axb_16\);
    
    \reg_g[16]\ : SLE
      port map(D => \next_reg_g[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[16]\);
    
    sum0_4_axb_19 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[19]\, B => \R1_data[19]\, C => 
        \R0_data[19]\, D => \SIG0[19]_net_1\, Y => 
        \sum0_4_axb_19\);
    
    \reg_c[26]\ : SLE
      port map(D => \next_reg_c[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[26]\);
    
    \reg_d[24]\ : SLE
      port map(D => \next_reg_d[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[24]\);
    
    sum3_4_cry_17 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[17]\, B => m207_1_0, C => m207_1_1, D
         => Kt_addr(5), FCI => \sum3_4_cry_16\, S => \sum3_4[17]\, 
        Y => OPEN, FCO => \sum3_4_cry_17\);
    
    \next_reg_g[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[3]\, B => N6_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[3]_net_1\);
    
    \reg_f[19]\ : SLE
      port map(D => \next_reg_f[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[19]\);
    
    next_reg_a_cry_12_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[12]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[12]\, D => N0_data(12), FCI => next_reg_a_cry_11, S
         => \next_reg_a[12]\, Y => OPEN, FCO => next_reg_a_cry_12);
    
    \reg_h[29]\ : SLE
      port map(D => \next_reg_h[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[29]\);
    
    \reg_f[22]\ : SLE
      port map(D => \next_reg_f[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[22]\);
    
    next_reg_a_cry_6_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[6]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[6]\, D => N0_data(6), FCI => next_reg_a_cry_5, S
         => \next_reg_a[6]\, Y => OPEN, FCO => next_reg_a_cry_6);
    
    \reg_f[21]\ : SLE
      port map(D => \next_reg_f[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[21]\);
    
    sum3_cry_12 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[12]\, B => Wt_data(12), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_11\, S => 
        \sum3[12]\, Y => OPEN, FCO => \sum3_cry_12\);
    
    \next_reg_c[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(30), B => \R1_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[30]_net_1\);
    
    sum0_4_cry_0_981 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[24]\, B => \R0_data[3]\, C => 
        \R0_data[12]\, Y => \SIG0_0[22]\);
    
    \reg_g[18]\ : SLE
      port map(D => \next_reg_g[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[18]\);
    
    sum0_4_axb_8 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[8]\, B => \R1_data[8]\, C => 
        \R0_data[8]\, D => \SIG0[8]_net_1\, Y => \sum0_4_axb_8\);
    
    \reg_c[28]\ : SLE
      port map(D => \next_reg_c[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[28]\);
    
    sum3_6_0_cry_4 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[4]\, B => \R4_data[4]\, C => 
        \R5_data[4]\, D => \R6_data[4]\, FCI => \sum3_6_0_cry_3\, 
        S => \sum3_6_0[4]\, Y => OPEN, FCO => \sum3_6_0_cry_4\);
    
    \next_reg_b[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(18), B => \R0_data[18]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[18]_net_1\);
    
    next_reg_a_cry_8_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[8]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[8]\, D => N0_data(8), FCI => next_reg_a_cry_7, S
         => \next_reg_a[8]\, Y => OPEN, FCO => next_reg_a_cry_8);
    
    sum3_6_0_cry_18 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[18]\, B => \R4_data[18]\, C => 
        \R5_data[18]\, D => \R6_data[18]\, FCI => 
        \sum3_6_0_cry_17\, S => \sum3_6_0[18]\, Y => OPEN, FCO
         => \sum3_6_0_cry_18\);
    
    \next_reg_c[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(16), B => \R1_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[16]_net_1\);
    
    \next_reg_d[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(17), B => \R2_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[17]_net_1\);
    
    sum0_4_axb_11 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[11]\, B => \R1_data[11]\, C => 
        \R0_data[11]\, D => \SIG0[11]_net_1\, Y => 
        \sum0_4_axb_11\);
    
    sum0_4_cry_2 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[2]\, C => 
        \sum0_4_axb_2\, D => GND_net_1, FCI => \sum0_4_cry_1\, S
         => \sum0_4[2]\, Y => OPEN, FCO => \sum0_4_cry_2\);
    
    sum0_4_cry_25 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[25]\, C => 
        \sum0_4_axb_25\, D => GND_net_1, FCI => \sum0_4_cry_24\, 
        S => \sum0_4[25]\, Y => OPEN, FCO => \sum0_4_cry_25\);
    
    \next_reg_d[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(15), B => \R2_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[15]_net_1\);
    
    \reg_c[10]\ : SLE
      port map(D => \next_reg_c[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[10]\);
    
    \next_reg_c[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(23), B => \R1_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[23]_net_1\);
    
    \reg_d[15]\ : SLE
      port map(D => \next_reg_d[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[15]\);
    
    \reg_a[5]\ : SLE
      port map(D => \next_reg_a[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[5]\);
    
    sum0_4_cry_0_982 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[11]\, C => 
        \R0_data[2]\, Y => \SIG0_0[21]\);
    
    \reg_b[1]\ : SLE
      port map(D => \next_reg_b[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[1]\);
    
    \reg_b[12]\ : SLE
      port map(D => \next_reg_b[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[12]\);
    
    \SIG0[2]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[24]\, B => \R0_data[15]\, C => 
        \R0_data[4]\, Y => \SIG0[2]_net_1\);
    
    sum0_4_axb_23 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[23]\, B => \R1_data[23]\, C => 
        \R0_data[23]\, D => \SIG0[23]_net_1\, Y => 
        \sum0_4_axb_23\);
    
    \next_reg_d[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(30), B => \R2_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[30]_net_1\);
    
    sum0_4_axb_5 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[5]\, B => \R1_data[5]\, C => 
        \R0_data[5]\, D => \SIG0[5]_net_1\, Y => \sum0_4_axb_5\);
    
    \reg_b[11]\ : SLE
      port map(D => \next_reg_b[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[11]\);
    
    \reg_f[26]\ : SLE
      port map(D => \next_reg_f[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[26]\);
    
    next_reg_e_cry_10_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[10]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(10), D => \R3_data[10]\, FCI => next_reg_e_cry_9, 
        S => \next_reg_e[10]\, Y => OPEN, FCO => 
        next_reg_e_cry_10);
    
    \reg_e[29]\ : SLE
      port map(D => \next_reg_e[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[29]\);
    
    \next_reg_b[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[2]\, B => N1_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[2]_net_1\);
    
    sum3_cry_8 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[8]\, B => Wt_data(8), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_7\, S => \sum3[8]\, Y
         => OPEN, FCO => \sum3_cry_8\);
    
    sum3_cry_23 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[23]\, B => Wt_data(23), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_22\, S => 
        \sum3[23]\, Y => OPEN, FCO => \sum3_cry_23\);
    
    sum0_4_axb_20 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[20]\, B => \R1_data[20]\, C => 
        \R0_data[20]\, D => \SIG0[20]_net_1\, Y => 
        \sum0_4_axb_20\);
    
    sum0_4_cry_0_973 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[20]\, B => \R0_data[11]\, C => 
        \R0_data[0]\, Y => \SIG0_0[30]\);
    
    next_reg_a_cry_25_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[25]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[25]\, D => N0_data(25), FCI => next_reg_a_cry_24, S
         => \next_reg_a[25]\, Y => OPEN, FCO => next_reg_a_cry_25);
    
    \next_reg_f[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(19), B => \R4_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[19]_net_1\);
    
    sum3_4_cry_21 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[21]\, B => m235_ns, C => m239, D => 
        Kt_addr(5), FCI => \sum3_4_cry_20\, S => \sum3_4[21]\, Y
         => OPEN, FCO => \sum3_4_cry_21\);
    
    \Maj[31]\ : CFG3
      generic map(INIT => x"E8")

      port map(A => \R2_data[31]\, B => \R1_data[31]\, C => 
        \R0_data[31]\, Y => \Maj[31]_net_1\);
    
    \SIG0[13]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[15]\, C => 
        \R0_data[3]\, Y => \SIG0[13]_net_1\);
    
    sum0_4_axb_12 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[12]\, B => \R1_data[12]\, C => 
        \R0_data[12]\, D => \SIG0[12]_net_1\, Y => 
        \sum0_4_axb_12\);
    
    sum3_cry_6 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[6]\, B => Wt_data(6), C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_cry_5\, S => \sum3[6]\, Y
         => OPEN, FCO => \sum3_cry_6\);
    
    \reg_f[28]\ : SLE
      port map(D => \next_reg_f[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[28]\);
    
    \reg_f[17]\ : SLE
      port map(D => \next_reg_f[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[17]\);
    
    sum3_4_cry_14 : ARI1
      generic map(INIT => x"5C53A")

      port map(A => \sum3_6[14]\, B => m172_ns, C => m177, D => 
        Kt_addr(5), FCI => \sum3_4_cry_13\, S => \sum3_4[14]\, Y
         => OPEN, FCO => \sum3_4_cry_14\);
    
    \reg_h[27]\ : SLE
      port map(D => \next_reg_h[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[27]\);
    
    \reg_b[16]\ : SLE
      port map(D => \next_reg_b[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[16]\);
    
    sum0_4_axb_15 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[15]\, B => \R1_data[15]\, C => 
        \R0_data[15]\, D => \SIG0[15]_net_1\, Y => 
        \sum0_4_axb_15\);
    
    \next_reg_b[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(16), B => \R0_data[16]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[16]_net_1\);
    
    \next_reg_h[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(14), B => \R6_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[14]_net_1\);
    
    sum0_4_cry_0_988 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[17]\, C => 
        \R0_data[5]\, Y => \SIG0_0[15]\);
    
    sum0_4_axb_9 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[9]\, B => \R1_data[9]\, C => 
        \R0_data[9]\, D => \SIG0[9]_net_1\, Y => \sum0_4_axb_9\);
    
    next_reg_a_cry_27_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[27]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[27]\, D => N0_data(27), FCI => next_reg_a_cry_26, S
         => \next_reg_a[27]\, Y => OPEN, FCO => next_reg_a_cry_27);
    
    next_reg_a_cry_15_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[15]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[15]\, D => N0_data(15), FCI => next_reg_a_cry_14, S
         => \next_reg_a[15]\, Y => OPEN, FCO => next_reg_a_cry_15);
    
    sum0_4_cry_0_976 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[29]\, B => \R0_data[17]\, C => 
        \R0_data[8]\, Y => \SIG0_0[27]\);
    
    \reg_d[29]\ : SLE
      port map(D => \next_reg_d[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[29]\);
    
    sum0_4_cry_5 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[5]\, C => 
        \sum0_4_axb_5\, D => GND_net_1, FCI => \sum0_4_cry_4\, S
         => \sum0_4[5]\, Y => OPEN, FCO => \sum0_4_cry_5\);
    
    next_reg_e_cry_1_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[1]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(1), D => \R3_data[1]\, FCI => next_reg_e_cry_0, S
         => \next_reg_e[1]\, Y => OPEN, FCO => next_reg_e_cry_1);
    
    \reg_b[9]\ : SLE
      port map(D => \next_reg_b[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[9]\);
    
    \next_reg_c[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(28), B => \R1_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[28]_net_1\);
    
    \reg_b[18]\ : SLE
      port map(D => \next_reg_b[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[18]\);
    
    \next_reg_g[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(19), B => \R5_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[19]_net_1\);
    
    sum0_4_cry_10 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[10]\, C => 
        \sum0_4_axb_10\, D => GND_net_1, FCI => \sum0_4_cry_9\, S
         => \sum0_4[10]\, Y => OPEN, FCO => \sum0_4_cry_10\);
    
    sum3_6_0_cry_8 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[8]\, B => \R4_data[8]\, C => 
        \R5_data[8]\, D => \R6_data[8]\, FCI => \sum3_6_0_cry_7\, 
        S => \sum3_6_0[8]\, Y => OPEN, FCO => \sum3_6_0_cry_8\);
    
    \next_reg_c[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[0]\, B => next_reg_H2_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_c[0]_net_1\);
    
    \reg_d[7]\ : SLE
      port map(D => \next_reg_d[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[7]\);
    
    \next_reg_d[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(10), B => \R2_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[10]_net_1\);
    
    \reg_d[10]\ : SLE
      port map(D => \next_reg_d[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[10]\);
    
    \SIG0[21]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[11]\, C => 
        \R0_data[2]\, Y => \SIG0[21]_net_1\);
    
    next_reg_e_cry_6_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[6]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(6), D => \R3_data[6]\, FCI => next_reg_e_cry_5, S
         => \next_reg_e[6]\, Y => OPEN, FCO => next_reg_e_cry_6);
    
    sum3_4_cry_9 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[9]\, B => m119_ns, C => m124, D => 
        Kt_addr(5), FCI => \sum3_4_cry_8\, S => \sum3_4[9]\, Y
         => OPEN, FCO => \sum3_4_cry_9\);
    
    \reg_e[27]\ : SLE
      port map(D => \next_reg_e[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[27]\);
    
    \reg_b[25]\ : SLE
      port map(D => \next_reg_b[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[25]\);
    
    \reg_g[3]\ : SLE
      port map(D => \next_reg_g[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[3]\);
    
    \next_reg_c[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[3]\, B => N2_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[3]_net_1\);
    
    next_reg_a_cry_17_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[17]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[17]\, D => N0_data(17), FCI => next_reg_a_cry_16, S
         => \next_reg_a[17]\, Y => OPEN, FCO => next_reg_a_cry_17);
    
    next_reg_e_cry_24_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[24]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(24), D => \R3_data[24]\, FCI => next_reg_e_cry_23, 
        S => \next_reg_e[24]\, Y => OPEN, FCO => 
        next_reg_e_cry_24);
    
    \next_reg_g[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(24), B => \R5_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[24]_net_1\);
    
    sum0_4_axb_0 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[0]\, B => \R1_data[0]\, C => 
        \R0_data[0]\, D => sum0_4, Y => \sum0_4[0]\);
    
    \next_reg_h[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(29), B => \R6_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[29]_net_1\);
    
    \reg_h[3]\ : SLE
      port map(D => \next_reg_h[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[3]\);
    
    next_reg_e_cry_13_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[13]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(13), D => \R3_data[13]\, FCI => next_reg_e_cry_12, 
        S => \next_reg_e[13]\, Y => OPEN, FCO => 
        next_reg_e_cry_13);
    
    sum0_4_cry_13 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[13]\, C => 
        \sum0_4_axb_13\, D => GND_net_1, FCI => \sum0_4_cry_12\, 
        S => \sum0_4[13]\, Y => OPEN, FCO => \sum0_4_cry_13\);
    
    sum0_4_axb_4 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[4]\, B => \R1_data[4]\, C => 
        \R0_data[4]\, D => \SIG0[4]_net_1\, Y => \sum0_4_axb_4\);
    
    sum0_4_cry_0_995 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[10]\, C => 
        \R0_data[21]\, Y => \SIG0_0[8]\);
    
    \reg_g[2]\ : SLE
      port map(D => \next_reg_g[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[2]\);
    
    \next_reg_d[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(12), B => \R2_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[12]_net_1\);
    
    sum3_s_31 : ARI1
      generic map(INIT => x"46600")

      port map(A => VCC_net_1, B => \sum3_4[31]\, C => 
        Wt_data(31), D => GND_net_1, FCI => \sum3_cry_30\, S => 
        \sum3[31]\, Y => OPEN, FCO => OPEN);
    
    sum3_6_0_cry_23 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[23]\, B => \R4_data[23]\, C => 
        \R5_data[23]\, D => \R6_data[23]\, FCI => 
        \sum3_6_0_cry_22\, S => \sum3_6_0[23]\, Y => OPEN, FCO
         => \sum3_6_0_cry_23\);
    
    sum3_6_cry_3 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[3]\, B => \R4_data[9]\, C => 
        \R4_data[14]\, D => \R4_data[28]\, FCI => \sum3_6_cry_2\, 
        S => \sum3_6[3]\, Y => OPEN, FCO => \sum3_6_cry_3\);
    
    sum3_6_0_cry_12 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[12]\, B => \R4_data[12]\, C => 
        \R5_data[12]\, D => \R6_data[12]\, FCI => 
        \sum3_6_0_cry_11\, S => \sum3_6_0[12]\, Y => OPEN, FCO
         => \sum3_6_0_cry_12\);
    
    \next_reg_f[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[2]\, B => N5_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[2]_net_1\);
    
    \SIG0[17]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[19]\, C => 
        \R0_data[7]\, Y => \SIG0[17]_net_1\);
    
    \reg_h[1]\ : SLE
      port map(D => \next_reg_h[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[1]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    sum3_6_cry_1 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[1]\, B => \R4_data[7]\, C => 
        \R4_data[12]\, D => \R4_data[26]\, FCI => \sum3_6_cry_0\, 
        S => \sum3_6[1]\, Y => OPEN, FCO => \sum3_6_cry_1\);
    
    \next_reg_d[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[5]\, B => N3_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[5]_net_1\);
    
    sum3_6_cry_15 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[15]\, B => \R4_data[8]\, C => 
        \R4_data[21]\, D => \R4_data[26]\, FCI => \sum3_6_cry_14\, 
        S => \sum3_6[15]\, Y => OPEN, FCO => \sum3_6_cry_15\);
    
    sum0_4_cry_18 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[18]\, C => 
        \sum0_4_axb_18\, D => GND_net_1, FCI => \sum0_4_cry_17\, 
        S => \sum0_4[18]\, Y => OPEN, FCO => \sum0_4_cry_18\);
    
    \reg_c[13]\ : SLE
      port map(D => \next_reg_c[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[13]\);
    
    \next_reg_c[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(26), B => \R1_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[26]_net_1\);
    
    next_reg_e_cry_29_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[29]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(29), D => \R3_data[29]\, FCI => next_reg_e_cry_28, 
        S => \next_reg_e[29]\, Y => OPEN, FCO => 
        next_reg_e_cry_29);
    
    \next_reg_h[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[2]\, B => N7_data(2), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[2]_net_1\);
    
    \next_reg_b[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(8), B => \R0_data[8]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[8]_net_1\);
    
    sum3_6_cry_21 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[21]\, B => \R4_data[0]\, C => 
        \R4_data[14]\, D => \R4_data[27]\, FCI => \sum3_6_cry_20\, 
        S => \sum3_6[21]\, Y => OPEN, FCO => \sum3_6_cry_21\);
    
    sum0_4_axb_2 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[2]\, B => \R1_data[2]\, C => 
        \R0_data[2]\, D => \SIG0[2]_net_1\, Y => \sum0_4_axb_2\);
    
    \reg_d[27]\ : SLE
      port map(D => \next_reg_d[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[27]\);
    
    sum0_4_axb_7 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[7]\, B => \R1_data[7]\, C => 
        \R0_data[7]\, D => \SIG0[7]_net_1\, Y => \sum0_4_axb_7\);
    
    \next_reg_d[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(23), B => \R2_data[23]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[23]_net_1\);
    
    \next_reg_c[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(31), B => \R1_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[31]_net_1\);
    
    \reg_a[12]\ : SLE
      port map(D => \next_reg_a[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[12]\);
    
    \next_reg_h[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(17), B => \R6_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[17]_net_1\);
    
    sum0_4_cry_0_997 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[28]\, B => \R0_data[19]\, C => 
        \R0_data[8]\, Y => \SIG0_0[6]\);
    
    \reg_a[11]\ : SLE
      port map(D => \next_reg_a[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[11]\);
    
    \next_reg_h[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[4]\, B => N7_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[4]_net_1\);
    
    \next_reg_h[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(15), B => \R6_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[15]_net_1\);
    
    sum3_6_cry_0 : ARI1
      generic map(INIT => x"56996")

      port map(A => sum3_6_0_cry_0_Y, B => \R4_data[6]\, C => 
        \R4_data[11]\, D => \R4_data[25]\, FCI => GND_net_1, S
         => OPEN, Y => sum3_6_cry_0_Y, FCO => \sum3_6_cry_0\);
    
    \reg_e[15]\ : SLE
      port map(D => \next_reg_e[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[15]\);
    
    \reg_a[22]\ : SLE
      port map(D => \next_reg_a[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[22]\);
    
    \next_reg_b[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[4]\, B => N1_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[4]_net_1\);
    
    sum0_4_axb_24 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[24]\, B => \R1_data[24]\, C => 
        \R0_data[24]\, D => \SIG0[24]_net_1\, Y => 
        \sum0_4_axb_24\);
    
    \reg_a[21]\ : SLE
      port map(D => \next_reg_a[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[21]\);
    
    sum3_cry_20 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[20]\, B => Wt_data(20), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_19\, S => 
        \sum3[20]\, Y => OPEN, FCO => \sum3_cry_20\);
    
    sum3_cry_11 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[11]\, B => Wt_data(11), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_10\, S => 
        \sum3[11]\, Y => OPEN, FCO => \sum3_cry_11\);
    
    \next_reg_b[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(29), B => \R0_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[29]_net_1\);
    
    \next_reg_f[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[4]\, B => N5_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[4]_net_1\);
    
    \reg_e[7]\ : SLE
      port map(D => \next_reg_e[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[7]\);
    
    sum3_6_0_cry_17 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[17]\, B => \R4_data[17]\, C => 
        \R5_data[17]\, D => \R6_data[17]\, FCI => 
        \sum3_6_0_cry_16\, S => \sum3_6_0[17]\, Y => OPEN, FCO
         => \sum3_6_0_cry_17\);
    
    \reg_c[14]\ : SLE
      port map(D => \next_reg_c[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[14]\);
    
    sum0_4_cry_0_983 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[10]\, B => \R0_data[1]\, C => 
        \R0_data[22]\, Y => \SIG0_0[20]\);
    
    \SIG0[10]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[23]\, B => \R0_data[0]\, C => 
        \R0_data[12]\, Y => \SIG0[10]_net_1\);
    
    next_reg_a_s_31 : ARI1
      generic map(INIT => x"47D28")

      port map(A => N0_data(31), B => oregs_ce_i_a2_0_a2, C => 
        \sum0_4[31]\, D => \sum3[31]\, FCI => next_reg_a_cry_30, 
        S => \next_reg_a[31]\, Y => OPEN, FCO => OPEN);
    
    \next_reg_d[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(31), B => \R2_data[31]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[31]_net_1\);
    
    \reg_b[20]\ : SLE
      port map(D => \next_reg_b[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[20]\);
    
    sum3_4_cry_20 : ARI1
      generic map(INIT => x"5C53A")

      port map(A => \sum3_6[20]\, B => m226_ns, C => m230, D => 
        Kt_addr(5), FCI => \sum3_4_cry_19\, S => \sum3_4[20]\, Y
         => OPEN, FCO => \sum3_4_cry_20\);
    
    \SIG0[24]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[26]\, B => \R0_data[14]\, C => 
        \R0_data[5]\, Y => \SIG0[24]_net_1\);
    
    \next_reg_f[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(29), B => \R4_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[29]_net_1\);
    
    \reg_h[12]\ : SLE
      port map(D => \next_reg_h[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[12]\);
    
    \next_reg_f[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(14), B => \R4_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[14]_net_1\);
    
    next_reg_e_cry_7_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[7]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(7), D => \R3_data[7]\, FCI => next_reg_e_cry_6, S
         => \next_reg_e[7]\, Y => OPEN, FCO => next_reg_e_cry_7);
    
    next_reg_a_cry_3_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[3]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[3]\, D => N0_data(3), FCI => next_reg_a_cry_2, S
         => \next_reg_a[3]\, Y => OPEN, FCO => next_reg_a_cry_3);
    
    \reg_h[11]\ : SLE
      port map(D => \next_reg_h[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[11]\);
    
    sum0_4_axb_27 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[27]\, B => \R1_data[27]\, C => 
        \R0_data[27]\, D => \SIG0[27]_net_1\, Y => 
        \sum0_4_axb_27\);
    
    \reg_a[16]\ : SLE
      port map(D => \next_reg_a[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[16]\);
    
    \reg_a[3]\ : SLE
      port map(D => \next_reg_a[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[3]\);
    
    \next_reg_d[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(9), B => \R2_data[9]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[9]_net_1\);
    
    \reg_g[30]\ : SLE
      port map(D => \next_reg_g[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[30]\);
    
    \reg_g[4]\ : SLE
      port map(D => \next_reg_g[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[4]\);
    
    sum3_4_cry_7 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[7]\, B => m104_am, C => m104_bm, D
         => Kt_addr(5), FCI => \sum3_4_cry_6\, S => \sum3_4[7]\, 
        Y => OPEN, FCO => \sum3_4_cry_7\);
    
    \next_reg_d[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[3]\, B => N3_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[3]_net_1\);
    
    \reg_a[26]\ : SLE
      port map(D => \next_reg_a[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[26]\);
    
    \next_reg_g[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(27), B => \R5_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[27]_net_1\);
    
    \next_reg_g[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(25), B => \R5_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[25]_net_1\);
    
    next_reg_e_cry_20_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[20]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(20), D => \R3_data[20]\, FCI => next_reg_e_cry_19, 
        S => \next_reg_e[20]\, Y => OPEN, FCO => 
        next_reg_e_cry_20);
    
    sum0_4_cry_30 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[30]\, C => 
        \sum0_4_axb_30\, D => GND_net_1, FCI => \sum0_4_cry_29\, 
        S => \sum0_4[30]\, Y => OPEN, FCO => \sum0_4_cry_30\);
    
    \next_reg_c[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R1_data[1]\, B => N2_data(1), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[1]_net_1\);
    
    sum3_4_cry_23 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[23]\, B => m254, C => m258_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_22\, S => \sum3_4[23]\, Y
         => OPEN, FCO => \sum3_4_cry_23\);
    
    \reg_a[7]\ : SLE
      port map(D => \next_reg_a[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[7]\);
    
    sum0_4_cry_0_986 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[30]\, B => \R0_data[19]\, C => 
        \R0_data[7]\, Y => \SIG0_0[17]\);
    
    \SIG0[18]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[20]\, C => 
        \R0_data[8]\, Y => \SIG0[18]_net_1\);
    
    \reg_a[18]\ : SLE
      port map(D => \next_reg_a[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[18]\);
    
    \reg_e[6]\ : SLE
      port map(D => \next_reg_e[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[6]\);
    
    \next_reg_d[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(28), B => \R2_data[28]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[28]_net_1\);
    
    \reg_d[13]\ : SLE
      port map(D => \next_reg_d[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[13]\);
    
    next_reg_a_cry_24_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[24]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[24]\, D => N0_data(24), FCI => next_reg_a_cry_23, S
         => \next_reg_a[24]\, Y => OPEN, FCO => next_reg_a_cry_24);
    
    sum0_4_cry_0_994 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[31]\, B => \R0_data[22]\, C => 
        \R0_data[11]\, Y => \SIG0_0[9]\);
    
    \reg_h[16]\ : SLE
      port map(D => \next_reg_h[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[16]\);
    
    sum3_4_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \sum3_6[1]\, B => m34, C => GND_net_1, D => 
        GND_net_1, FCI => \sum3_4_cry_0\, S => \sum3_4[1]\, Y => 
        OPEN, FCO => \sum3_4_cry_1\);
    
    sum0_4_axb_13 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[13]\, B => \R1_data[13]\, C => 
        \R0_data[13]\, D => \SIG0[13]_net_1\, Y => 
        \sum0_4_axb_13\);
    
    \reg_c[6]\ : SLE
      port map(D => \next_reg_c[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[6]\);
    
    sum3_4_cry_15 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_6[15]\, B => Kt_data_0, C => GND_net_1, 
        D => GND_net_1, FCI => \sum3_4_cry_14\, S => \sum3_4[15]\, 
        Y => OPEN, FCO => \sum3_4_cry_15\);
    
    sum3_4_cry_0 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => sum3_4_0, C => \sum3_4[0]\, D
         => GND_net_1, FCI => GND_net_1, S => OPEN, Y => 
        sum3_4_cry_0_Y, FCO => \sum3_4_cry_0\);
    
    \next_reg_f[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[3]\, B => N5_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[3]_net_1\);
    
    \reg_g[15]\ : SLE
      port map(D => \next_reg_g[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[15]\);
    
    sum0_4_cry_19 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[19]\, C => 
        \sum0_4_axb_19\, D => GND_net_1, FCI => \sum0_4_cry_18\, 
        S => \sum0_4[19]\, Y => OPEN, FCO => \sum0_4_cry_19\);
    
    \reg_a[28]\ : SLE
      port map(D => \next_reg_a[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[28]\);
    
    \reg_c[25]\ : SLE
      port map(D => \next_reg_c[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[25]\);
    
    sum0_4_axb_10 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[10]\, B => \R1_data[10]\, C => 
        \R0_data[10]\, D => \SIG0[10]_net_1\, Y => 
        \sum0_4_axb_10\);
    
    \reg_c[3]\ : SLE
      port map(D => \next_reg_c[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[3]\);
    
    sum3_4_cry_28 : ARI1
      generic map(INIT => x"53AC5")

      port map(A => \sum3_6[28]\, B => m296, C => m300_ns, D => 
        Kt_addr(5), FCI => \sum3_4_cry_27\, S => \sum3_4[28]\, Y
         => OPEN, FCO => \sum3_4_cry_28\);
    
    sum3_6_0_cry_0 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[0]\, B => \R4_data[0]\, C => 
        \R5_data[0]\, D => \R6_data[0]\, FCI => GND_net_1, S => 
        OPEN, Y => sum3_6_0_cry_0_Y, FCO => \sum3_6_0_cry_0\);
    
    \next_reg_g[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(14), B => \R5_data[14]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[14]_net_1\);
    
    \SIG0[25]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[15]\, C => 
        \R0_data[6]\, Y => \SIG0[25]_net_1\);
    
    \next_reg_h[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[3]\, B => N7_data(3), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[3]_net_1\);
    
    \next_reg_b[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R0_data[6]\, B => N1_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[6]_net_1\);
    
    sum0_4_cry_16 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[16]\, C => 
        \sum0_4_axb_16\, D => GND_net_1, FCI => \sum0_4_cry_15\, 
        S => \sum0_4[16]\, Y => OPEN, FCO => \sum0_4_cry_16\);
    
    \next_reg_h[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(10), B => \R6_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[10]_net_1\);
    
    sum3_cry_29 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[29]\, B => Wt_data(29), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_28\, S => 
        \sum3[29]\, Y => OPEN, FCO => \sum3_cry_29\);
    
    \reg_e[10]\ : SLE
      port map(D => \next_reg_e[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[10]\);
    
    next_reg_e_s_31 : ARI1
      generic map(INIT => x"472D8")

      port map(A => \R3_data[31]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[31]\, D => N4_data(31), FCI => next_reg_e_cry_30, S
         => \next_reg_e[31]\, Y => OPEN, FCO => OPEN);
    
    sum3_cry_28 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[28]\, B => Wt_data(28), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_27\, S => 
        \sum3[28]\, Y => OPEN, FCO => \sum3_cry_28\);
    
    \reg_h[18]\ : SLE
      port map(D => \next_reg_h[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[18]\);
    
    next_reg_a_cry_29_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[29]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[29]\, D => N0_data(29), FCI => next_reg_a_cry_28, S
         => \next_reg_a[29]\, Y => OPEN, FCO => next_reg_a_cry_29);
    
    sum3_6_s_31 : ARI1
      generic map(INIT => x"46996")

      port map(A => \R4_data[24]\, B => \sum3_6_0[31]\, C => 
        \R4_data[5]\, D => \R4_data[10]\, FCI => \sum3_6_cry_30\, 
        S => \sum3_6[31]\, Y => OPEN, FCO => OPEN);
    
    \next_reg_d[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(11), B => \R2_data[11]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[11]_net_1\);
    
    \next_reg_c[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(19), B => \R1_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[19]_net_1\);
    
    sum0_4_cry_0_991 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[14]\, C => 
        \R0_data[2]\, Y => \SIG0_0[12]\);
    
    \reg_c[1]\ : SLE
      port map(D => \next_reg_c[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[1]\);
    
    \next_reg_h[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(7), B => \R6_data[7]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[7]_net_1\);
    
    \reg_h[6]\ : SLE
      port map(D => \next_reg_h[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[6]\);
    
    \reg_d[14]\ : SLE
      port map(D => \next_reg_d[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[14]\);
    
    next_reg_a_cry_14_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[14]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[14]\, D => N0_data(14), FCI => next_reg_a_cry_13, S
         => \next_reg_a[14]\, Y => OPEN, FCO => next_reg_a_cry_14);
    
    next_reg_a_cry_2_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[2]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[2]\, D => N0_data(2), FCI => next_reg_a_cry_1, S
         => \next_reg_a[2]\, Y => OPEN, FCO => next_reg_a_cry_2);
    
    \reg_g[0]\ : SLE
      port map(D => \next_reg_g[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[0]\);
    
    \next_reg_h[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(24), B => \R6_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[24]_net_1\);
    
    \reg_h[2]\ : SLE
      port map(D => \next_reg_h[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[2]\);
    
    \reg_b[30]\ : SLE
      port map(D => \next_reg_b[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[30]\);
    
    \reg_c[19]\ : SLE
      port map(D => \next_reg_c[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[19]\);
    
    \next_reg_h[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(12), B => \R6_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[12]_net_1\);
    
    sum3_6_cry_9 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[9]\, B => \R4_data[2]\, C => 
        \R4_data[15]\, D => \R4_data[20]\, FCI => \sum3_6_cry_8\, 
        S => \sum3_6[9]\, Y => OPEN, FCO => \sum3_6_cry_9\);
    
    \next_reg_d[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N3_data(26), B => \R2_data[26]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[26]_net_1\);
    
    \reg_d[30]\ : SLE
      port map(D => \next_reg_d[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[30]\);
    
    sum3_6_0_cry_19 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[19]\, B => \R4_data[19]\, C => 
        \R5_data[19]\, D => \R6_data[19]\, FCI => 
        \sum3_6_0_cry_18\, S => \sum3_6_0[19]\, Y => OPEN, FCO
         => \sum3_6_0_cry_19\);
    
    sum0_4_cry_0_992 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[13]\, B => \R0_data[1]\, C => 
        \R0_data[24]\, Y => \SIG0_0[11]\);
    
    \reg_f[25]\ : SLE
      port map(D => \next_reg_f[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[25]\);
    
    \next_reg_f[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(17), B => \R4_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[17]_net_1\);
    
    \next_reg_h[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R6_data[0]\, B => next_reg_H7_cry_0_0_Y, C
         => oregs_ce_i_a2_0_a2, Y => \next_reg_h[0]_net_1\);
    
    \next_reg_f[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(15), B => \R4_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[15]_net_1\);
    
    sum0_4_cry_21 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[21]\, C => 
        \sum0_4_axb_21\, D => GND_net_1, FCI => \sum0_4_cry_20\, 
        S => \sum0_4[21]\, Y => OPEN, FCO => \sum0_4_cry_21\);
    
    sum0_4_cry_12 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[12]\, C => 
        \sum0_4_axb_12\, D => GND_net_1, FCI => \sum0_4_cry_11\, 
        S => \sum0_4[12]\, Y => OPEN, FCO => \sum0_4_cry_12\);
    
    sum3_6_0_cry_20 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[20]\, B => \R4_data[20]\, C => 
        \R5_data[20]\, D => \R6_data[20]\, FCI => 
        \sum3_6_0_cry_19\, S => \sum3_6_0[20]\, Y => OPEN, FCO
         => \sum3_6_0_cry_20\);
    
    sum3_cry_0 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \Wt_data_0[0]\, C => 
        \sum3[0]\, D => GND_net_1, FCI => GND_net_1, S => OPEN, Y
         => sum3_cry_0_Y, FCO => \sum3_cry_0\);
    
    sum3_6_0_cry_26 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[26]\, B => \R4_data[26]\, C => 
        \R5_data[26]\, D => \R6_data[26]\, FCI => 
        \sum3_6_0_cry_25\, S => \sum3_6_0[26]\, Y => OPEN, FCO
         => \sum3_6_0_cry_26\);
    
    sum0_4_cry_9 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \SIG0_0[9]\, C => 
        \sum0_4_axb_9\, D => GND_net_1, FCI => \sum0_4_cry_8\, S
         => \sum0_4[9]\, Y => OPEN, FCO => \sum0_4_cry_9\);
    
    next_reg_a_cry_19_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[19]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[19]\, D => N0_data(19), FCI => next_reg_a_cry_18, S
         => \next_reg_a[19]\, Y => OPEN, FCO => next_reg_a_cry_19);
    
    \reg_g[8]\ : SLE
      port map(D => \next_reg_g[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[8]\);
    
    \reg_d[1]\ : SLE
      port map(D => \next_reg_d[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[1]\);
    
    sum3_6_cry_20 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[20]\, B => \R4_data[13]\, C => 
        \R4_data[26]\, D => \R4_data[31]\, FCI => \sum3_6_cry_19\, 
        S => \sum3_6[20]\, Y => OPEN, FCO => \sum3_6_cry_20\);
    
    \next_reg_g[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(20), B => \R5_data[20]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[20]_net_1\);
    
    \next_reg_g[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(30), B => \R5_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[30]_net_1\);
    
    \reg_b[8]\ : SLE
      port map(D => \next_reg_b[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[8]\);
    
    next_reg_e_cry_23_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[23]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(23), D => \R3_data[23]\, FCI => next_reg_e_cry_22, 
        S => \next_reg_e[23]\, Y => OPEN, FCO => 
        next_reg_e_cry_23);
    
    \reg_h[30]\ : SLE
      port map(D => \next_reg_h[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[30]\);
    
    \next_reg_d[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[6]\, B => N3_data(6), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[6]_net_1\);
    
    \reg_g[10]\ : SLE
      port map(D => \next_reg_g[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[10]\);
    
    \reg_e[2]\ : SLE
      port map(D => \next_reg_e[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[2]\);
    
    \reg_c[20]\ : SLE
      port map(D => \next_reg_c[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[20]\);
    
    \next_reg_b[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(19), B => \R0_data[19]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[19]_net_1\);
    
    \reg_b[23]\ : SLE
      port map(D => \next_reg_b[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[23]\);
    
    \next_reg_f[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(30), B => \R4_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[30]_net_1\);
    
    \reg_g[22]\ : SLE
      port map(D => \next_reg_g[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[22]\);
    
    \reg_c[8]\ : SLE
      port map(D => \next_reg_c[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[8]\);
    
    \reg_b[15]\ : SLE
      port map(D => \next_reg_b[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[15]\);
    
    \reg_g[21]\ : SLE
      port map(D => \next_reg_g[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[21]\);
    
    \reg_h[7]\ : SLE
      port map(D => \next_reg_h[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[7]\);
    
    next_reg_a_cry_20_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[20]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[20]\, D => N0_data(20), FCI => next_reg_a_cry_19, S
         => \next_reg_a[20]\, Y => OPEN, FCO => next_reg_a_cry_20);
    
    sum0_4_cry_0_998 : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[18]\, C => 
        \R0_data[7]\, Y => \SIG0_0[5]\);
    
    sum3_cry_25 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[25]\, B => Wt_data(25), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_24\, S => 
        \sum3[25]\, Y => OPEN, FCO => \sum3_cry_25\);
    
    \next_reg_g[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R5_data[4]\, B => N6_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[4]_net_1\);
    
    sum3_4_cry_29 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[29]\, B => m304, C => i3_mux_1, D => 
        Kt_addr(5), FCI => \sum3_4_cry_28\, S => \sum3_4[29]\, Y
         => OPEN, FCO => \sum3_4_cry_29\);
    
    sum3_6_cry_23 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[23]\, B => \R4_data[2]\, C => 
        \R4_data[16]\, D => \R4_data[29]\, FCI => \sum3_6_cry_22\, 
        S => \sum3_6[23]\, Y => OPEN, FCO => \sum3_6_cry_23\);
    
    \next_reg_g[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(22), B => \R5_data[22]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[22]_net_1\);
    
    \next_reg_b[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N1_data(24), B => \R0_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_b[24]_net_1\);
    
    \reg_e[3]\ : SLE
      port map(D => \next_reg_e[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[3]\);
    
    \SIG0[5]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[27]\, B => \R0_data[18]\, C => 
        \R0_data[7]\, Y => \SIG0[5]_net_1\);
    
    \next_reg_g[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(17), B => \R5_data[17]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[17]_net_1\);
    
    \next_reg_g[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N6_data(15), B => \R5_data[15]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_g[15]_net_1\);
    
    sum3_6_0_cry_7 : ARI1
      generic map(INIT => x"527D8")

      port map(A => \R7_data[7]\, B => \R4_data[7]\, C => 
        \R5_data[7]\, D => \R6_data[7]\, FCI => \sum3_6_0_cry_6\, 
        S => \sum3_6_0[7]\, Y => OPEN, FCO => \sum3_6_0_cry_7\);
    
    sum3_4_cry_26 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[26]\, B => m281_ns, C => m285, D => 
        Kt_addr(5), FCI => \sum3_4_cry_25\, S => \sum3_4[26]\, Y
         => OPEN, FCO => \sum3_4_cry_26\);
    
    \next_reg_f[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(24), B => \R4_data[24]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[24]_net_1\);
    
    \reg_f[6]\ : SLE
      port map(D => \next_reg_f[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[6]\);
    
    sum3_axb_0 : CFG2
      generic map(INIT => x"6")

      port map(A => Wt_data(0), B => sum3_4_cry_0_Y, Y => 
        \sum3[0]\);
    
    \next_reg_h[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(30), B => \R6_data[30]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[30]_net_1\);
    
    sum3_6_cry_28 : ARI1
      generic map(INIT => x"56996")

      port map(A => \sum3_6_0[28]\, B => \R4_data[2]\, C => 
        \R4_data[7]\, D => \R4_data[21]\, FCI => \sum3_6_cry_27\, 
        S => \sum3_6[28]\, Y => OPEN, FCO => \sum3_6_cry_28\);
    
    \reg_a[9]\ : SLE
      port map(D => \next_reg_a[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[9]\);
    
    \SIG0[3]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[25]\, B => \R0_data[16]\, C => 
        \R0_data[5]\, Y => \SIG0[3]_net_1\);
    
    \reg_c[17]\ : SLE
      port map(D => \next_reg_c[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[17]\);
    
    \reg_b[24]\ : SLE
      port map(D => \next_reg_b[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[24]\);
    
    sum0_4_axb_1 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[1]\, B => \R1_data[1]\, C => 
        \R0_data[1]\, D => \SIG0[1]_net_1\, Y => \sum0_4_axb_1\);
    
    \reg_g[26]\ : SLE
      port map(D => \next_reg_g[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[26]\);
    
    \reg_a[6]\ : SLE
      port map(D => \next_reg_a[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[6]\);
    
    \SIG0[22]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[24]\, B => \R0_data[3]\, C => 
        \R0_data[12]\, Y => \SIG0[22]_net_1\);
    
    \reg_d[19]\ : SLE
      port map(D => \next_reg_d[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[19]\);
    
    \reg_d[5]\ : SLE
      port map(D => \next_reg_d[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R3_data[5]\);
    
    \reg_a[4]\ : SLE
      port map(D => \next_reg_a[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[4]\);
    
    \reg_f[20]\ : SLE
      port map(D => \next_reg_f[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[20]\);
    
    next_reg_a_cry_10_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[10]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[10]\, D => N0_data(10), FCI => next_reg_a_cry_9, S
         => \next_reg_a[10]\, Y => OPEN, FCO => next_reg_a_cry_10);
    
    \next_reg_h[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(27), B => \R6_data[27]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[27]_net_1\);
    
    next_reg_e_cry_30_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[30]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(30), D => \R3_data[30]\, FCI => next_reg_e_cry_29, 
        S => \next_reg_e[30]\, Y => OPEN, FCO => 
        next_reg_e_cry_30);
    
    \reg_c[0]\ : SLE
      port map(D => \next_reg_c[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R2_data[0]\);
    
    \next_reg_h[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N7_data(25), B => \R6_data[25]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_h[25]_net_1\);
    
    \next_reg_d[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R2_data[4]\, B => N3_data(4), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_d[4]_net_1\);
    
    \next_reg_f[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(10), B => \R4_data[10]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[10]_net_1\);
    
    \reg_g[7]\ : SLE
      port map(D => \next_reg_g[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[7]\);
    
    sum0_4_axb_14 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[14]\, B => \R1_data[14]\, C => 
        \R0_data[14]\, D => \SIG0[14]_net_1\, Y => 
        \sum0_4_axb_14\);
    
    sum3_cry_13 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum3_4[13]\, B => Wt_data(13), C => 
        GND_net_1, D => GND_net_1, FCI => \sum3_cry_12\, S => 
        \sum3[13]\, Y => OPEN, FCO => \sum3_cry_13\);
    
    \reg_e[13]\ : SLE
      port map(D => \next_reg_e[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R4_data[13]\);
    
    next_reg_a_cry_9_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[9]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[9]\, D => N0_data(9), FCI => next_reg_a_cry_8, S
         => \next_reg_a[9]\, Y => OPEN, FCO => next_reg_a_cry_9);
    
    next_reg_a_cry_30_0 : ARI1
      generic map(INIT => x"572D8")

      port map(A => \sum0_4[30]\, B => oregs_ce_i_a2_0_a2, C => 
        \sum3[30]\, D => N0_data(30), FCI => next_reg_a_cry_29, S
         => \next_reg_a[30]\, Y => OPEN, FCO => next_reg_a_cry_30);
    
    sum3_4_axb_0 : CFG4
      generic map(INIT => x"3AC5")

      port map(A => m10_ns, B => m19, C => Kt_addr(5), D => 
        sum3_6_cry_0_Y, Y => \sum3_4[0]\);
    
    \reg_g[28]\ : SLE
      port map(D => \next_reg_g[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R6_data[28]\);
    
    next_reg_e_cry_16_0 : ARI1
      generic map(INIT => x"54EE4")

      port map(A => \sum3[16]\, B => oregs_ce_i_a2_0_a2, C => 
        N4_data(16), D => \R3_data[16]\, FCI => next_reg_e_cry_15, 
        S => \next_reg_e[16]\, Y => OPEN, FCO => 
        next_reg_e_cry_16);
    
    \reg_h[5]\ : SLE
      port map(D => \next_reg_h[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R7_data[5]\);
    
    \next_reg_f[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \R4_data[5]\, B => N5_data(5), C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[5]_net_1\);
    
    sum3_4_cry_22 : ARI1
      generic map(INIT => x"5CA35")

      port map(A => \sum3_6[22]\, B => m250_am, C => m250_bm, D
         => Kt_addr(5), FCI => \sum3_4_cry_21\, S => \sum3_4[22]\, 
        Y => OPEN, FCO => \sum3_4_cry_22\);
    
    \SIG0[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \R0_data[13]\, B => \R0_data[1]\, C => 
        \R0_data[24]\, Y => \SIG0[11]_net_1\);
    
    \reg_f[31]\ : SLE
      port map(D => \next_reg_f[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R5_data[31]\);
    
    \next_reg_c[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N2_data(29), B => \R1_data[29]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_c[29]_net_1\);
    
    \reg_b[10]\ : SLE
      port map(D => \next_reg_b[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R1_data[10]\);
    
    \reg_a[1]\ : SLE
      port map(D => \next_reg_a[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        core_ce_o_iv_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R0_data[1]\);
    
    sum0_4_axb_17 : CFG4
      generic map(INIT => x"17E8")

      port map(A => \R2_data[17]\, B => \R1_data[17]\, C => 
        \R0_data[17]\, D => \SIG0[17]_net_1\, Y => 
        \sum0_4_axb_17\);
    
    sum3_4_cry_3 : ARI1
      generic map(INIT => x"535CA")

      port map(A => \sum3_6[3]\, B => m62_am, C => m62_bm, D => 
        Kt_addr(5), FCI => \sum3_4_cry_2\, S => \sum3_4[3]\, Y
         => OPEN, FCO => \sum3_4_cry_3\);
    
    \next_reg_f[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N5_data(12), B => \R4_data[12]\, C => 
        oregs_ce_i_a2_0_a2, Y => \next_reg_f[12]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_regs is

    port( SHA256_BLOCK_0_H0_o                  : out   std_logic_vector(31 downto 0);
          N0_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H1_o                  : out   std_logic_vector(31 downto 0);
          N1_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H2_o                  : out   std_logic_vector(31 downto 0);
          N2_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H3_o                  : out   std_logic_vector(31 downto 0);
          N3_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H4_o                  : out   std_logic_vector(31 downto 0);
          N4_data                              : out   std_logic_vector(31 downto 1);
          N5_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H5_o                  : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o                  : out   std_logic_vector(31 downto 0);
          N6_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H7_o                  : out   std_logic_vector(31 downto 0);
          N7_data                              : out   std_logic_vector(31 downto 1);
          hash_control_st_reg_i                : in    std_logic_vector(6 to 6);
          R0_data                              : in    std_logic_vector(31 downto 0);
          R1_data                              : in    std_logic_vector(31 downto 0);
          R2_data                              : in    std_logic_vector(31 downto 0);
          R3_data                              : in    std_logic_vector(31 downto 0);
          R4_data                              : in    std_logic_vector(31 downto 0);
          R5_data                              : in    std_logic_vector(31 downto 0);
          R6_data                              : in    std_logic_vector(31 downto 0);
          R7_data                              : in    std_logic_vector(31 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          N_168_i_0                            : in    std_logic;
          next_reg_H0_cry_0_0_Y                : out   std_logic;
          next_reg_H1_cry_0_0_Y                : out   std_logic;
          next_reg_H2_cry_0_0_Y                : out   std_logic;
          next_reg_H3_cry_0_0_Y                : out   std_logic;
          next_reg_H4_cry_0_0_Y                : out   std_logic;
          next_reg_H5_cry_0_0_Y                : out   std_logic;
          next_reg_H6_cry_0_0_Y                : out   std_logic;
          next_reg_H7_cry_0_0_Y                : out   std_logic
        );

end sha256_regs;

architecture DEF_ARCH of sha256_regs is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \SHA256_BLOCK_0_H0_o[21]\, VCC_net_1, \N0_data[21]\, 
        GND_net_1, \SHA256_BLOCK_0_H0_o[22]\, \N0_data[22]\, 
        \SHA256_BLOCK_0_H0_o[23]\, \N0_data[23]\, 
        \SHA256_BLOCK_0_H0_o[24]\, \N0_data[24]\, 
        \SHA256_BLOCK_0_H0_o[25]\, \N0_data[25]\, 
        \SHA256_BLOCK_0_H0_o[26]\, \N0_data[26]\, 
        \SHA256_BLOCK_0_H0_o[27]\, \N0_data[27]\, 
        \SHA256_BLOCK_0_H0_o[28]\, \N0_data[28]\, 
        \SHA256_BLOCK_0_H0_o[29]\, \N0_data[29]\, 
        \SHA256_BLOCK_0_H0_o[30]\, \N0_data[30]\, 
        \SHA256_BLOCK_0_H0_o[31]\, \N0_data[31]\, 
        \SHA256_BLOCK_0_H0_o[6]\, \N0_data[6]\, 
        \SHA256_BLOCK_0_H0_o[7]\, \N0_data[7]\, 
        \SHA256_BLOCK_0_H0_o[8]\, \N0_data[8]\, 
        \SHA256_BLOCK_0_H0_o[9]\, \N0_data[9]\, 
        \SHA256_BLOCK_0_H0_o[10]\, \N0_data[10]\, 
        \SHA256_BLOCK_0_H0_o[11]\, \N0_data[11]\, 
        \SHA256_BLOCK_0_H0_o[12]\, \N0_data[12]\, 
        \SHA256_BLOCK_0_H0_o[13]\, \N0_data[13]\, 
        \SHA256_BLOCK_0_H0_o[14]\, \N0_data[14]\, 
        \SHA256_BLOCK_0_H0_o[15]\, \N0_data[15]\, 
        \SHA256_BLOCK_0_H0_o[16]\, \N0_data[16]\, 
        \SHA256_BLOCK_0_H0_o[17]\, \N0_data[17]\, 
        \SHA256_BLOCK_0_H0_o[18]\, \N0_data[18]\, 
        \SHA256_BLOCK_0_H0_o[19]\, \N0_data[19]\, 
        \SHA256_BLOCK_0_H0_o[20]\, \N0_data[20]\, 
        \SHA256_BLOCK_0_H1_o[23]\, \N1_data[23]\, 
        \SHA256_BLOCK_0_H1_o[24]\, \N1_data[24]\, 
        \SHA256_BLOCK_0_H1_o[25]\, \N1_data[25]\, 
        \SHA256_BLOCK_0_H1_o[26]\, \N1_data[26]\, 
        \SHA256_BLOCK_0_H1_o[27]\, \N1_data[27]\, 
        \SHA256_BLOCK_0_H1_o[28]\, \N1_data[28]\, 
        \SHA256_BLOCK_0_H1_o[29]\, \N1_data[29]\, 
        \SHA256_BLOCK_0_H1_o[30]\, \N1_data[30]\, 
        \SHA256_BLOCK_0_H1_o[31]\, \N1_data[31]\, 
        \SHA256_BLOCK_0_H0_o[0]\, \next_reg_H0_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H0_o[1]\, \N0_data[1]\, 
        \SHA256_BLOCK_0_H0_o[2]\, \N0_data[2]\, 
        \SHA256_BLOCK_0_H0_o[3]\, \N0_data[3]\, 
        \SHA256_BLOCK_0_H0_o[4]\, \N0_data[4]\, 
        \SHA256_BLOCK_0_H0_o[5]\, \N0_data[5]\, 
        \SHA256_BLOCK_0_H1_o[8]\, \N1_data[8]\, 
        \SHA256_BLOCK_0_H1_o[9]\, \N1_data[9]\, 
        \SHA256_BLOCK_0_H1_o[10]\, \N1_data[10]\, 
        \SHA256_BLOCK_0_H1_o[11]\, \N1_data[11]\, 
        \SHA256_BLOCK_0_H1_o[12]\, \N1_data[12]\, 
        \SHA256_BLOCK_0_H1_o[13]\, \N1_data[13]\, 
        \SHA256_BLOCK_0_H1_o[14]\, \N1_data[14]\, 
        \SHA256_BLOCK_0_H1_o[15]\, \N1_data[15]\, 
        \SHA256_BLOCK_0_H1_o[16]\, \N1_data[16]\, 
        \SHA256_BLOCK_0_H1_o[17]\, \N1_data[17]\, 
        \SHA256_BLOCK_0_H1_o[18]\, \N1_data[18]\, 
        \SHA256_BLOCK_0_H1_o[19]\, \N1_data[19]\, 
        \SHA256_BLOCK_0_H1_o[20]\, \N1_data[20]\, 
        \SHA256_BLOCK_0_H1_o[21]\, \N1_data[21]\, 
        \SHA256_BLOCK_0_H1_o[22]\, \N1_data[22]\, 
        \SHA256_BLOCK_0_H2_o[25]\, \N2_data[25]\, 
        \SHA256_BLOCK_0_H2_o[26]\, \N2_data[26]\, 
        \SHA256_BLOCK_0_H2_o[27]\, \N2_data[27]\, 
        \SHA256_BLOCK_0_H2_o[28]\, \N2_data[28]\, 
        \SHA256_BLOCK_0_H2_o[29]\, \N2_data[29]\, 
        \SHA256_BLOCK_0_H2_o[30]\, \N2_data[30]\, 
        \SHA256_BLOCK_0_H2_o[31]\, \N2_data[31]\, 
        \SHA256_BLOCK_0_H1_o[0]\, \next_reg_H1_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H1_o[1]\, \N1_data[1]\, 
        \SHA256_BLOCK_0_H1_o[2]\, \N1_data[2]\, 
        \SHA256_BLOCK_0_H1_o[3]\, \N1_data[3]\, 
        \SHA256_BLOCK_0_H1_o[4]\, \N1_data[4]\, 
        \SHA256_BLOCK_0_H1_o[5]\, \N1_data[5]\, 
        \SHA256_BLOCK_0_H1_o[6]\, \N1_data[6]\, 
        \SHA256_BLOCK_0_H1_o[7]\, \N1_data[7]\, 
        \SHA256_BLOCK_0_H2_o[10]\, \N2_data[10]\, 
        \SHA256_BLOCK_0_H2_o[11]\, \N2_data[11]\, 
        \SHA256_BLOCK_0_H2_o[12]\, \N2_data[12]\, 
        \SHA256_BLOCK_0_H2_o[13]\, \N2_data[13]\, 
        \SHA256_BLOCK_0_H2_o[14]\, \N2_data[14]\, 
        \SHA256_BLOCK_0_H2_o[15]\, \N2_data[15]\, 
        \SHA256_BLOCK_0_H2_o[16]\, \N2_data[16]\, 
        \SHA256_BLOCK_0_H2_o[17]\, \N2_data[17]\, 
        \SHA256_BLOCK_0_H2_o[18]\, \N2_data[18]\, 
        \SHA256_BLOCK_0_H2_o[19]\, \N2_data[19]\, 
        \SHA256_BLOCK_0_H2_o[20]\, \N2_data[20]\, 
        \SHA256_BLOCK_0_H2_o[21]\, \N2_data[21]\, 
        \SHA256_BLOCK_0_H2_o[22]\, \N2_data[22]\, 
        \SHA256_BLOCK_0_H2_o[23]\, \N2_data[23]\, 
        \SHA256_BLOCK_0_H2_o[24]\, \N2_data[24]\, 
        \SHA256_BLOCK_0_H3_o[27]\, \N3_data[27]\, 
        \SHA256_BLOCK_0_H3_o[28]\, \N3_data[28]\, 
        \SHA256_BLOCK_0_H3_o[29]\, \N3_data[29]\, 
        \SHA256_BLOCK_0_H3_o[30]\, \N3_data[30]\, 
        \SHA256_BLOCK_0_H3_o[31]\, \N3_data[31]\, 
        \SHA256_BLOCK_0_H2_o[0]\, \next_reg_H2_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H2_o[1]\, \N2_data[1]\, 
        \SHA256_BLOCK_0_H2_o[2]\, \N2_data[2]\, 
        \SHA256_BLOCK_0_H2_o[3]\, \N2_data[3]\, 
        \SHA256_BLOCK_0_H2_o[4]\, \N2_data[4]\, 
        \SHA256_BLOCK_0_H2_o[5]\, \N2_data[5]\, 
        \SHA256_BLOCK_0_H2_o[6]\, \N2_data[6]\, 
        \SHA256_BLOCK_0_H2_o[7]\, \N2_data[7]\, 
        \SHA256_BLOCK_0_H2_o[8]\, \N2_data[8]\, 
        \SHA256_BLOCK_0_H2_o[9]\, \N2_data[9]\, 
        \SHA256_BLOCK_0_H3_o[12]\, \N3_data[12]\, 
        \SHA256_BLOCK_0_H3_o[13]\, \N3_data[13]\, 
        \SHA256_BLOCK_0_H3_o[14]\, \N3_data[14]\, 
        \SHA256_BLOCK_0_H3_o[15]\, \N3_data[15]\, 
        \SHA256_BLOCK_0_H3_o[16]\, \N3_data[16]\, 
        \SHA256_BLOCK_0_H3_o[17]\, \N3_data[17]\, 
        \SHA256_BLOCK_0_H3_o[18]\, \N3_data[18]\, 
        \SHA256_BLOCK_0_H3_o[19]\, \N3_data[19]\, 
        \SHA256_BLOCK_0_H3_o[20]\, \N3_data[20]\, 
        \SHA256_BLOCK_0_H3_o[21]\, \N3_data[21]\, 
        \SHA256_BLOCK_0_H3_o[22]\, \N3_data[22]\, 
        \SHA256_BLOCK_0_H3_o[23]\, \N3_data[23]\, 
        \SHA256_BLOCK_0_H3_o[24]\, \N3_data[24]\, 
        \SHA256_BLOCK_0_H3_o[25]\, \N3_data[25]\, 
        \SHA256_BLOCK_0_H3_o[26]\, \N3_data[26]\, 
        \SHA256_BLOCK_0_H4_o[29]\, \N4_data[29]\, 
        \SHA256_BLOCK_0_H4_o[30]\, \N4_data[30]\, 
        \SHA256_BLOCK_0_H4_o[31]\, \N4_data[31]\, 
        \SHA256_BLOCK_0_H3_o[0]\, \next_reg_H3_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H3_o[1]\, \N3_data[1]\, 
        \SHA256_BLOCK_0_H3_o[2]\, \N3_data[2]\, 
        \SHA256_BLOCK_0_H3_o[3]\, \N3_data[3]\, 
        \SHA256_BLOCK_0_H3_o[4]\, \N3_data[4]\, 
        \SHA256_BLOCK_0_H3_o[5]\, \N3_data[5]\, 
        \SHA256_BLOCK_0_H3_o[6]\, \N3_data[6]\, 
        \SHA256_BLOCK_0_H3_o[7]\, \N3_data[7]\, 
        \SHA256_BLOCK_0_H3_o[8]\, \N3_data[8]\, 
        \SHA256_BLOCK_0_H3_o[9]\, \N3_data[9]\, 
        \SHA256_BLOCK_0_H3_o[10]\, \N3_data[10]\, 
        \SHA256_BLOCK_0_H3_o[11]\, \N3_data[11]\, 
        \SHA256_BLOCK_0_H4_o[14]\, \N4_data[14]\, 
        \SHA256_BLOCK_0_H4_o[15]\, \N4_data[15]\, 
        \SHA256_BLOCK_0_H4_o[16]\, \N4_data[16]\, 
        \SHA256_BLOCK_0_H4_o[17]\, \N4_data[17]\, 
        \SHA256_BLOCK_0_H4_o[18]\, \N4_data[18]\, 
        \SHA256_BLOCK_0_H4_o[19]\, \N4_data[19]\, 
        \SHA256_BLOCK_0_H4_o[20]\, \N4_data[20]\, 
        \SHA256_BLOCK_0_H4_o[21]\, \N4_data[21]\, 
        \SHA256_BLOCK_0_H4_o[22]\, \N4_data[22]\, 
        \SHA256_BLOCK_0_H4_o[23]\, \N4_data[23]\, 
        \SHA256_BLOCK_0_H4_o[24]\, \N4_data[24]\, 
        \SHA256_BLOCK_0_H4_o[25]\, \N4_data[25]\, 
        \SHA256_BLOCK_0_H4_o[26]\, \N4_data[26]\, 
        \SHA256_BLOCK_0_H4_o[27]\, \N4_data[27]\, 
        \SHA256_BLOCK_0_H4_o[28]\, \N4_data[28]\, 
        \SHA256_BLOCK_0_H5_o[31]\, \N5_data[31]\, 
        \SHA256_BLOCK_0_H4_o[0]\, \next_reg_H4_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H4_o[1]\, \N4_data[1]\, 
        \SHA256_BLOCK_0_H4_o[2]\, \N4_data[2]\, 
        \SHA256_BLOCK_0_H4_o[3]\, \N4_data[3]\, 
        \SHA256_BLOCK_0_H4_o[4]\, \N4_data[4]\, 
        \SHA256_BLOCK_0_H4_o[5]\, \N4_data[5]\, 
        \SHA256_BLOCK_0_H4_o[6]\, \N4_data[6]\, 
        \SHA256_BLOCK_0_H4_o[7]\, \N4_data[7]\, 
        \SHA256_BLOCK_0_H4_o[8]\, \N4_data[8]\, 
        \SHA256_BLOCK_0_H4_o[9]\, \N4_data[9]\, 
        \SHA256_BLOCK_0_H4_o[10]\, \N4_data[10]\, 
        \SHA256_BLOCK_0_H4_o[11]\, \N4_data[11]\, 
        \SHA256_BLOCK_0_H4_o[12]\, \N4_data[12]\, 
        \SHA256_BLOCK_0_H4_o[13]\, \N4_data[13]\, 
        \SHA256_BLOCK_0_H5_o[16]\, \N5_data[16]\, 
        \SHA256_BLOCK_0_H5_o[17]\, \N5_data[17]\, 
        \SHA256_BLOCK_0_H5_o[18]\, \N5_data[18]\, 
        \SHA256_BLOCK_0_H5_o[19]\, \N5_data[19]\, 
        \SHA256_BLOCK_0_H5_o[20]\, \N5_data[20]\, 
        \SHA256_BLOCK_0_H5_o[21]\, \N5_data[21]\, 
        \SHA256_BLOCK_0_H5_o[22]\, \N5_data[22]\, 
        \SHA256_BLOCK_0_H5_o[23]\, \N5_data[23]\, 
        \SHA256_BLOCK_0_H5_o[24]\, \N5_data[24]\, 
        \SHA256_BLOCK_0_H5_o[25]\, \N5_data[25]\, 
        \SHA256_BLOCK_0_H5_o[26]\, \N5_data[26]\, 
        \SHA256_BLOCK_0_H5_o[27]\, \N5_data[27]\, 
        \SHA256_BLOCK_0_H5_o[28]\, \N5_data[28]\, 
        \SHA256_BLOCK_0_H5_o[29]\, \N5_data[29]\, 
        \SHA256_BLOCK_0_H5_o[30]\, \N5_data[30]\, 
        \SHA256_BLOCK_0_H5_o[1]\, \N5_data[1]\, 
        \SHA256_BLOCK_0_H5_o[2]\, \N5_data[2]\, 
        \SHA256_BLOCK_0_H5_o[3]\, \N5_data[3]\, 
        \SHA256_BLOCK_0_H5_o[4]\, \N5_data[4]\, 
        \SHA256_BLOCK_0_H5_o[5]\, \N5_data[5]\, 
        \SHA256_BLOCK_0_H5_o[6]\, \N5_data[6]\, 
        \SHA256_BLOCK_0_H5_o[7]\, \N5_data[7]\, 
        \SHA256_BLOCK_0_H5_o[8]\, \N5_data[8]\, 
        \SHA256_BLOCK_0_H5_o[9]\, \N5_data[9]\, 
        \SHA256_BLOCK_0_H5_o[10]\, \N5_data[10]\, 
        \SHA256_BLOCK_0_H5_o[11]\, \N5_data[11]\, 
        \SHA256_BLOCK_0_H5_o[12]\, \N5_data[12]\, 
        \SHA256_BLOCK_0_H5_o[13]\, \N5_data[13]\, 
        \SHA256_BLOCK_0_H5_o[14]\, \N5_data[14]\, 
        \SHA256_BLOCK_0_H5_o[15]\, \N5_data[15]\, 
        \SHA256_BLOCK_0_H6_o[18]\, \N6_data[18]\, 
        \SHA256_BLOCK_0_H6_o[19]\, \N6_data[19]\, 
        \SHA256_BLOCK_0_H6_o[20]\, \N6_data[20]\, 
        \SHA256_BLOCK_0_H6_o[21]\, \N6_data[21]\, 
        \SHA256_BLOCK_0_H6_o[22]\, \N6_data[22]\, 
        \SHA256_BLOCK_0_H6_o[23]\, \N6_data[23]\, 
        \SHA256_BLOCK_0_H6_o[24]\, \N6_data[24]\, 
        \SHA256_BLOCK_0_H6_o[25]\, \N6_data[25]\, 
        \SHA256_BLOCK_0_H6_o[26]\, \N6_data[26]\, 
        \SHA256_BLOCK_0_H6_o[27]\, \N6_data[27]\, 
        \SHA256_BLOCK_0_H6_o[28]\, \N6_data[28]\, 
        \SHA256_BLOCK_0_H6_o[29]\, \N6_data[29]\, 
        \SHA256_BLOCK_0_H6_o[30]\, \N6_data[30]\, 
        \SHA256_BLOCK_0_H6_o[31]\, \N6_data[31]\, 
        \SHA256_BLOCK_0_H5_o[0]\, \next_reg_H5_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H6_o[3]\, \N6_data[3]\, 
        \SHA256_BLOCK_0_H6_o[4]\, \N6_data[4]\, 
        \SHA256_BLOCK_0_H6_o[5]\, \N6_data[5]\, 
        \SHA256_BLOCK_0_H6_o[6]\, \N6_data[6]\, 
        \SHA256_BLOCK_0_H6_o[7]\, \N6_data[7]\, 
        \SHA256_BLOCK_0_H6_o[8]\, \N6_data[8]\, 
        \SHA256_BLOCK_0_H6_o[9]\, \N6_data[9]\, 
        \SHA256_BLOCK_0_H6_o[10]\, \N6_data[10]\, 
        \SHA256_BLOCK_0_H6_o[11]\, \N6_data[11]\, 
        \SHA256_BLOCK_0_H6_o[12]\, \N6_data[12]\, 
        \SHA256_BLOCK_0_H6_o[13]\, \N6_data[13]\, 
        \SHA256_BLOCK_0_H6_o[14]\, \N6_data[14]\, 
        \SHA256_BLOCK_0_H6_o[15]\, \N6_data[15]\, 
        \SHA256_BLOCK_0_H6_o[16]\, \N6_data[16]\, 
        \SHA256_BLOCK_0_H6_o[17]\, \N6_data[17]\, 
        \SHA256_BLOCK_0_H7_o[20]\, \N7_data[20]\, 
        \SHA256_BLOCK_0_H7_o[21]\, \N7_data[21]\, 
        \SHA256_BLOCK_0_H7_o[22]\, \N7_data[22]\, 
        \SHA256_BLOCK_0_H7_o[23]\, \N7_data[23]\, 
        \SHA256_BLOCK_0_H7_o[24]\, \N7_data[24]\, 
        \SHA256_BLOCK_0_H7_o[25]\, \N7_data[25]\, 
        \SHA256_BLOCK_0_H7_o[26]\, \N7_data[26]\, 
        \SHA256_BLOCK_0_H7_o[27]\, \N7_data[27]\, 
        \SHA256_BLOCK_0_H7_o[28]\, \N7_data[28]\, 
        \SHA256_BLOCK_0_H7_o[29]\, \N7_data[29]\, 
        \SHA256_BLOCK_0_H7_o[30]\, \N7_data[30]\, 
        \SHA256_BLOCK_0_H7_o[31]\, \N7_data[31]\, 
        \SHA256_BLOCK_0_H6_o[0]\, \next_reg_H6_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H6_o[1]\, \N6_data[1]\, 
        \SHA256_BLOCK_0_H6_o[2]\, \N6_data[2]\, 
        \SHA256_BLOCK_0_H7_o[5]\, \N7_data[5]\, 
        \SHA256_BLOCK_0_H7_o[6]\, \N7_data[6]\, 
        \SHA256_BLOCK_0_H7_o[7]\, \N7_data[7]\, 
        \SHA256_BLOCK_0_H7_o[8]\, \N7_data[8]\, 
        \SHA256_BLOCK_0_H7_o[9]\, \N7_data[9]\, 
        \SHA256_BLOCK_0_H7_o[10]\, \N7_data[10]\, 
        \SHA256_BLOCK_0_H7_o[11]\, \N7_data[11]\, 
        \SHA256_BLOCK_0_H7_o[12]\, \N7_data[12]\, 
        \SHA256_BLOCK_0_H7_o[13]\, \N7_data[13]\, 
        \SHA256_BLOCK_0_H7_o[14]\, \N7_data[14]\, 
        \SHA256_BLOCK_0_H7_o[15]\, \N7_data[15]\, 
        \SHA256_BLOCK_0_H7_o[16]\, \N7_data[16]\, 
        \SHA256_BLOCK_0_H7_o[17]\, \N7_data[17]\, 
        \SHA256_BLOCK_0_H7_o[18]\, \N7_data[18]\, 
        \SHA256_BLOCK_0_H7_o[19]\, \N7_data[19]\, 
        \SHA256_BLOCK_0_H7_o[0]\, \next_reg_H7_cry_0_0_Y\, 
        \SHA256_BLOCK_0_H7_o[1]\, \N7_data[1]\, 
        \SHA256_BLOCK_0_H7_o[2]\, \N7_data[2]\, 
        \SHA256_BLOCK_0_H7_o[3]\, \N7_data[3]\, 
        \SHA256_BLOCK_0_H7_o[4]\, \N7_data[4]\, next_reg_H0_cry_0, 
        next_reg_H0_cry_1, next_reg_H0_cry_2, next_reg_H0_cry_3, 
        next_reg_H0_cry_4, next_reg_H0_cry_5, next_reg_H0_cry_6, 
        next_reg_H0_cry_7, next_reg_H0_cry_8, next_reg_H0_cry_9, 
        next_reg_H0_cry_10, next_reg_H0_cry_11, 
        next_reg_H0_cry_12, next_reg_H0_cry_13, 
        next_reg_H0_cry_14, next_reg_H0_cry_15, 
        next_reg_H0_cry_16, next_reg_H0_cry_17, 
        next_reg_H0_cry_18, next_reg_H0_cry_19, 
        next_reg_H0_cry_20, next_reg_H0_cry_21, 
        next_reg_H0_cry_22, next_reg_H0_cry_23, 
        next_reg_H0_cry_24, next_reg_H0_cry_25, 
        next_reg_H0_cry_26, next_reg_H0_cry_27, 
        next_reg_H0_cry_28, next_reg_H0_cry_29, 
        next_reg_H0_cry_30, next_reg_H1_cry_0, next_reg_H1_cry_1, 
        next_reg_H1_cry_2, next_reg_H1_cry_3, next_reg_H1_cry_4, 
        next_reg_H1_cry_5, next_reg_H1_cry_6, next_reg_H1_cry_7, 
        next_reg_H1_cry_8, next_reg_H1_cry_9, next_reg_H1_cry_10, 
        next_reg_H1_cry_11, next_reg_H1_cry_12, 
        next_reg_H1_cry_13, next_reg_H1_cry_14, 
        next_reg_H1_cry_15, next_reg_H1_cry_16, 
        next_reg_H1_cry_17, next_reg_H1_cry_18, 
        next_reg_H1_cry_19, next_reg_H1_cry_20, 
        next_reg_H1_cry_21, next_reg_H1_cry_22, 
        next_reg_H1_cry_23, next_reg_H1_cry_24, 
        next_reg_H1_cry_25, next_reg_H1_cry_26, 
        next_reg_H1_cry_27, next_reg_H1_cry_28, 
        next_reg_H1_cry_29, next_reg_H1_cry_30, next_reg_H2_cry_0, 
        next_reg_H2_cry_1, next_reg_H2_cry_2, next_reg_H2_cry_3, 
        next_reg_H2_cry_4, next_reg_H2_cry_5, next_reg_H2_cry_6, 
        next_reg_H2_cry_7, next_reg_H2_cry_8, next_reg_H2_cry_9, 
        next_reg_H2_cry_10, next_reg_H2_cry_11, 
        next_reg_H2_cry_12, next_reg_H2_cry_13, 
        next_reg_H2_cry_14, next_reg_H2_cry_15, 
        next_reg_H2_cry_16, next_reg_H2_cry_17, 
        next_reg_H2_cry_18, next_reg_H2_cry_19, 
        next_reg_H2_cry_20, next_reg_H2_cry_21, 
        next_reg_H2_cry_22, next_reg_H2_cry_23, 
        next_reg_H2_cry_24, next_reg_H2_cry_25, 
        next_reg_H2_cry_26, next_reg_H2_cry_27, 
        next_reg_H2_cry_28, next_reg_H2_cry_29, 
        next_reg_H2_cry_30, next_reg_H3_cry_0, next_reg_H3_cry_1, 
        next_reg_H3_cry_2, next_reg_H3_cry_3, next_reg_H3_cry_4, 
        next_reg_H3_cry_5, next_reg_H3_cry_6, next_reg_H3_cry_7, 
        next_reg_H3_cry_8, next_reg_H3_cry_9, next_reg_H3_cry_10, 
        next_reg_H3_cry_11, next_reg_H3_cry_12, 
        next_reg_H3_cry_13, next_reg_H3_cry_14, 
        next_reg_H3_cry_15, next_reg_H3_cry_16, 
        next_reg_H3_cry_17, next_reg_H3_cry_18, 
        next_reg_H3_cry_19, next_reg_H3_cry_20, 
        next_reg_H3_cry_21, next_reg_H3_cry_22, 
        next_reg_H3_cry_23, next_reg_H3_cry_24, 
        next_reg_H3_cry_25, next_reg_H3_cry_26, 
        next_reg_H3_cry_27, next_reg_H3_cry_28, 
        next_reg_H3_cry_29, next_reg_H3_cry_30, next_reg_H4_cry_0, 
        next_reg_H4_cry_1, next_reg_H4_cry_2, next_reg_H4_cry_3, 
        next_reg_H4_cry_4, next_reg_H4_cry_5, next_reg_H4_cry_6, 
        next_reg_H4_cry_7, next_reg_H4_cry_8, next_reg_H4_cry_9, 
        next_reg_H4_cry_10, next_reg_H4_cry_11, 
        next_reg_H4_cry_12, next_reg_H4_cry_13, 
        next_reg_H4_cry_14, next_reg_H4_cry_15, 
        next_reg_H4_cry_16, next_reg_H4_cry_17, 
        next_reg_H4_cry_18, next_reg_H4_cry_19, 
        next_reg_H4_cry_20, next_reg_H4_cry_21, 
        next_reg_H4_cry_22, next_reg_H4_cry_23, 
        next_reg_H4_cry_24, next_reg_H4_cry_25, 
        next_reg_H4_cry_26, next_reg_H4_cry_27, 
        next_reg_H4_cry_28, next_reg_H4_cry_29, 
        next_reg_H4_cry_30, next_reg_H5_cry_0, next_reg_H5_cry_1, 
        next_reg_H5_cry_2, next_reg_H5_cry_3, next_reg_H5_cry_4, 
        next_reg_H5_cry_5, next_reg_H5_cry_6, next_reg_H5_cry_7, 
        next_reg_H5_cry_8, next_reg_H5_cry_9, next_reg_H5_cry_10, 
        next_reg_H5_cry_11, next_reg_H5_cry_12, 
        next_reg_H5_cry_13, next_reg_H5_cry_14, 
        next_reg_H5_cry_15, next_reg_H5_cry_16, 
        next_reg_H5_cry_17, next_reg_H5_cry_18, 
        next_reg_H5_cry_19, next_reg_H5_cry_20, 
        next_reg_H5_cry_21, next_reg_H5_cry_22, 
        next_reg_H5_cry_23, next_reg_H5_cry_24, 
        next_reg_H5_cry_25, next_reg_H5_cry_26, 
        next_reg_H5_cry_27, next_reg_H5_cry_28, 
        next_reg_H5_cry_29, next_reg_H5_cry_30, next_reg_H6_cry_0, 
        next_reg_H6_cry_1, next_reg_H6_cry_2, next_reg_H6_cry_3, 
        next_reg_H6_cry_4, next_reg_H6_cry_5, next_reg_H6_cry_6, 
        next_reg_H6_cry_7, next_reg_H6_cry_8, next_reg_H6_cry_9, 
        next_reg_H6_cry_10, next_reg_H6_cry_11, 
        next_reg_H6_cry_12, next_reg_H6_cry_13, 
        next_reg_H6_cry_14, next_reg_H6_cry_15, 
        next_reg_H6_cry_16, next_reg_H6_cry_17, 
        next_reg_H6_cry_18, next_reg_H6_cry_19, 
        next_reg_H6_cry_20, next_reg_H6_cry_21, 
        next_reg_H6_cry_22, next_reg_H6_cry_23, 
        next_reg_H6_cry_24, next_reg_H6_cry_25, 
        next_reg_H6_cry_26, next_reg_H6_cry_27, 
        next_reg_H6_cry_28, next_reg_H6_cry_29, 
        next_reg_H6_cry_30, next_reg_H7_cry_0, next_reg_H7_cry_1, 
        next_reg_H7_cry_2, next_reg_H7_cry_3, next_reg_H7_cry_4, 
        next_reg_H7_cry_5, next_reg_H7_cry_6, next_reg_H7_cry_7, 
        next_reg_H7_cry_8, next_reg_H7_cry_9, next_reg_H7_cry_10, 
        next_reg_H7_cry_11, next_reg_H7_cry_12, 
        next_reg_H7_cry_13, next_reg_H7_cry_14, 
        next_reg_H7_cry_15, next_reg_H7_cry_16, 
        next_reg_H7_cry_17, next_reg_H7_cry_18, 
        next_reg_H7_cry_19, next_reg_H7_cry_20, 
        next_reg_H7_cry_21, next_reg_H7_cry_22, 
        next_reg_H7_cry_23, next_reg_H7_cry_24, 
        next_reg_H7_cry_25, next_reg_H7_cry_26, 
        next_reg_H7_cry_27, next_reg_H7_cry_28, 
        next_reg_H7_cry_29, next_reg_H7_cry_30 : std_logic;

begin 

    SHA256_BLOCK_0_H0_o(31) <= \SHA256_BLOCK_0_H0_o[31]\;
    SHA256_BLOCK_0_H0_o(30) <= \SHA256_BLOCK_0_H0_o[30]\;
    SHA256_BLOCK_0_H0_o(29) <= \SHA256_BLOCK_0_H0_o[29]\;
    SHA256_BLOCK_0_H0_o(28) <= \SHA256_BLOCK_0_H0_o[28]\;
    SHA256_BLOCK_0_H0_o(27) <= \SHA256_BLOCK_0_H0_o[27]\;
    SHA256_BLOCK_0_H0_o(26) <= \SHA256_BLOCK_0_H0_o[26]\;
    SHA256_BLOCK_0_H0_o(25) <= \SHA256_BLOCK_0_H0_o[25]\;
    SHA256_BLOCK_0_H0_o(24) <= \SHA256_BLOCK_0_H0_o[24]\;
    SHA256_BLOCK_0_H0_o(23) <= \SHA256_BLOCK_0_H0_o[23]\;
    SHA256_BLOCK_0_H0_o(22) <= \SHA256_BLOCK_0_H0_o[22]\;
    SHA256_BLOCK_0_H0_o(21) <= \SHA256_BLOCK_0_H0_o[21]\;
    SHA256_BLOCK_0_H0_o(20) <= \SHA256_BLOCK_0_H0_o[20]\;
    SHA256_BLOCK_0_H0_o(19) <= \SHA256_BLOCK_0_H0_o[19]\;
    SHA256_BLOCK_0_H0_o(18) <= \SHA256_BLOCK_0_H0_o[18]\;
    SHA256_BLOCK_0_H0_o(17) <= \SHA256_BLOCK_0_H0_o[17]\;
    SHA256_BLOCK_0_H0_o(16) <= \SHA256_BLOCK_0_H0_o[16]\;
    SHA256_BLOCK_0_H0_o(15) <= \SHA256_BLOCK_0_H0_o[15]\;
    SHA256_BLOCK_0_H0_o(14) <= \SHA256_BLOCK_0_H0_o[14]\;
    SHA256_BLOCK_0_H0_o(13) <= \SHA256_BLOCK_0_H0_o[13]\;
    SHA256_BLOCK_0_H0_o(12) <= \SHA256_BLOCK_0_H0_o[12]\;
    SHA256_BLOCK_0_H0_o(11) <= \SHA256_BLOCK_0_H0_o[11]\;
    SHA256_BLOCK_0_H0_o(10) <= \SHA256_BLOCK_0_H0_o[10]\;
    SHA256_BLOCK_0_H0_o(9) <= \SHA256_BLOCK_0_H0_o[9]\;
    SHA256_BLOCK_0_H0_o(8) <= \SHA256_BLOCK_0_H0_o[8]\;
    SHA256_BLOCK_0_H0_o(7) <= \SHA256_BLOCK_0_H0_o[7]\;
    SHA256_BLOCK_0_H0_o(6) <= \SHA256_BLOCK_0_H0_o[6]\;
    SHA256_BLOCK_0_H0_o(5) <= \SHA256_BLOCK_0_H0_o[5]\;
    SHA256_BLOCK_0_H0_o(4) <= \SHA256_BLOCK_0_H0_o[4]\;
    SHA256_BLOCK_0_H0_o(3) <= \SHA256_BLOCK_0_H0_o[3]\;
    SHA256_BLOCK_0_H0_o(2) <= \SHA256_BLOCK_0_H0_o[2]\;
    SHA256_BLOCK_0_H0_o(1) <= \SHA256_BLOCK_0_H0_o[1]\;
    SHA256_BLOCK_0_H0_o(0) <= \SHA256_BLOCK_0_H0_o[0]\;
    N0_data(31) <= \N0_data[31]\;
    N0_data(30) <= \N0_data[30]\;
    N0_data(29) <= \N0_data[29]\;
    N0_data(28) <= \N0_data[28]\;
    N0_data(27) <= \N0_data[27]\;
    N0_data(26) <= \N0_data[26]\;
    N0_data(25) <= \N0_data[25]\;
    N0_data(24) <= \N0_data[24]\;
    N0_data(23) <= \N0_data[23]\;
    N0_data(22) <= \N0_data[22]\;
    N0_data(21) <= \N0_data[21]\;
    N0_data(20) <= \N0_data[20]\;
    N0_data(19) <= \N0_data[19]\;
    N0_data(18) <= \N0_data[18]\;
    N0_data(17) <= \N0_data[17]\;
    N0_data(16) <= \N0_data[16]\;
    N0_data(15) <= \N0_data[15]\;
    N0_data(14) <= \N0_data[14]\;
    N0_data(13) <= \N0_data[13]\;
    N0_data(12) <= \N0_data[12]\;
    N0_data(11) <= \N0_data[11]\;
    N0_data(10) <= \N0_data[10]\;
    N0_data(9) <= \N0_data[9]\;
    N0_data(8) <= \N0_data[8]\;
    N0_data(7) <= \N0_data[7]\;
    N0_data(6) <= \N0_data[6]\;
    N0_data(5) <= \N0_data[5]\;
    N0_data(4) <= \N0_data[4]\;
    N0_data(3) <= \N0_data[3]\;
    N0_data(2) <= \N0_data[2]\;
    N0_data(1) <= \N0_data[1]\;
    SHA256_BLOCK_0_H1_o(31) <= \SHA256_BLOCK_0_H1_o[31]\;
    SHA256_BLOCK_0_H1_o(30) <= \SHA256_BLOCK_0_H1_o[30]\;
    SHA256_BLOCK_0_H1_o(29) <= \SHA256_BLOCK_0_H1_o[29]\;
    SHA256_BLOCK_0_H1_o(28) <= \SHA256_BLOCK_0_H1_o[28]\;
    SHA256_BLOCK_0_H1_o(27) <= \SHA256_BLOCK_0_H1_o[27]\;
    SHA256_BLOCK_0_H1_o(26) <= \SHA256_BLOCK_0_H1_o[26]\;
    SHA256_BLOCK_0_H1_o(25) <= \SHA256_BLOCK_0_H1_o[25]\;
    SHA256_BLOCK_0_H1_o(24) <= \SHA256_BLOCK_0_H1_o[24]\;
    SHA256_BLOCK_0_H1_o(23) <= \SHA256_BLOCK_0_H1_o[23]\;
    SHA256_BLOCK_0_H1_o(22) <= \SHA256_BLOCK_0_H1_o[22]\;
    SHA256_BLOCK_0_H1_o(21) <= \SHA256_BLOCK_0_H1_o[21]\;
    SHA256_BLOCK_0_H1_o(20) <= \SHA256_BLOCK_0_H1_o[20]\;
    SHA256_BLOCK_0_H1_o(19) <= \SHA256_BLOCK_0_H1_o[19]\;
    SHA256_BLOCK_0_H1_o(18) <= \SHA256_BLOCK_0_H1_o[18]\;
    SHA256_BLOCK_0_H1_o(17) <= \SHA256_BLOCK_0_H1_o[17]\;
    SHA256_BLOCK_0_H1_o(16) <= \SHA256_BLOCK_0_H1_o[16]\;
    SHA256_BLOCK_0_H1_o(15) <= \SHA256_BLOCK_0_H1_o[15]\;
    SHA256_BLOCK_0_H1_o(14) <= \SHA256_BLOCK_0_H1_o[14]\;
    SHA256_BLOCK_0_H1_o(13) <= \SHA256_BLOCK_0_H1_o[13]\;
    SHA256_BLOCK_0_H1_o(12) <= \SHA256_BLOCK_0_H1_o[12]\;
    SHA256_BLOCK_0_H1_o(11) <= \SHA256_BLOCK_0_H1_o[11]\;
    SHA256_BLOCK_0_H1_o(10) <= \SHA256_BLOCK_0_H1_o[10]\;
    SHA256_BLOCK_0_H1_o(9) <= \SHA256_BLOCK_0_H1_o[9]\;
    SHA256_BLOCK_0_H1_o(8) <= \SHA256_BLOCK_0_H1_o[8]\;
    SHA256_BLOCK_0_H1_o(7) <= \SHA256_BLOCK_0_H1_o[7]\;
    SHA256_BLOCK_0_H1_o(6) <= \SHA256_BLOCK_0_H1_o[6]\;
    SHA256_BLOCK_0_H1_o(5) <= \SHA256_BLOCK_0_H1_o[5]\;
    SHA256_BLOCK_0_H1_o(4) <= \SHA256_BLOCK_0_H1_o[4]\;
    SHA256_BLOCK_0_H1_o(3) <= \SHA256_BLOCK_0_H1_o[3]\;
    SHA256_BLOCK_0_H1_o(2) <= \SHA256_BLOCK_0_H1_o[2]\;
    SHA256_BLOCK_0_H1_o(1) <= \SHA256_BLOCK_0_H1_o[1]\;
    SHA256_BLOCK_0_H1_o(0) <= \SHA256_BLOCK_0_H1_o[0]\;
    N1_data(31) <= \N1_data[31]\;
    N1_data(30) <= \N1_data[30]\;
    N1_data(29) <= \N1_data[29]\;
    N1_data(28) <= \N1_data[28]\;
    N1_data(27) <= \N1_data[27]\;
    N1_data(26) <= \N1_data[26]\;
    N1_data(25) <= \N1_data[25]\;
    N1_data(24) <= \N1_data[24]\;
    N1_data(23) <= \N1_data[23]\;
    N1_data(22) <= \N1_data[22]\;
    N1_data(21) <= \N1_data[21]\;
    N1_data(20) <= \N1_data[20]\;
    N1_data(19) <= \N1_data[19]\;
    N1_data(18) <= \N1_data[18]\;
    N1_data(17) <= \N1_data[17]\;
    N1_data(16) <= \N1_data[16]\;
    N1_data(15) <= \N1_data[15]\;
    N1_data(14) <= \N1_data[14]\;
    N1_data(13) <= \N1_data[13]\;
    N1_data(12) <= \N1_data[12]\;
    N1_data(11) <= \N1_data[11]\;
    N1_data(10) <= \N1_data[10]\;
    N1_data(9) <= \N1_data[9]\;
    N1_data(8) <= \N1_data[8]\;
    N1_data(7) <= \N1_data[7]\;
    N1_data(6) <= \N1_data[6]\;
    N1_data(5) <= \N1_data[5]\;
    N1_data(4) <= \N1_data[4]\;
    N1_data(3) <= \N1_data[3]\;
    N1_data(2) <= \N1_data[2]\;
    N1_data(1) <= \N1_data[1]\;
    SHA256_BLOCK_0_H2_o(31) <= \SHA256_BLOCK_0_H2_o[31]\;
    SHA256_BLOCK_0_H2_o(30) <= \SHA256_BLOCK_0_H2_o[30]\;
    SHA256_BLOCK_0_H2_o(29) <= \SHA256_BLOCK_0_H2_o[29]\;
    SHA256_BLOCK_0_H2_o(28) <= \SHA256_BLOCK_0_H2_o[28]\;
    SHA256_BLOCK_0_H2_o(27) <= \SHA256_BLOCK_0_H2_o[27]\;
    SHA256_BLOCK_0_H2_o(26) <= \SHA256_BLOCK_0_H2_o[26]\;
    SHA256_BLOCK_0_H2_o(25) <= \SHA256_BLOCK_0_H2_o[25]\;
    SHA256_BLOCK_0_H2_o(24) <= \SHA256_BLOCK_0_H2_o[24]\;
    SHA256_BLOCK_0_H2_o(23) <= \SHA256_BLOCK_0_H2_o[23]\;
    SHA256_BLOCK_0_H2_o(22) <= \SHA256_BLOCK_0_H2_o[22]\;
    SHA256_BLOCK_0_H2_o(21) <= \SHA256_BLOCK_0_H2_o[21]\;
    SHA256_BLOCK_0_H2_o(20) <= \SHA256_BLOCK_0_H2_o[20]\;
    SHA256_BLOCK_0_H2_o(19) <= \SHA256_BLOCK_0_H2_o[19]\;
    SHA256_BLOCK_0_H2_o(18) <= \SHA256_BLOCK_0_H2_o[18]\;
    SHA256_BLOCK_0_H2_o(17) <= \SHA256_BLOCK_0_H2_o[17]\;
    SHA256_BLOCK_0_H2_o(16) <= \SHA256_BLOCK_0_H2_o[16]\;
    SHA256_BLOCK_0_H2_o(15) <= \SHA256_BLOCK_0_H2_o[15]\;
    SHA256_BLOCK_0_H2_o(14) <= \SHA256_BLOCK_0_H2_o[14]\;
    SHA256_BLOCK_0_H2_o(13) <= \SHA256_BLOCK_0_H2_o[13]\;
    SHA256_BLOCK_0_H2_o(12) <= \SHA256_BLOCK_0_H2_o[12]\;
    SHA256_BLOCK_0_H2_o(11) <= \SHA256_BLOCK_0_H2_o[11]\;
    SHA256_BLOCK_0_H2_o(10) <= \SHA256_BLOCK_0_H2_o[10]\;
    SHA256_BLOCK_0_H2_o(9) <= \SHA256_BLOCK_0_H2_o[9]\;
    SHA256_BLOCK_0_H2_o(8) <= \SHA256_BLOCK_0_H2_o[8]\;
    SHA256_BLOCK_0_H2_o(7) <= \SHA256_BLOCK_0_H2_o[7]\;
    SHA256_BLOCK_0_H2_o(6) <= \SHA256_BLOCK_0_H2_o[6]\;
    SHA256_BLOCK_0_H2_o(5) <= \SHA256_BLOCK_0_H2_o[5]\;
    SHA256_BLOCK_0_H2_o(4) <= \SHA256_BLOCK_0_H2_o[4]\;
    SHA256_BLOCK_0_H2_o(3) <= \SHA256_BLOCK_0_H2_o[3]\;
    SHA256_BLOCK_0_H2_o(2) <= \SHA256_BLOCK_0_H2_o[2]\;
    SHA256_BLOCK_0_H2_o(1) <= \SHA256_BLOCK_0_H2_o[1]\;
    SHA256_BLOCK_0_H2_o(0) <= \SHA256_BLOCK_0_H2_o[0]\;
    N2_data(31) <= \N2_data[31]\;
    N2_data(30) <= \N2_data[30]\;
    N2_data(29) <= \N2_data[29]\;
    N2_data(28) <= \N2_data[28]\;
    N2_data(27) <= \N2_data[27]\;
    N2_data(26) <= \N2_data[26]\;
    N2_data(25) <= \N2_data[25]\;
    N2_data(24) <= \N2_data[24]\;
    N2_data(23) <= \N2_data[23]\;
    N2_data(22) <= \N2_data[22]\;
    N2_data(21) <= \N2_data[21]\;
    N2_data(20) <= \N2_data[20]\;
    N2_data(19) <= \N2_data[19]\;
    N2_data(18) <= \N2_data[18]\;
    N2_data(17) <= \N2_data[17]\;
    N2_data(16) <= \N2_data[16]\;
    N2_data(15) <= \N2_data[15]\;
    N2_data(14) <= \N2_data[14]\;
    N2_data(13) <= \N2_data[13]\;
    N2_data(12) <= \N2_data[12]\;
    N2_data(11) <= \N2_data[11]\;
    N2_data(10) <= \N2_data[10]\;
    N2_data(9) <= \N2_data[9]\;
    N2_data(8) <= \N2_data[8]\;
    N2_data(7) <= \N2_data[7]\;
    N2_data(6) <= \N2_data[6]\;
    N2_data(5) <= \N2_data[5]\;
    N2_data(4) <= \N2_data[4]\;
    N2_data(3) <= \N2_data[3]\;
    N2_data(2) <= \N2_data[2]\;
    N2_data(1) <= \N2_data[1]\;
    SHA256_BLOCK_0_H3_o(31) <= \SHA256_BLOCK_0_H3_o[31]\;
    SHA256_BLOCK_0_H3_o(30) <= \SHA256_BLOCK_0_H3_o[30]\;
    SHA256_BLOCK_0_H3_o(29) <= \SHA256_BLOCK_0_H3_o[29]\;
    SHA256_BLOCK_0_H3_o(28) <= \SHA256_BLOCK_0_H3_o[28]\;
    SHA256_BLOCK_0_H3_o(27) <= \SHA256_BLOCK_0_H3_o[27]\;
    SHA256_BLOCK_0_H3_o(26) <= \SHA256_BLOCK_0_H3_o[26]\;
    SHA256_BLOCK_0_H3_o(25) <= \SHA256_BLOCK_0_H3_o[25]\;
    SHA256_BLOCK_0_H3_o(24) <= \SHA256_BLOCK_0_H3_o[24]\;
    SHA256_BLOCK_0_H3_o(23) <= \SHA256_BLOCK_0_H3_o[23]\;
    SHA256_BLOCK_0_H3_o(22) <= \SHA256_BLOCK_0_H3_o[22]\;
    SHA256_BLOCK_0_H3_o(21) <= \SHA256_BLOCK_0_H3_o[21]\;
    SHA256_BLOCK_0_H3_o(20) <= \SHA256_BLOCK_0_H3_o[20]\;
    SHA256_BLOCK_0_H3_o(19) <= \SHA256_BLOCK_0_H3_o[19]\;
    SHA256_BLOCK_0_H3_o(18) <= \SHA256_BLOCK_0_H3_o[18]\;
    SHA256_BLOCK_0_H3_o(17) <= \SHA256_BLOCK_0_H3_o[17]\;
    SHA256_BLOCK_0_H3_o(16) <= \SHA256_BLOCK_0_H3_o[16]\;
    SHA256_BLOCK_0_H3_o(15) <= \SHA256_BLOCK_0_H3_o[15]\;
    SHA256_BLOCK_0_H3_o(14) <= \SHA256_BLOCK_0_H3_o[14]\;
    SHA256_BLOCK_0_H3_o(13) <= \SHA256_BLOCK_0_H3_o[13]\;
    SHA256_BLOCK_0_H3_o(12) <= \SHA256_BLOCK_0_H3_o[12]\;
    SHA256_BLOCK_0_H3_o(11) <= \SHA256_BLOCK_0_H3_o[11]\;
    SHA256_BLOCK_0_H3_o(10) <= \SHA256_BLOCK_0_H3_o[10]\;
    SHA256_BLOCK_0_H3_o(9) <= \SHA256_BLOCK_0_H3_o[9]\;
    SHA256_BLOCK_0_H3_o(8) <= \SHA256_BLOCK_0_H3_o[8]\;
    SHA256_BLOCK_0_H3_o(7) <= \SHA256_BLOCK_0_H3_o[7]\;
    SHA256_BLOCK_0_H3_o(6) <= \SHA256_BLOCK_0_H3_o[6]\;
    SHA256_BLOCK_0_H3_o(5) <= \SHA256_BLOCK_0_H3_o[5]\;
    SHA256_BLOCK_0_H3_o(4) <= \SHA256_BLOCK_0_H3_o[4]\;
    SHA256_BLOCK_0_H3_o(3) <= \SHA256_BLOCK_0_H3_o[3]\;
    SHA256_BLOCK_0_H3_o(2) <= \SHA256_BLOCK_0_H3_o[2]\;
    SHA256_BLOCK_0_H3_o(1) <= \SHA256_BLOCK_0_H3_o[1]\;
    SHA256_BLOCK_0_H3_o(0) <= \SHA256_BLOCK_0_H3_o[0]\;
    N3_data(31) <= \N3_data[31]\;
    N3_data(30) <= \N3_data[30]\;
    N3_data(29) <= \N3_data[29]\;
    N3_data(28) <= \N3_data[28]\;
    N3_data(27) <= \N3_data[27]\;
    N3_data(26) <= \N3_data[26]\;
    N3_data(25) <= \N3_data[25]\;
    N3_data(24) <= \N3_data[24]\;
    N3_data(23) <= \N3_data[23]\;
    N3_data(22) <= \N3_data[22]\;
    N3_data(21) <= \N3_data[21]\;
    N3_data(20) <= \N3_data[20]\;
    N3_data(19) <= \N3_data[19]\;
    N3_data(18) <= \N3_data[18]\;
    N3_data(17) <= \N3_data[17]\;
    N3_data(16) <= \N3_data[16]\;
    N3_data(15) <= \N3_data[15]\;
    N3_data(14) <= \N3_data[14]\;
    N3_data(13) <= \N3_data[13]\;
    N3_data(12) <= \N3_data[12]\;
    N3_data(11) <= \N3_data[11]\;
    N3_data(10) <= \N3_data[10]\;
    N3_data(9) <= \N3_data[9]\;
    N3_data(8) <= \N3_data[8]\;
    N3_data(7) <= \N3_data[7]\;
    N3_data(6) <= \N3_data[6]\;
    N3_data(5) <= \N3_data[5]\;
    N3_data(4) <= \N3_data[4]\;
    N3_data(3) <= \N3_data[3]\;
    N3_data(2) <= \N3_data[2]\;
    N3_data(1) <= \N3_data[1]\;
    SHA256_BLOCK_0_H4_o(31) <= \SHA256_BLOCK_0_H4_o[31]\;
    SHA256_BLOCK_0_H4_o(30) <= \SHA256_BLOCK_0_H4_o[30]\;
    SHA256_BLOCK_0_H4_o(29) <= \SHA256_BLOCK_0_H4_o[29]\;
    SHA256_BLOCK_0_H4_o(28) <= \SHA256_BLOCK_0_H4_o[28]\;
    SHA256_BLOCK_0_H4_o(27) <= \SHA256_BLOCK_0_H4_o[27]\;
    SHA256_BLOCK_0_H4_o(26) <= \SHA256_BLOCK_0_H4_o[26]\;
    SHA256_BLOCK_0_H4_o(25) <= \SHA256_BLOCK_0_H4_o[25]\;
    SHA256_BLOCK_0_H4_o(24) <= \SHA256_BLOCK_0_H4_o[24]\;
    SHA256_BLOCK_0_H4_o(23) <= \SHA256_BLOCK_0_H4_o[23]\;
    SHA256_BLOCK_0_H4_o(22) <= \SHA256_BLOCK_0_H4_o[22]\;
    SHA256_BLOCK_0_H4_o(21) <= \SHA256_BLOCK_0_H4_o[21]\;
    SHA256_BLOCK_0_H4_o(20) <= \SHA256_BLOCK_0_H4_o[20]\;
    SHA256_BLOCK_0_H4_o(19) <= \SHA256_BLOCK_0_H4_o[19]\;
    SHA256_BLOCK_0_H4_o(18) <= \SHA256_BLOCK_0_H4_o[18]\;
    SHA256_BLOCK_0_H4_o(17) <= \SHA256_BLOCK_0_H4_o[17]\;
    SHA256_BLOCK_0_H4_o(16) <= \SHA256_BLOCK_0_H4_o[16]\;
    SHA256_BLOCK_0_H4_o(15) <= \SHA256_BLOCK_0_H4_o[15]\;
    SHA256_BLOCK_0_H4_o(14) <= \SHA256_BLOCK_0_H4_o[14]\;
    SHA256_BLOCK_0_H4_o(13) <= \SHA256_BLOCK_0_H4_o[13]\;
    SHA256_BLOCK_0_H4_o(12) <= \SHA256_BLOCK_0_H4_o[12]\;
    SHA256_BLOCK_0_H4_o(11) <= \SHA256_BLOCK_0_H4_o[11]\;
    SHA256_BLOCK_0_H4_o(10) <= \SHA256_BLOCK_0_H4_o[10]\;
    SHA256_BLOCK_0_H4_o(9) <= \SHA256_BLOCK_0_H4_o[9]\;
    SHA256_BLOCK_0_H4_o(8) <= \SHA256_BLOCK_0_H4_o[8]\;
    SHA256_BLOCK_0_H4_o(7) <= \SHA256_BLOCK_0_H4_o[7]\;
    SHA256_BLOCK_0_H4_o(6) <= \SHA256_BLOCK_0_H4_o[6]\;
    SHA256_BLOCK_0_H4_o(5) <= \SHA256_BLOCK_0_H4_o[5]\;
    SHA256_BLOCK_0_H4_o(4) <= \SHA256_BLOCK_0_H4_o[4]\;
    SHA256_BLOCK_0_H4_o(3) <= \SHA256_BLOCK_0_H4_o[3]\;
    SHA256_BLOCK_0_H4_o(2) <= \SHA256_BLOCK_0_H4_o[2]\;
    SHA256_BLOCK_0_H4_o(1) <= \SHA256_BLOCK_0_H4_o[1]\;
    SHA256_BLOCK_0_H4_o(0) <= \SHA256_BLOCK_0_H4_o[0]\;
    N4_data(31) <= \N4_data[31]\;
    N4_data(30) <= \N4_data[30]\;
    N4_data(29) <= \N4_data[29]\;
    N4_data(28) <= \N4_data[28]\;
    N4_data(27) <= \N4_data[27]\;
    N4_data(26) <= \N4_data[26]\;
    N4_data(25) <= \N4_data[25]\;
    N4_data(24) <= \N4_data[24]\;
    N4_data(23) <= \N4_data[23]\;
    N4_data(22) <= \N4_data[22]\;
    N4_data(21) <= \N4_data[21]\;
    N4_data(20) <= \N4_data[20]\;
    N4_data(19) <= \N4_data[19]\;
    N4_data(18) <= \N4_data[18]\;
    N4_data(17) <= \N4_data[17]\;
    N4_data(16) <= \N4_data[16]\;
    N4_data(15) <= \N4_data[15]\;
    N4_data(14) <= \N4_data[14]\;
    N4_data(13) <= \N4_data[13]\;
    N4_data(12) <= \N4_data[12]\;
    N4_data(11) <= \N4_data[11]\;
    N4_data(10) <= \N4_data[10]\;
    N4_data(9) <= \N4_data[9]\;
    N4_data(8) <= \N4_data[8]\;
    N4_data(7) <= \N4_data[7]\;
    N4_data(6) <= \N4_data[6]\;
    N4_data(5) <= \N4_data[5]\;
    N4_data(4) <= \N4_data[4]\;
    N4_data(3) <= \N4_data[3]\;
    N4_data(2) <= \N4_data[2]\;
    N4_data(1) <= \N4_data[1]\;
    N5_data(31) <= \N5_data[31]\;
    N5_data(30) <= \N5_data[30]\;
    N5_data(29) <= \N5_data[29]\;
    N5_data(28) <= \N5_data[28]\;
    N5_data(27) <= \N5_data[27]\;
    N5_data(26) <= \N5_data[26]\;
    N5_data(25) <= \N5_data[25]\;
    N5_data(24) <= \N5_data[24]\;
    N5_data(23) <= \N5_data[23]\;
    N5_data(22) <= \N5_data[22]\;
    N5_data(21) <= \N5_data[21]\;
    N5_data(20) <= \N5_data[20]\;
    N5_data(19) <= \N5_data[19]\;
    N5_data(18) <= \N5_data[18]\;
    N5_data(17) <= \N5_data[17]\;
    N5_data(16) <= \N5_data[16]\;
    N5_data(15) <= \N5_data[15]\;
    N5_data(14) <= \N5_data[14]\;
    N5_data(13) <= \N5_data[13]\;
    N5_data(12) <= \N5_data[12]\;
    N5_data(11) <= \N5_data[11]\;
    N5_data(10) <= \N5_data[10]\;
    N5_data(9) <= \N5_data[9]\;
    N5_data(8) <= \N5_data[8]\;
    N5_data(7) <= \N5_data[7]\;
    N5_data(6) <= \N5_data[6]\;
    N5_data(5) <= \N5_data[5]\;
    N5_data(4) <= \N5_data[4]\;
    N5_data(3) <= \N5_data[3]\;
    N5_data(2) <= \N5_data[2]\;
    N5_data(1) <= \N5_data[1]\;
    SHA256_BLOCK_0_H5_o(31) <= \SHA256_BLOCK_0_H5_o[31]\;
    SHA256_BLOCK_0_H5_o(30) <= \SHA256_BLOCK_0_H5_o[30]\;
    SHA256_BLOCK_0_H5_o(29) <= \SHA256_BLOCK_0_H5_o[29]\;
    SHA256_BLOCK_0_H5_o(28) <= \SHA256_BLOCK_0_H5_o[28]\;
    SHA256_BLOCK_0_H5_o(27) <= \SHA256_BLOCK_0_H5_o[27]\;
    SHA256_BLOCK_0_H5_o(26) <= \SHA256_BLOCK_0_H5_o[26]\;
    SHA256_BLOCK_0_H5_o(25) <= \SHA256_BLOCK_0_H5_o[25]\;
    SHA256_BLOCK_0_H5_o(24) <= \SHA256_BLOCK_0_H5_o[24]\;
    SHA256_BLOCK_0_H5_o(23) <= \SHA256_BLOCK_0_H5_o[23]\;
    SHA256_BLOCK_0_H5_o(22) <= \SHA256_BLOCK_0_H5_o[22]\;
    SHA256_BLOCK_0_H5_o(21) <= \SHA256_BLOCK_0_H5_o[21]\;
    SHA256_BLOCK_0_H5_o(20) <= \SHA256_BLOCK_0_H5_o[20]\;
    SHA256_BLOCK_0_H5_o(19) <= \SHA256_BLOCK_0_H5_o[19]\;
    SHA256_BLOCK_0_H5_o(18) <= \SHA256_BLOCK_0_H5_o[18]\;
    SHA256_BLOCK_0_H5_o(17) <= \SHA256_BLOCK_0_H5_o[17]\;
    SHA256_BLOCK_0_H5_o(16) <= \SHA256_BLOCK_0_H5_o[16]\;
    SHA256_BLOCK_0_H5_o(15) <= \SHA256_BLOCK_0_H5_o[15]\;
    SHA256_BLOCK_0_H5_o(14) <= \SHA256_BLOCK_0_H5_o[14]\;
    SHA256_BLOCK_0_H5_o(13) <= \SHA256_BLOCK_0_H5_o[13]\;
    SHA256_BLOCK_0_H5_o(12) <= \SHA256_BLOCK_0_H5_o[12]\;
    SHA256_BLOCK_0_H5_o(11) <= \SHA256_BLOCK_0_H5_o[11]\;
    SHA256_BLOCK_0_H5_o(10) <= \SHA256_BLOCK_0_H5_o[10]\;
    SHA256_BLOCK_0_H5_o(9) <= \SHA256_BLOCK_0_H5_o[9]\;
    SHA256_BLOCK_0_H5_o(8) <= \SHA256_BLOCK_0_H5_o[8]\;
    SHA256_BLOCK_0_H5_o(7) <= \SHA256_BLOCK_0_H5_o[7]\;
    SHA256_BLOCK_0_H5_o(6) <= \SHA256_BLOCK_0_H5_o[6]\;
    SHA256_BLOCK_0_H5_o(5) <= \SHA256_BLOCK_0_H5_o[5]\;
    SHA256_BLOCK_0_H5_o(4) <= \SHA256_BLOCK_0_H5_o[4]\;
    SHA256_BLOCK_0_H5_o(3) <= \SHA256_BLOCK_0_H5_o[3]\;
    SHA256_BLOCK_0_H5_o(2) <= \SHA256_BLOCK_0_H5_o[2]\;
    SHA256_BLOCK_0_H5_o(1) <= \SHA256_BLOCK_0_H5_o[1]\;
    SHA256_BLOCK_0_H5_o(0) <= \SHA256_BLOCK_0_H5_o[0]\;
    SHA256_BLOCK_0_H6_o(31) <= \SHA256_BLOCK_0_H6_o[31]\;
    SHA256_BLOCK_0_H6_o(30) <= \SHA256_BLOCK_0_H6_o[30]\;
    SHA256_BLOCK_0_H6_o(29) <= \SHA256_BLOCK_0_H6_o[29]\;
    SHA256_BLOCK_0_H6_o(28) <= \SHA256_BLOCK_0_H6_o[28]\;
    SHA256_BLOCK_0_H6_o(27) <= \SHA256_BLOCK_0_H6_o[27]\;
    SHA256_BLOCK_0_H6_o(26) <= \SHA256_BLOCK_0_H6_o[26]\;
    SHA256_BLOCK_0_H6_o(25) <= \SHA256_BLOCK_0_H6_o[25]\;
    SHA256_BLOCK_0_H6_o(24) <= \SHA256_BLOCK_0_H6_o[24]\;
    SHA256_BLOCK_0_H6_o(23) <= \SHA256_BLOCK_0_H6_o[23]\;
    SHA256_BLOCK_0_H6_o(22) <= \SHA256_BLOCK_0_H6_o[22]\;
    SHA256_BLOCK_0_H6_o(21) <= \SHA256_BLOCK_0_H6_o[21]\;
    SHA256_BLOCK_0_H6_o(20) <= \SHA256_BLOCK_0_H6_o[20]\;
    SHA256_BLOCK_0_H6_o(19) <= \SHA256_BLOCK_0_H6_o[19]\;
    SHA256_BLOCK_0_H6_o(18) <= \SHA256_BLOCK_0_H6_o[18]\;
    SHA256_BLOCK_0_H6_o(17) <= \SHA256_BLOCK_0_H6_o[17]\;
    SHA256_BLOCK_0_H6_o(16) <= \SHA256_BLOCK_0_H6_o[16]\;
    SHA256_BLOCK_0_H6_o(15) <= \SHA256_BLOCK_0_H6_o[15]\;
    SHA256_BLOCK_0_H6_o(14) <= \SHA256_BLOCK_0_H6_o[14]\;
    SHA256_BLOCK_0_H6_o(13) <= \SHA256_BLOCK_0_H6_o[13]\;
    SHA256_BLOCK_0_H6_o(12) <= \SHA256_BLOCK_0_H6_o[12]\;
    SHA256_BLOCK_0_H6_o(11) <= \SHA256_BLOCK_0_H6_o[11]\;
    SHA256_BLOCK_0_H6_o(10) <= \SHA256_BLOCK_0_H6_o[10]\;
    SHA256_BLOCK_0_H6_o(9) <= \SHA256_BLOCK_0_H6_o[9]\;
    SHA256_BLOCK_0_H6_o(8) <= \SHA256_BLOCK_0_H6_o[8]\;
    SHA256_BLOCK_0_H6_o(7) <= \SHA256_BLOCK_0_H6_o[7]\;
    SHA256_BLOCK_0_H6_o(6) <= \SHA256_BLOCK_0_H6_o[6]\;
    SHA256_BLOCK_0_H6_o(5) <= \SHA256_BLOCK_0_H6_o[5]\;
    SHA256_BLOCK_0_H6_o(4) <= \SHA256_BLOCK_0_H6_o[4]\;
    SHA256_BLOCK_0_H6_o(3) <= \SHA256_BLOCK_0_H6_o[3]\;
    SHA256_BLOCK_0_H6_o(2) <= \SHA256_BLOCK_0_H6_o[2]\;
    SHA256_BLOCK_0_H6_o(1) <= \SHA256_BLOCK_0_H6_o[1]\;
    SHA256_BLOCK_0_H6_o(0) <= \SHA256_BLOCK_0_H6_o[0]\;
    N6_data(31) <= \N6_data[31]\;
    N6_data(30) <= \N6_data[30]\;
    N6_data(29) <= \N6_data[29]\;
    N6_data(28) <= \N6_data[28]\;
    N6_data(27) <= \N6_data[27]\;
    N6_data(26) <= \N6_data[26]\;
    N6_data(25) <= \N6_data[25]\;
    N6_data(24) <= \N6_data[24]\;
    N6_data(23) <= \N6_data[23]\;
    N6_data(22) <= \N6_data[22]\;
    N6_data(21) <= \N6_data[21]\;
    N6_data(20) <= \N6_data[20]\;
    N6_data(19) <= \N6_data[19]\;
    N6_data(18) <= \N6_data[18]\;
    N6_data(17) <= \N6_data[17]\;
    N6_data(16) <= \N6_data[16]\;
    N6_data(15) <= \N6_data[15]\;
    N6_data(14) <= \N6_data[14]\;
    N6_data(13) <= \N6_data[13]\;
    N6_data(12) <= \N6_data[12]\;
    N6_data(11) <= \N6_data[11]\;
    N6_data(10) <= \N6_data[10]\;
    N6_data(9) <= \N6_data[9]\;
    N6_data(8) <= \N6_data[8]\;
    N6_data(7) <= \N6_data[7]\;
    N6_data(6) <= \N6_data[6]\;
    N6_data(5) <= \N6_data[5]\;
    N6_data(4) <= \N6_data[4]\;
    N6_data(3) <= \N6_data[3]\;
    N6_data(2) <= \N6_data[2]\;
    N6_data(1) <= \N6_data[1]\;
    SHA256_BLOCK_0_H7_o(31) <= \SHA256_BLOCK_0_H7_o[31]\;
    SHA256_BLOCK_0_H7_o(30) <= \SHA256_BLOCK_0_H7_o[30]\;
    SHA256_BLOCK_0_H7_o(29) <= \SHA256_BLOCK_0_H7_o[29]\;
    SHA256_BLOCK_0_H7_o(28) <= \SHA256_BLOCK_0_H7_o[28]\;
    SHA256_BLOCK_0_H7_o(27) <= \SHA256_BLOCK_0_H7_o[27]\;
    SHA256_BLOCK_0_H7_o(26) <= \SHA256_BLOCK_0_H7_o[26]\;
    SHA256_BLOCK_0_H7_o(25) <= \SHA256_BLOCK_0_H7_o[25]\;
    SHA256_BLOCK_0_H7_o(24) <= \SHA256_BLOCK_0_H7_o[24]\;
    SHA256_BLOCK_0_H7_o(23) <= \SHA256_BLOCK_0_H7_o[23]\;
    SHA256_BLOCK_0_H7_o(22) <= \SHA256_BLOCK_0_H7_o[22]\;
    SHA256_BLOCK_0_H7_o(21) <= \SHA256_BLOCK_0_H7_o[21]\;
    SHA256_BLOCK_0_H7_o(20) <= \SHA256_BLOCK_0_H7_o[20]\;
    SHA256_BLOCK_0_H7_o(19) <= \SHA256_BLOCK_0_H7_o[19]\;
    SHA256_BLOCK_0_H7_o(18) <= \SHA256_BLOCK_0_H7_o[18]\;
    SHA256_BLOCK_0_H7_o(17) <= \SHA256_BLOCK_0_H7_o[17]\;
    SHA256_BLOCK_0_H7_o(16) <= \SHA256_BLOCK_0_H7_o[16]\;
    SHA256_BLOCK_0_H7_o(15) <= \SHA256_BLOCK_0_H7_o[15]\;
    SHA256_BLOCK_0_H7_o(14) <= \SHA256_BLOCK_0_H7_o[14]\;
    SHA256_BLOCK_0_H7_o(13) <= \SHA256_BLOCK_0_H7_o[13]\;
    SHA256_BLOCK_0_H7_o(12) <= \SHA256_BLOCK_0_H7_o[12]\;
    SHA256_BLOCK_0_H7_o(11) <= \SHA256_BLOCK_0_H7_o[11]\;
    SHA256_BLOCK_0_H7_o(10) <= \SHA256_BLOCK_0_H7_o[10]\;
    SHA256_BLOCK_0_H7_o(9) <= \SHA256_BLOCK_0_H7_o[9]\;
    SHA256_BLOCK_0_H7_o(8) <= \SHA256_BLOCK_0_H7_o[8]\;
    SHA256_BLOCK_0_H7_o(7) <= \SHA256_BLOCK_0_H7_o[7]\;
    SHA256_BLOCK_0_H7_o(6) <= \SHA256_BLOCK_0_H7_o[6]\;
    SHA256_BLOCK_0_H7_o(5) <= \SHA256_BLOCK_0_H7_o[5]\;
    SHA256_BLOCK_0_H7_o(4) <= \SHA256_BLOCK_0_H7_o[4]\;
    SHA256_BLOCK_0_H7_o(3) <= \SHA256_BLOCK_0_H7_o[3]\;
    SHA256_BLOCK_0_H7_o(2) <= \SHA256_BLOCK_0_H7_o[2]\;
    SHA256_BLOCK_0_H7_o(1) <= \SHA256_BLOCK_0_H7_o[1]\;
    SHA256_BLOCK_0_H7_o(0) <= \SHA256_BLOCK_0_H7_o[0]\;
    N7_data(31) <= \N7_data[31]\;
    N7_data(30) <= \N7_data[30]\;
    N7_data(29) <= \N7_data[29]\;
    N7_data(28) <= \N7_data[28]\;
    N7_data(27) <= \N7_data[27]\;
    N7_data(26) <= \N7_data[26]\;
    N7_data(25) <= \N7_data[25]\;
    N7_data(24) <= \N7_data[24]\;
    N7_data(23) <= \N7_data[23]\;
    N7_data(22) <= \N7_data[22]\;
    N7_data(21) <= \N7_data[21]\;
    N7_data(20) <= \N7_data[20]\;
    N7_data(19) <= \N7_data[19]\;
    N7_data(18) <= \N7_data[18]\;
    N7_data(17) <= \N7_data[17]\;
    N7_data(16) <= \N7_data[16]\;
    N7_data(15) <= \N7_data[15]\;
    N7_data(14) <= \N7_data[14]\;
    N7_data(13) <= \N7_data[13]\;
    N7_data(12) <= \N7_data[12]\;
    N7_data(11) <= \N7_data[11]\;
    N7_data(10) <= \N7_data[10]\;
    N7_data(9) <= \N7_data[9]\;
    N7_data(8) <= \N7_data[8]\;
    N7_data(7) <= \N7_data[7]\;
    N7_data(6) <= \N7_data[6]\;
    N7_data(5) <= \N7_data[5]\;
    N7_data(4) <= \N7_data[4]\;
    N7_data(3) <= \N7_data[3]\;
    N7_data(2) <= \N7_data[2]\;
    N7_data(1) <= \N7_data[1]\;
    next_reg_H0_cry_0_0_Y <= \next_reg_H0_cry_0_0_Y\;
    next_reg_H1_cry_0_0_Y <= \next_reg_H1_cry_0_0_Y\;
    next_reg_H2_cry_0_0_Y <= \next_reg_H2_cry_0_0_Y\;
    next_reg_H3_cry_0_0_Y <= \next_reg_H3_cry_0_0_Y\;
    next_reg_H4_cry_0_0_Y <= \next_reg_H4_cry_0_0_Y\;
    next_reg_H5_cry_0_0_Y <= \next_reg_H5_cry_0_0_Y\;
    next_reg_H6_cry_0_0_Y <= \next_reg_H6_cry_0_0_Y\;
    next_reg_H7_cry_0_0_Y <= \next_reg_H7_cry_0_0_Y\;

    \reg_H7[31]\ : SLE
      port map(D => \N7_data[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[31]\);
    
    next_reg_H2_cry_21_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[21]\, B => 
        hash_control_st_reg_i(6), C => R2_data(21), D => 
        GND_net_1, FCI => next_reg_H2_cry_20, S => \N2_data[21]\, 
        Y => OPEN, FCO => next_reg_H2_cry_21);
    
    \reg_H4[12]\ : SLE
      port map(D => \N4_data[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[12]\);
    
    next_reg_H1_cry_8_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[8]\, B => 
        hash_control_st_reg_i(6), C => R1_data(8), D => GND_net_1, 
        FCI => next_reg_H1_cry_7, S => \N1_data[8]\, Y => OPEN, 
        FCO => next_reg_H1_cry_8);
    
    \reg_H3[4]\ : SLE
      port map(D => \N3_data[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[4]\);
    
    next_reg_H7_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[14]\, B => 
        hash_control_st_reg_i(6), C => R7_data(14), D => 
        GND_net_1, FCI => next_reg_H7_cry_13, S => \N7_data[14]\, 
        Y => OPEN, FCO => next_reg_H7_cry_14);
    
    \reg_H4[17]\ : SLE
      port map(D => \N4_data[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[17]\);
    
    next_reg_H4_cry_22_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[22]\, B => 
        hash_control_st_reg_i(6), C => R4_data(22), D => 
        GND_net_1, FCI => next_reg_H4_cry_21, S => \N4_data[22]\, 
        Y => OPEN, FCO => next_reg_H4_cry_22);
    
    \reg_H1[2]\ : SLE
      port map(D => \N1_data[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[2]\);
    
    next_reg_H7_cry_25_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[25]\, B => 
        hash_control_st_reg_i(6), C => R7_data(25), D => 
        GND_net_1, FCI => next_reg_H7_cry_24, S => \N7_data[25]\, 
        Y => OPEN, FCO => next_reg_H7_cry_25);
    
    next_reg_H4_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[20]\, B => 
        hash_control_st_reg_i(6), C => R4_data(20), D => 
        GND_net_1, FCI => next_reg_H4_cry_19, S => \N4_data[20]\, 
        Y => OPEN, FCO => next_reg_H4_cry_20);
    
    \reg_H6[5]\ : SLE
      port map(D => \N6_data[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[5]\);
    
    next_reg_H0_cry_11_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[11]\, B => 
        hash_control_st_reg_i(6), C => R0_data(11), D => 
        GND_net_1, FCI => next_reg_H0_cry_10, S => \N0_data[11]\, 
        Y => OPEN, FCO => next_reg_H0_cry_11);
    
    \reg_H1[5]\ : SLE
      port map(D => \N1_data[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[5]\);
    
    next_reg_H5_cry_25_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[25]\, B => 
        hash_control_st_reg_i(6), C => R5_data(25), D => 
        GND_net_1, FCI => next_reg_H5_cry_24, S => \N5_data[25]\, 
        Y => OPEN, FCO => next_reg_H5_cry_25);
    
    \reg_H5[12]\ : SLE
      port map(D => \N5_data[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[12]\);
    
    \reg_H3[20]\ : SLE
      port map(D => \N3_data[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[20]\);
    
    next_reg_H5_s_31 : ARI1
      generic map(INIT => x"47D00")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R5_data(31), D => \SHA256_BLOCK_0_H5_o[31]\, FCI => 
        next_reg_H5_cry_30, S => \N5_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    \reg_H0[16]\ : SLE
      port map(D => \N0_data[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[16]\);
    
    next_reg_H3_cry_11_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[11]\, B => 
        hash_control_st_reg_i(6), C => R3_data(11), D => 
        GND_net_1, FCI => next_reg_H3_cry_10, S => \N3_data[11]\, 
        Y => OPEN, FCO => next_reg_H3_cry_11);
    
    \reg_H5[17]\ : SLE
      port map(D => \N5_data[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[17]\);
    
    next_reg_H5_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[14]\, B => 
        hash_control_st_reg_i(6), C => R5_data(14), D => 
        GND_net_1, FCI => next_reg_H5_cry_13, S => \N5_data[14]\, 
        Y => OPEN, FCO => next_reg_H5_cry_14);
    
    next_reg_H1_cry_13_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[13]\, B => 
        hash_control_st_reg_i(6), C => R1_data(13), D => 
        GND_net_1, FCI => next_reg_H1_cry_12, S => \N1_data[13]\, 
        Y => OPEN, FCO => next_reg_H1_cry_13);
    
    \reg_H3[30]\ : SLE
      port map(D => \N3_data[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[30]\);
    
    next_reg_H3_cry_29_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[29]\, B => 
        hash_control_st_reg_i(6), C => R3_data(29), D => 
        GND_net_1, FCI => next_reg_H3_cry_28, S => \N3_data[29]\, 
        Y => OPEN, FCO => next_reg_H3_cry_29);
    
    \reg_H1[8]\ : SLE
      port map(D => \N1_data[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[8]\);
    
    next_reg_H7_cry_4_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[4]\, B => 
        hash_control_st_reg_i(6), C => R7_data(4), D => GND_net_1, 
        FCI => next_reg_H7_cry_3, S => \N7_data[4]\, Y => OPEN, 
        FCO => next_reg_H7_cry_4);
    
    \reg_H5[22]\ : SLE
      port map(D => \N5_data[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[22]\);
    
    next_reg_H6_cry_18_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[18]\, B => 
        hash_control_st_reg_i(6), C => R6_data(18), D => 
        GND_net_1, FCI => next_reg_H6_cry_17, S => \N6_data[18]\, 
        Y => OPEN, FCO => next_reg_H6_cry_18);
    
    \reg_H1[4]\ : SLE
      port map(D => \N1_data[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[4]\);
    
    \reg_H1[21]\ : SLE
      port map(D => \N1_data[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[21]\);
    
    next_reg_H5_cry_9_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[9]\, B => 
        hash_control_st_reg_i(6), C => R5_data(9), D => GND_net_1, 
        FCI => next_reg_H5_cry_8, S => \N5_data[9]\, Y => OPEN, 
        FCO => next_reg_H5_cry_9);
    
    next_reg_H2_cry_0_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[0]\, B => 
        hash_control_st_reg_i(6), C => R2_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H2_cry_0_0_Y\, 
        FCO => next_reg_H2_cry_0);
    
    next_reg_H6_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[24]\, B => 
        hash_control_st_reg_i(6), C => R6_data(24), D => 
        GND_net_1, FCI => next_reg_H6_cry_23, S => \N6_data[24]\, 
        Y => OPEN, FCO => next_reg_H6_cry_24);
    
    \reg_H7[28]\ : SLE
      port map(D => \N7_data[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[28]\);
    
    \reg_H5[31]\ : SLE
      port map(D => \N5_data[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[31]\);
    
    \reg_H5[27]\ : SLE
      port map(D => \N5_data[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[27]\);
    
    next_reg_H7_cry_30_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[30]\, B => 
        hash_control_st_reg_i(6), C => R7_data(30), D => 
        GND_net_1, FCI => next_reg_H7_cry_29, S => \N7_data[30]\, 
        Y => OPEN, FCO => next_reg_H7_cry_30);
    
    \reg_H7[0]\ : SLE
      port map(D => \next_reg_H7_cry_0_0_Y\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[0]\);
    
    \reg_H6[20]\ : SLE
      port map(D => \N6_data[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[20]\);
    
    next_reg_H2_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[15]\, B => 
        hash_control_st_reg_i(6), C => R2_data(15), D => 
        GND_net_1, FCI => next_reg_H2_cry_14, S => \N2_data[15]\, 
        Y => OPEN, FCO => next_reg_H2_cry_15);
    
    \reg_H6[6]\ : SLE
      port map(D => \N6_data[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[6]\);
    
    next_reg_H6_cry_4_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[4]\, B => 
        hash_control_st_reg_i(6), C => R6_data(4), D => GND_net_1, 
        FCI => next_reg_H6_cry_3, S => \N6_data[4]\, Y => OPEN, 
        FCO => next_reg_H6_cry_4);
    
    \reg_H4[7]\ : SLE
      port map(D => \N4_data[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[7]\);
    
    \reg_H4[13]\ : SLE
      port map(D => \N4_data[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[13]\);
    
    next_reg_H4_cry_13_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[13]\, B => 
        hash_control_st_reg_i(6), C => R4_data(13), D => 
        GND_net_1, FCI => next_reg_H4_cry_12, S => \N4_data[13]\, 
        Y => OPEN, FCO => next_reg_H4_cry_13);
    
    next_reg_H0_cry_9_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[9]\, B => 
        hash_control_st_reg_i(6), C => R0_data(9), D => GND_net_1, 
        FCI => next_reg_H0_cry_8, S => \N0_data[9]\, Y => OPEN, 
        FCO => next_reg_H0_cry_9);
    
    \reg_H4[14]\ : SLE
      port map(D => \N4_data[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[14]\);
    
    \reg_H2[9]\ : SLE
      port map(D => \N2_data[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[9]\);
    
    next_reg_H1_cry_25_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[25]\, B => 
        hash_control_st_reg_i(6), C => R1_data(25), D => 
        GND_net_1, FCI => next_reg_H1_cry_24, S => \N1_data[25]\, 
        Y => OPEN, FCO => next_reg_H1_cry_25);
    
    \reg_H2[22]\ : SLE
      port map(D => \N2_data[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[22]\);
    
    \reg_H3[29]\ : SLE
      port map(D => \N3_data[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[29]\);
    
    \reg_H7[25]\ : SLE
      port map(D => \N7_data[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[25]\);
    
    \reg_H0[20]\ : SLE
      port map(D => \N0_data[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[20]\);
    
    \reg_H4[4]\ : SLE
      port map(D => \N4_data[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[4]\);
    
    \reg_H2[27]\ : SLE
      port map(D => \N2_data[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[27]\);
    
    next_reg_H6_cry_30_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[30]\, B => 
        hash_control_st_reg_i(6), C => R6_data(30), D => 
        GND_net_1, FCI => next_reg_H6_cry_29, S => \N6_data[30]\, 
        Y => OPEN, FCO => next_reg_H6_cry_30);
    
    \reg_H1[26]\ : SLE
      port map(D => \N1_data[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[26]\);
    
    next_reg_H7_cry_2_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[2]\, B => 
        hash_control_st_reg_i(6), C => R7_data(2), D => GND_net_1, 
        FCI => next_reg_H7_cry_1, S => \N7_data[2]\, Y => OPEN, 
        FCO => next_reg_H7_cry_2);
    
    next_reg_H3_cry_2_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[2]\, B => 
        hash_control_st_reg_i(6), C => R3_data(2), D => GND_net_1, 
        FCI => next_reg_H3_cry_1, S => \N3_data[2]\, Y => OPEN, 
        FCO => next_reg_H3_cry_2);
    
    next_reg_H0_cry_6_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[6]\, B => 
        hash_control_st_reg_i(6), C => R0_data(6), D => GND_net_1, 
        FCI => next_reg_H0_cry_5, S => \N0_data[6]\, Y => OPEN, 
        FCO => next_reg_H0_cry_6);
    
    next_reg_H7_cry_18_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[18]\, B => 
        hash_control_st_reg_i(6), C => R7_data(18), D => 
        GND_net_1, FCI => next_reg_H7_cry_17, S => \N7_data[18]\, 
        Y => OPEN, FCO => next_reg_H7_cry_18);
    
    next_reg_H6_cry_11_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[11]\, B => 
        hash_control_st_reg_i(6), C => R6_data(11), D => 
        GND_net_1, FCI => next_reg_H6_cry_10, S => \N6_data[11]\, 
        Y => OPEN, FCO => next_reg_H6_cry_11);
    
    next_reg_H3_cry_9_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[9]\, B => 
        hash_control_st_reg_i(6), C => R3_data(9), D => GND_net_1, 
        FCI => next_reg_H3_cry_8, S => \N3_data[9]\, Y => OPEN, 
        FCO => next_reg_H3_cry_9);
    
    \reg_H5[13]\ : SLE
      port map(D => \N5_data[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[13]\);
    
    \reg_H0[1]\ : SLE
      port map(D => \N0_data[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[1]\);
    
    \reg_H5[14]\ : SLE
      port map(D => \N5_data[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[14]\);
    
    \reg_H4[2]\ : SLE
      port map(D => \N4_data[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[2]\);
    
    next_reg_H2_cry_25_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[25]\, B => 
        hash_control_st_reg_i(6), C => R2_data(25), D => 
        GND_net_1, FCI => next_reg_H2_cry_24, S => \N2_data[25]\, 
        Y => OPEN, FCO => next_reg_H2_cry_25);
    
    \reg_H3[8]\ : SLE
      port map(D => \N3_data[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[8]\);
    
    \reg_H6[29]\ : SLE
      port map(D => \N6_data[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[29]\);
    
    \reg_H5[23]\ : SLE
      port map(D => \N5_data[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[23]\);
    
    \reg_H0[12]\ : SLE
      port map(D => \N0_data[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[12]\);
    
    \reg_H5[24]\ : SLE
      port map(D => \N5_data[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[24]\);
    
    next_reg_H5_cry_2_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[2]\, B => 
        hash_control_st_reg_i(6), C => R5_data(2), D => GND_net_1, 
        FCI => next_reg_H5_cry_1, S => \N5_data[2]\, Y => OPEN, 
        FCO => next_reg_H5_cry_2);
    
    next_reg_H0_cry_26_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[26]\, B => 
        hash_control_st_reg_i(6), C => R0_data(26), D => 
        GND_net_1, FCI => next_reg_H0_cry_25, S => \N0_data[26]\, 
        Y => OPEN, FCO => next_reg_H0_cry_26);
    
    next_reg_H0_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[15]\, B => 
        hash_control_st_reg_i(6), C => R0_data(15), D => 
        GND_net_1, FCI => next_reg_H0_cry_14, S => \N0_data[15]\, 
        Y => OPEN, FCO => next_reg_H0_cry_15);
    
    \reg_H7[18]\ : SLE
      port map(D => \N7_data[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[18]\);
    
    \reg_H0[17]\ : SLE
      port map(D => \N0_data[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[17]\);
    
    next_reg_H1_cry_30_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[30]\, B => 
        hash_control_st_reg_i(6), C => R1_data(30), D => 
        GND_net_1, FCI => next_reg_H1_cry_29, S => \N1_data[30]\, 
        Y => OPEN, FCO => next_reg_H1_cry_30);
    
    next_reg_H1_cry_17_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[17]\, B => 
        hash_control_st_reg_i(6), C => R1_data(17), D => 
        GND_net_1, FCI => next_reg_H1_cry_16, S => \N1_data[17]\, 
        Y => OPEN, FCO => next_reg_H1_cry_17);
    
    \reg_H1[1]\ : SLE
      port map(D => \N1_data[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[1]\);
    
    \reg_H1[18]\ : SLE
      port map(D => \N1_data[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[18]\);
    
    next_reg_H5_cry_18_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[18]\, B => 
        hash_control_st_reg_i(6), C => R5_data(18), D => 
        GND_net_1, FCI => next_reg_H5_cry_17, S => \N5_data[18]\, 
        Y => OPEN, FCO => next_reg_H5_cry_18);
    
    next_reg_H3_cry_22_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[22]\, B => 
        hash_control_st_reg_i(6), C => R3_data(22), D => 
        GND_net_1, FCI => next_reg_H3_cry_21, S => \N3_data[22]\, 
        Y => OPEN, FCO => next_reg_H3_cry_22);
    
    next_reg_H7_cry_3_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[3]\, B => 
        hash_control_st_reg_i(6), C => R7_data(3), D => GND_net_1, 
        FCI => next_reg_H7_cry_2, S => \N7_data[3]\, Y => OPEN, 
        FCO => next_reg_H7_cry_3);
    
    next_reg_H3_cry_8_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[8]\, B => 
        hash_control_st_reg_i(6), C => R3_data(8), D => GND_net_1, 
        FCI => next_reg_H3_cry_7, S => \N3_data[8]\, Y => OPEN, 
        FCO => next_reg_H3_cry_8);
    
    next_reg_H3_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[15]\, B => 
        hash_control_st_reg_i(6), C => R3_data(15), D => 
        GND_net_1, FCI => next_reg_H3_cry_14, S => \N3_data[15]\, 
        Y => OPEN, FCO => next_reg_H3_cry_15);
    
    \reg_H0[29]\ : SLE
      port map(D => \N0_data[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[29]\);
    
    next_reg_H4_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[23]\, B => 
        hash_control_st_reg_i(6), C => R4_data(23), D => 
        GND_net_1, FCI => next_reg_H4_cry_22, S => \N4_data[23]\, 
        Y => OPEN, FCO => next_reg_H4_cry_23);
    
    next_reg_H3_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[20]\, B => 
        hash_control_st_reg_i(6), C => R3_data(20), D => 
        GND_net_1, FCI => next_reg_H3_cry_19, S => \N3_data[20]\, 
        Y => OPEN, FCO => next_reg_H3_cry_20);
    
    next_reg_H7_cry_11_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[11]\, B => 
        hash_control_st_reg_i(6), C => R7_data(11), D => 
        GND_net_1, FCI => next_reg_H7_cry_10, S => \N7_data[11]\, 
        Y => OPEN, FCO => next_reg_H7_cry_11);
    
    next_reg_H6_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[28]\, B => 
        hash_control_st_reg_i(6), C => R6_data(28), D => 
        GND_net_1, FCI => next_reg_H6_cry_27, S => \N6_data[28]\, 
        Y => OPEN, FCO => next_reg_H6_cry_28);
    
    \reg_H4[30]\ : SLE
      port map(D => \N4_data[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[30]\);
    
    next_reg_H6_cry_7_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[7]\, B => 
        hash_control_st_reg_i(6), C => R6_data(7), D => GND_net_1, 
        FCI => next_reg_H6_cry_6, S => \N6_data[7]\, Y => OPEN, 
        FCO => next_reg_H6_cry_7);
    
    \reg_H2[23]\ : SLE
      port map(D => \N2_data[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[23]\);
    
    next_reg_H7_cry_26_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[26]\, B => 
        hash_control_st_reg_i(6), C => R7_data(26), D => 
        GND_net_1, FCI => next_reg_H7_cry_25, S => \N7_data[26]\, 
        Y => OPEN, FCO => next_reg_H7_cry_26);
    
    \reg_H2[24]\ : SLE
      port map(D => \N2_data[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[24]\);
    
    \reg_H7[21]\ : SLE
      port map(D => \N7_data[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[21]\);
    
    next_reg_H5_cry_26_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[26]\, B => 
        hash_control_st_reg_i(6), C => R5_data(26), D => 
        GND_net_1, FCI => next_reg_H5_cry_25, S => \N5_data[26]\, 
        Y => OPEN, FCO => next_reg_H5_cry_26);
    
    \reg_H7[15]\ : SLE
      port map(D => \N7_data[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[15]\);
    
    next_reg_H4_cry_17_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[17]\, B => 
        hash_control_st_reg_i(6), C => R4_data(17), D => 
        GND_net_1, FCI => next_reg_H4_cry_16, S => \N4_data[17]\, 
        Y => OPEN, FCO => next_reg_H4_cry_17);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \reg_H5[9]\ : SLE
      port map(D => \N5_data[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[9]\);
    
    \reg_H1[15]\ : SLE
      port map(D => \N1_data[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[15]\);
    
    \reg_H6[9]\ : SLE
      port map(D => \N6_data[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[9]\);
    
    \reg_H6[8]\ : SLE
      port map(D => \N6_data[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[8]\);
    
    \reg_H5[0]\ : SLE
      port map(D => \next_reg_H5_cry_0_0_Y\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[0]\);
    
    \reg_H3[3]\ : SLE
      port map(D => \N3_data[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[3]\);
    
    \reg_H2[18]\ : SLE
      port map(D => \N2_data[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[18]\);
    
    \reg_H1[22]\ : SLE
      port map(D => \N1_data[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[22]\);
    
    \reg_H6[2]\ : SLE
      port map(D => \N6_data[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[2]\);
    
    \reg_H6[18]\ : SLE
      port map(D => \N6_data[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[18]\);
    
    next_reg_H5_cry_3_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[3]\, B => 
        hash_control_st_reg_i(6), C => R5_data(3), D => GND_net_1, 
        FCI => next_reg_H5_cry_2, S => \N5_data[3]\, Y => OPEN, 
        FCO => next_reg_H5_cry_3);
    
    next_reg_H0_cry_29_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[29]\, B => 
        hash_control_st_reg_i(6), C => R0_data(29), D => 
        GND_net_1, FCI => next_reg_H0_cry_28, S => \N0_data[29]\, 
        Y => OPEN, FCO => next_reg_H0_cry_29);
    
    \reg_H0[2]\ : SLE
      port map(D => \N0_data[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[2]\);
    
    next_reg_H5_cry_11_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[11]\, B => 
        hash_control_st_reg_i(6), C => R5_data(11), D => 
        GND_net_1, FCI => next_reg_H5_cry_10, S => \N5_data[11]\, 
        Y => OPEN, FCO => next_reg_H5_cry_11);
    
    \reg_H3[0]\ : SLE
      port map(D => \next_reg_H3_cry_0_0_Y\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[0]\);
    
    \reg_H1[27]\ : SLE
      port map(D => \N1_data[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[27]\);
    
    next_reg_H0_cry_30_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[30]\, B => 
        hash_control_st_reg_i(6), C => R0_data(30), D => 
        GND_net_1, FCI => next_reg_H0_cry_29, S => \N0_data[30]\, 
        Y => OPEN, FCO => next_reg_H0_cry_30);
    
    \reg_H4[28]\ : SLE
      port map(D => \N4_data[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[28]\);
    
    next_reg_H1_cry_14_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[14]\, B => 
        hash_control_st_reg_i(6), C => R1_data(14), D => 
        GND_net_1, FCI => next_reg_H1_cry_13, S => \N1_data[14]\, 
        Y => OPEN, FCO => next_reg_H1_cry_14);
    
    \reg_H0[13]\ : SLE
      port map(D => \N0_data[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[13]\);
    
    \reg_H0[14]\ : SLE
      port map(D => \N0_data[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[14]\);
    
    next_reg_H2_cry_2_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[2]\, B => 
        hash_control_st_reg_i(6), C => R2_data(2), D => GND_net_1, 
        FCI => next_reg_H2_cry_1, S => \N2_data[2]\, Y => OPEN, 
        FCO => next_reg_H2_cry_2);
    
    \reg_H7[26]\ : SLE
      port map(D => \N7_data[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[26]\);
    
    next_reg_H6_cry_21_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[21]\, B => 
        hash_control_st_reg_i(6), C => R6_data(21), D => 
        GND_net_1, FCI => next_reg_H6_cry_20, S => \N6_data[21]\, 
        Y => OPEN, FCO => next_reg_H6_cry_21);
    
    next_reg_H2_cry_16_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[16]\, B => 
        hash_control_st_reg_i(6), C => R2_data(16), D => 
        GND_net_1, FCI => next_reg_H2_cry_15, S => \N2_data[16]\, 
        Y => OPEN, FCO => next_reg_H2_cry_16);
    
    next_reg_H6_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[15]\, B => 
        hash_control_st_reg_i(6), C => R6_data(15), D => 
        GND_net_1, FCI => next_reg_H6_cry_14, S => \N6_data[15]\, 
        Y => OPEN, FCO => next_reg_H6_cry_15);
    
    \reg_H4[10]\ : SLE
      port map(D => \N4_data[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[10]\);
    
    \reg_H0[8]\ : SLE
      port map(D => \N0_data[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[8]\);
    
    \reg_H7[4]\ : SLE
      port map(D => \N7_data[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[4]\);
    
    \reg_H2[15]\ : SLE
      port map(D => \N2_data[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[15]\);
    
    \reg_H6[15]\ : SLE
      port map(D => \N6_data[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[15]\);
    
    next_reg_H7_cry_29_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[29]\, B => 
        hash_control_st_reg_i(6), C => R7_data(29), D => 
        GND_net_1, FCI => next_reg_H7_cry_28, S => \N7_data[29]\, 
        Y => OPEN, FCO => next_reg_H7_cry_29);
    
    next_reg_H1_cry_26_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[26]\, B => 
        hash_control_st_reg_i(6), C => R1_data(26), D => 
        GND_net_1, FCI => next_reg_H1_cry_25, S => \N1_data[26]\, 
        Y => OPEN, FCO => next_reg_H1_cry_26);
    
    next_reg_H5_cry_29_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[29]\, B => 
        hash_control_st_reg_i(6), C => R5_data(29), D => 
        GND_net_1, FCI => next_reg_H5_cry_28, S => \N5_data[29]\, 
        Y => OPEN, FCO => next_reg_H5_cry_29);
    
    next_reg_H1_s_31 : ARI1
      generic map(INIT => x"47D00")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R1_data(31), D => \SHA256_BLOCK_0_H1_o[31]\, FCI => 
        next_reg_H1_cry_30, S => \N1_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    \reg_H4[25]\ : SLE
      port map(D => \N4_data[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[25]\);
    
    next_reg_H4_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[14]\, B => 
        hash_control_st_reg_i(6), C => R4_data(14), D => 
        GND_net_1, FCI => next_reg_H4_cry_13, S => \N4_data[14]\, 
        Y => OPEN, FCO => next_reg_H4_cry_14);
    
    next_reg_H0_cry_5_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[5]\, B => 
        hash_control_st_reg_i(6), C => R0_data(5), D => GND_net_1, 
        FCI => next_reg_H0_cry_4, S => \N0_data[5]\, Y => OPEN, 
        FCO => next_reg_H0_cry_5);
    
    next_reg_H2_cry_5_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[5]\, B => 
        hash_control_st_reg_i(6), C => R2_data(5), D => GND_net_1, 
        FCI => next_reg_H2_cry_4, S => \N2_data[5]\, Y => OPEN, 
        FCO => next_reg_H2_cry_5);
    
    \reg_H2[0]\ : SLE
      port map(D => \next_reg_H2_cry_0_0_Y\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[0]\);
    
    \reg_H7[11]\ : SLE
      port map(D => \N7_data[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[11]\);
    
    next_reg_H6_cry_8_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[8]\, B => 
        hash_control_st_reg_i(6), C => R6_data(8), D => GND_net_1, 
        FCI => next_reg_H6_cry_7, S => \N6_data[8]\, Y => OPEN, 
        FCO => next_reg_H6_cry_8);
    
    next_reg_H4_cry_27_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[27]\, B => 
        hash_control_st_reg_i(6), C => R4_data(27), D => 
        GND_net_1, FCI => next_reg_H4_cry_26, S => \N4_data[27]\, 
        Y => OPEN, FCO => next_reg_H4_cry_27);
    
    \reg_H4[0]\ : SLE
      port map(D => \next_reg_H4_cry_0_0_Y\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[0]\);
    
    \reg_H1[11]\ : SLE
      port map(D => \N1_data[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[11]\);
    
    \reg_H6[31]\ : SLE
      port map(D => \N6_data[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[31]\);
    
    \reg_H5[10]\ : SLE
      port map(D => \N5_data[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[10]\);
    
    \reg_H6[1]\ : SLE
      port map(D => \N6_data[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[1]\);
    
    \reg_H2[30]\ : SLE
      port map(D => \N2_data[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[30]\);
    
    next_reg_H6_cry_2_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[2]\, B => 
        hash_control_st_reg_i(6), C => R6_data(2), D => GND_net_1, 
        FCI => next_reg_H6_cry_1, S => \N6_data[2]\, Y => OPEN, 
        FCO => next_reg_H6_cry_2);
    
    next_reg_H2_cry_26_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[26]\, B => 
        hash_control_st_reg_i(6), C => R2_data(26), D => 
        GND_net_1, FCI => next_reg_H2_cry_25, S => \N2_data[26]\, 
        Y => OPEN, FCO => next_reg_H2_cry_26);
    
    \reg_H7[7]\ : SLE
      port map(D => \N7_data[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[7]\);
    
    \reg_H0[31]\ : SLE
      port map(D => \N0_data[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[31]\);
    
    \reg_H1[23]\ : SLE
      port map(D => \N1_data[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[23]\);
    
    \reg_H1[24]\ : SLE
      port map(D => \N1_data[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[24]\);
    
    next_reg_H7_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[15]\, B => 
        hash_control_st_reg_i(6), C => R7_data(15), D => 
        GND_net_1, FCI => next_reg_H7_cry_14, S => \N7_data[15]\, 
        Y => OPEN, FCO => next_reg_H7_cry_15);
    
    \reg_H5[20]\ : SLE
      port map(D => \N5_data[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[20]\);
    
    \reg_H4[8]\ : SLE
      port map(D => \N4_data[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[8]\);
    
    next_reg_H2_cry_19_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[19]\, B => 
        hash_control_st_reg_i(6), C => R2_data(19), D => 
        GND_net_1, FCI => next_reg_H2_cry_18, S => \N2_data[19]\, 
        Y => OPEN, FCO => next_reg_H2_cry_19);
    
    \reg_H7[5]\ : SLE
      port map(D => \N7_data[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[5]\);
    
    next_reg_H0_cry_16_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[16]\, B => 
        hash_control_st_reg_i(6), C => R0_data(16), D => 
        GND_net_1, FCI => next_reg_H0_cry_15, S => \N0_data[16]\, 
        Y => OPEN, FCO => next_reg_H0_cry_16);
    
    \reg_H4[19]\ : SLE
      port map(D => \N4_data[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[19]\);
    
    \reg_H0[4]\ : SLE
      port map(D => \N0_data[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[4]\);
    
    next_reg_H5_cry_0_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[0]\, B => 
        hash_control_st_reg_i(6), C => R5_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H5_cry_0_0_Y\, 
        FCO => next_reg_H5_cry_0);
    
    next_reg_H1_cry_6_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[6]\, B => 
        hash_control_st_reg_i(6), C => R1_data(6), D => GND_net_1, 
        FCI => next_reg_H1_cry_5, S => \N1_data[6]\, Y => OPEN, 
        FCO => next_reg_H1_cry_6);
    
    next_reg_H1_cry_1_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[1]\, B => 
        hash_control_st_reg_i(6), C => R1_data(1), D => GND_net_1, 
        FCI => next_reg_H1_cry_0, S => \N1_data[1]\, Y => OPEN, 
        FCO => next_reg_H1_cry_1);
    
    \reg_H7[16]\ : SLE
      port map(D => \N7_data[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[16]\);
    
    next_reg_H3_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[23]\, B => 
        hash_control_st_reg_i(6), C => R3_data(23), D => 
        GND_net_1, FCI => next_reg_H3_cry_22, S => \N3_data[23]\, 
        Y => OPEN, FCO => next_reg_H3_cry_23);
    
    \reg_H1[16]\ : SLE
      port map(D => \N1_data[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[16]\);
    
    next_reg_H3_cry_6_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[6]\, B => 
        hash_control_st_reg_i(6), C => R3_data(6), D => GND_net_1, 
        FCI => next_reg_H3_cry_5, S => \N3_data[6]\, Y => OPEN, 
        FCO => next_reg_H3_cry_6);
    
    next_reg_H1_cry_29_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[29]\, B => 
        hash_control_st_reg_i(6), C => R1_data(29), D => 
        GND_net_1, FCI => next_reg_H1_cry_28, S => \N1_data[29]\, 
        Y => OPEN, FCO => next_reg_H1_cry_29);
    
    next_reg_H0_cry_22_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[22]\, B => 
        hash_control_st_reg_i(6), C => R0_data(22), D => 
        GND_net_1, FCI => next_reg_H0_cry_21, S => \N0_data[22]\, 
        Y => OPEN, FCO => next_reg_H0_cry_22);
    
    next_reg_H3_cry_16_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[16]\, B => 
        hash_control_st_reg_i(6), C => R3_data(16), D => 
        GND_net_1, FCI => next_reg_H3_cry_15, S => \N3_data[16]\, 
        Y => OPEN, FCO => next_reg_H3_cry_16);
    
    \reg_H2[11]\ : SLE
      port map(D => \N2_data[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[11]\);
    
    \reg_H6[3]\ : SLE
      port map(D => \N6_data[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[3]\);
    
    \reg_H6[11]\ : SLE
      port map(D => \N6_data[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[11]\);
    
    next_reg_H1_cry_18_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[18]\, B => 
        hash_control_st_reg_i(6), C => R1_data(18), D => 
        GND_net_1, FCI => next_reg_H1_cry_17, S => \N1_data[18]\, 
        Y => OPEN, FCO => next_reg_H1_cry_18);
    
    next_reg_H0_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[20]\, B => 
        hash_control_st_reg_i(6), C => R0_data(20), D => 
        GND_net_1, FCI => next_reg_H0_cry_19, S => \N0_data[20]\, 
        Y => OPEN, FCO => next_reg_H0_cry_20);
    
    \reg_H7[22]\ : SLE
      port map(D => \N7_data[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[22]\);
    
    \reg_H3[7]\ : SLE
      port map(D => \N3_data[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[7]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \reg_H2[20]\ : SLE
      port map(D => \N2_data[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[20]\);
    
    next_reg_H5_cry_15_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[15]\, B => 
        hash_control_st_reg_i(6), C => R5_data(15), D => 
        GND_net_1, FCI => next_reg_H5_cry_14, S => \N5_data[15]\, 
        Y => OPEN, FCO => next_reg_H5_cry_15);
    
    \reg_H4[21]\ : SLE
      port map(D => \N4_data[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[21]\);
    
    next_reg_H4_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[24]\, B => 
        hash_control_st_reg_i(6), C => R4_data(24), D => 
        GND_net_1, FCI => next_reg_H4_cry_23, S => \N4_data[24]\, 
        Y => OPEN, FCO => next_reg_H4_cry_24);
    
    \reg_H7[27]\ : SLE
      port map(D => \N7_data[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[27]\);
    
    \reg_H5[19]\ : SLE
      port map(D => \N5_data[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[19]\);
    
    next_reg_H1_cry_2_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[2]\, B => 
        hash_control_st_reg_i(6), C => R1_data(2), D => GND_net_1, 
        FCI => next_reg_H1_cry_1, S => \N1_data[2]\, Y => OPEN, 
        FCO => next_reg_H1_cry_2);
    
    \reg_H1[31]\ : SLE
      port map(D => \N1_data[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[31]\);
    
    next_reg_H2_cry_29_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[29]\, B => 
        hash_control_st_reg_i(6), C => R2_data(29), D => 
        GND_net_1, FCI => next_reg_H2_cry_28, S => \N2_data[29]\, 
        Y => OPEN, FCO => next_reg_H2_cry_29);
    
    next_reg_H6_cry_25_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[25]\, B => 
        hash_control_st_reg_i(6), C => R6_data(25), D => 
        GND_net_1, FCI => next_reg_H6_cry_24, S => \N6_data[25]\, 
        Y => OPEN, FCO => next_reg_H6_cry_25);
    
    \reg_H3[18]\ : SLE
      port map(D => \N3_data[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[18]\);
    
    next_reg_H7_cry_22_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[22]\, B => 
        hash_control_st_reg_i(6), C => R7_data(22), D => 
        GND_net_1, FCI => next_reg_H7_cry_21, S => \N7_data[22]\, 
        Y => OPEN, FCO => next_reg_H7_cry_22);
    
    next_reg_H2_cry_4_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[4]\, B => 
        hash_control_st_reg_i(6), C => R2_data(4), D => GND_net_1, 
        FCI => next_reg_H2_cry_3, S => \N2_data[4]\, Y => OPEN, 
        FCO => next_reg_H2_cry_4);
    
    \reg_H5[29]\ : SLE
      port map(D => \N5_data[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[29]\);
    
    next_reg_H5_cry_22_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[22]\, B => 
        hash_control_st_reg_i(6), C => R5_data(22), D => 
        GND_net_1, FCI => next_reg_H5_cry_21, S => \N5_data[22]\, 
        Y => OPEN, FCO => next_reg_H5_cry_22);
    
    next_reg_H3_cry_5_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[5]\, B => 
        hash_control_st_reg_i(6), C => R3_data(5), D => GND_net_1, 
        FCI => next_reg_H3_cry_4, S => \N3_data[5]\, Y => OPEN, 
        FCO => next_reg_H3_cry_5);
    
    next_reg_H7_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[20]\, B => 
        hash_control_st_reg_i(6), C => R7_data(20), D => 
        GND_net_1, FCI => next_reg_H7_cry_19, S => \N7_data[20]\, 
        Y => OPEN, FCO => next_reg_H7_cry_20);
    
    next_reg_H4_cry_18_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[18]\, B => 
        hash_control_st_reg_i(6), C => R4_data(18), D => 
        GND_net_1, FCI => next_reg_H4_cry_17, S => \N4_data[18]\, 
        Y => OPEN, FCO => next_reg_H4_cry_18);
    
    next_reg_H0_cry_4_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[4]\, B => 
        hash_control_st_reg_i(6), C => R0_data(4), D => GND_net_1, 
        FCI => next_reg_H0_cry_3, S => \N0_data[4]\, Y => OPEN, 
        FCO => next_reg_H0_cry_4);
    
    \reg_H1[3]\ : SLE
      port map(D => \N1_data[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[3]\);
    
    next_reg_H7_cry_5_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[5]\, B => 
        hash_control_st_reg_i(6), C => R7_data(5), D => GND_net_1, 
        FCI => next_reg_H7_cry_4, S => \N7_data[5]\, Y => OPEN, 
        FCO => next_reg_H7_cry_5);
    
    \reg_H5[6]\ : SLE
      port map(D => \N5_data[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[6]\);
    
    next_reg_H5_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[20]\, B => 
        hash_control_st_reg_i(6), C => R5_data(20), D => 
        GND_net_1, FCI => next_reg_H5_cry_19, S => \N5_data[20]\, 
        Y => OPEN, FCO => next_reg_H5_cry_20);
    
    \reg_H2[16]\ : SLE
      port map(D => \N2_data[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[16]\);
    
    next_reg_H4_cry_9_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[9]\, B => 
        hash_control_st_reg_i(6), C => R4_data(9), D => GND_net_1, 
        FCI => next_reg_H4_cry_8, S => \N4_data[9]\, Y => OPEN, 
        FCO => next_reg_H4_cry_9);
    
    next_reg_H0_cry_19_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[19]\, B => 
        hash_control_st_reg_i(6), C => R0_data(19), D => 
        GND_net_1, FCI => next_reg_H0_cry_18, S => \N0_data[19]\, 
        Y => OPEN, FCO => next_reg_H0_cry_19);
    
    \reg_H6[16]\ : SLE
      port map(D => \N6_data[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[16]\);
    
    \reg_H1[6]\ : SLE
      port map(D => \N1_data[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[6]\);
    
    \reg_H0[10]\ : SLE
      port map(D => \N0_data[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[10]\);
    
    next_reg_H2_cry_9_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[9]\, B => 
        hash_control_st_reg_i(6), C => R2_data(9), D => GND_net_1, 
        FCI => next_reg_H2_cry_8, S => \N2_data[9]\, Y => OPEN, 
        FCO => next_reg_H2_cry_9);
    
    \reg_H7[30]\ : SLE
      port map(D => \N7_data[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[30]\);
    
    \reg_H6[4]\ : SLE
      port map(D => \N6_data[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[4]\);
    
    \reg_H4[26]\ : SLE
      port map(D => \N4_data[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[26]\);
    
    next_reg_H7_s_31 : ARI1
      generic map(INIT => x"42800")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R7_data(31), D => \SHA256_BLOCK_0_H7_o[31]\, FCI => 
        next_reg_H7_cry_30, S => \N7_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_H1_cry_11_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[11]\, B => 
        hash_control_st_reg_i(6), C => R1_data(11), D => 
        GND_net_1, FCI => next_reg_H1_cry_10, S => \N1_data[11]\, 
        Y => OPEN, FCO => next_reg_H1_cry_11);
    
    \reg_H4[5]\ : SLE
      port map(D => \N4_data[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[5]\);
    
    \reg_H3[15]\ : SLE
      port map(D => \N3_data[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[15]\);
    
    next_reg_H5_cry_8_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[8]\, B => 
        hash_control_st_reg_i(6), C => R5_data(8), D => GND_net_1, 
        FCI => next_reg_H5_cry_7, S => \N5_data[8]\, Y => OPEN, 
        FCO => next_reg_H5_cry_8);
    
    next_reg_H3_cry_19_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[19]\, B => 
        hash_control_st_reg_i(6), C => R3_data(19), D => 
        GND_net_1, FCI => next_reg_H3_cry_18, S => \N3_data[19]\, 
        Y => OPEN, FCO => next_reg_H3_cry_19);
    
    next_reg_H6_cry_16_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[16]\, B => 
        hash_control_st_reg_i(6), C => R6_data(16), D => 
        GND_net_1, FCI => next_reg_H6_cry_15, S => \N6_data[16]\, 
        Y => OPEN, FCO => next_reg_H6_cry_16);
    
    \reg_H2[29]\ : SLE
      port map(D => \N2_data[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[29]\);
    
    next_reg_H4_cry_4_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[4]\, B => 
        hash_control_st_reg_i(6), C => R4_data(4), D => GND_net_1, 
        FCI => next_reg_H4_cry_3, S => \N4_data[4]\, Y => OPEN, 
        FCO => next_reg_H4_cry_4);
    
    \reg_H3[6]\ : SLE
      port map(D => \N3_data[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[6]\);
    
    next_reg_H0_cry_7_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[7]\, B => 
        hash_control_st_reg_i(6), C => R0_data(7), D => GND_net_1, 
        FCI => next_reg_H0_cry_6, S => \N0_data[7]\, Y => OPEN, 
        FCO => next_reg_H0_cry_7);
    
    next_reg_H2_cry_8_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[8]\, B => 
        hash_control_st_reg_i(6), C => R2_data(8), D => GND_net_1, 
        FCI => next_reg_H2_cry_7, S => \N2_data[8]\, Y => OPEN, 
        FCO => next_reg_H2_cry_8);
    
    next_reg_H2_cry_12_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[12]\, B => 
        hash_control_st_reg_i(6), C => R2_data(12), D => 
        GND_net_1, FCI => next_reg_H2_cry_11, S => \N2_data[12]\, 
        Y => OPEN, FCO => next_reg_H2_cry_12);
    
    \reg_H7[23]\ : SLE
      port map(D => \N7_data[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[23]\);
    
    \reg_H7[12]\ : SLE
      port map(D => \N7_data[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[12]\);
    
    \reg_H4[1]\ : SLE
      port map(D => \N4_data[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[1]\);
    
    \reg_H0[6]\ : SLE
      port map(D => \N0_data[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[6]\);
    
    \reg_H7[24]\ : SLE
      port map(D => \N7_data[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[24]\);
    
    next_reg_H3_cry_27_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[27]\, B => 
        hash_control_st_reg_i(6), C => R3_data(27), D => 
        GND_net_1, FCI => next_reg_H3_cry_26, S => \N3_data[27]\, 
        Y => OPEN, FCO => next_reg_H3_cry_27);
    
    \reg_H1[12]\ : SLE
      port map(D => \N1_data[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[12]\);
    
    next_reg_H2_cry_10_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[10]\, B => 
        hash_control_st_reg_i(6), C => R2_data(10), D => 
        GND_net_1, FCI => next_reg_H2_cry_9, S => \N2_data[10]\, 
        Y => OPEN, FCO => next_reg_H2_cry_10);
    
    \reg_H7[17]\ : SLE
      port map(D => \N7_data[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[17]\);
    
    next_reg_H4_cry_11_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[11]\, B => 
        hash_control_st_reg_i(6), C => R4_data(11), D => 
        GND_net_1, FCI => next_reg_H4_cry_10, S => \N4_data[11]\, 
        Y => OPEN, FCO => next_reg_H4_cry_11);
    
    \reg_H1[17]\ : SLE
      port map(D => \N1_data[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[17]\);
    
    next_reg_H1_cry_22_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[22]\, B => 
        hash_control_st_reg_i(6), C => R1_data(22), D => 
        GND_net_1, FCI => next_reg_H1_cry_21, S => \N1_data[22]\, 
        Y => OPEN, FCO => next_reg_H1_cry_22);
    
    next_reg_H1_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[20]\, B => 
        hash_control_st_reg_i(6), C => R1_data(20), D => 
        GND_net_1, FCI => next_reg_H1_cry_19, S => \N1_data[20]\, 
        Y => OPEN, FCO => next_reg_H1_cry_20);
    
    next_reg_H4_cry_0_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[0]\, B => 
        hash_control_st_reg_i(6), C => R4_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H4_cry_0_0_Y\, 
        FCO => next_reg_H4_cry_0);
    
    next_reg_H3_cry_1_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[1]\, B => 
        hash_control_st_reg_i(6), C => R3_data(1), D => GND_net_1, 
        FCI => next_reg_H3_cry_0, S => \N3_data[1]\, Y => OPEN, 
        FCO => next_reg_H3_cry_1);
    
    \reg_H3[2]\ : SLE
      port map(D => \N3_data[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[2]\);
    
    \reg_H0[19]\ : SLE
      port map(D => \N0_data[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[19]\);
    
    next_reg_H4_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[28]\, B => 
        hash_control_st_reg_i(6), C => R4_data(28), D => 
        GND_net_1, FCI => next_reg_H4_cry_27, S => \N4_data[28]\, 
        Y => OPEN, FCO => next_reg_H4_cry_28);
    
    \reg_H1[20]\ : SLE
      port map(D => \N1_data[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[20]\);
    
    \reg_H5[30]\ : SLE
      port map(D => \N5_data[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[30]\);
    
    next_reg_H7_cry_16_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[16]\, B => 
        hash_control_st_reg_i(6), C => R7_data(16), D => 
        GND_net_1, FCI => next_reg_H7_cry_15, S => \N7_data[16]\, 
        Y => OPEN, FCO => next_reg_H7_cry_16);
    
    next_reg_H4_cry_1_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[1]\, B => 
        hash_control_st_reg_i(6), C => R4_data(1), D => GND_net_1, 
        FCI => next_reg_H4_cry_0, S => \N4_data[1]\, Y => OPEN, 
        FCO => next_reg_H4_cry_1);
    
    next_reg_H2_cry_22_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[22]\, B => 
        hash_control_st_reg_i(6), C => R2_data(22), D => 
        GND_net_1, FCI => next_reg_H2_cry_21, S => \N2_data[22]\, 
        Y => OPEN, FCO => next_reg_H2_cry_22);
    
    next_reg_H6_cry_19_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[19]\, B => 
        hash_control_st_reg_i(6), C => R6_data(19), D => 
        GND_net_1, FCI => next_reg_H6_cry_18, S => \N6_data[19]\, 
        Y => OPEN, FCO => next_reg_H6_cry_19);
    
    next_reg_H2_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[20]\, B => 
        hash_control_st_reg_i(6), C => R2_data(20), D => 
        GND_net_1, FCI => next_reg_H2_cry_19, S => \N2_data[20]\, 
        Y => OPEN, FCO => next_reg_H2_cry_20);
    
    \reg_H3[11]\ : SLE
      port map(D => \N3_data[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[11]\);
    
    \reg_H2[12]\ : SLE
      port map(D => \N2_data[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[12]\);
    
    \reg_H6[12]\ : SLE
      port map(D => \N6_data[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[12]\);
    
    next_reg_H0_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[23]\, B => 
        hash_control_st_reg_i(6), C => R0_data(23), D => 
        GND_net_1, FCI => next_reg_H0_cry_22, S => \N0_data[23]\, 
        Y => OPEN, FCO => next_reg_H0_cry_23);
    
    \reg_H2[17]\ : SLE
      port map(D => \N2_data[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[17]\);
    
    next_reg_H0_cry_12_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[12]\, B => 
        hash_control_st_reg_i(6), C => R0_data(12), D => 
        GND_net_1, FCI => next_reg_H0_cry_11, S => \N0_data[12]\, 
        Y => OPEN, FCO => next_reg_H0_cry_12);
    
    \reg_H6[17]\ : SLE
      port map(D => \N6_data[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[17]\);
    
    \reg_H4[22]\ : SLE
      port map(D => \N4_data[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[22]\);
    
    \reg_H3[28]\ : SLE
      port map(D => \N3_data[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[28]\);
    
    next_reg_H3_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[24]\, B => 
        hash_control_st_reg_i(6), C => R3_data(24), D => 
        GND_net_1, FCI => next_reg_H3_cry_23, S => \N3_data[24]\, 
        Y => OPEN, FCO => next_reg_H3_cry_24);
    
    next_reg_H0_cry_10_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[10]\, B => 
        hash_control_st_reg_i(6), C => R0_data(10), D => 
        GND_net_1, FCI => next_reg_H0_cry_9, S => \N0_data[10]\, 
        Y => OPEN, FCO => next_reg_H0_cry_10);
    
    next_reg_H5_cry_1_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[1]\, B => 
        hash_control_st_reg_i(6), C => R5_data(1), D => GND_net_1, 
        FCI => next_reg_H5_cry_0, S => \N5_data[1]\, Y => OPEN, 
        FCO => next_reg_H5_cry_1);
    
    \reg_H4[27]\ : SLE
      port map(D => \N4_data[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[27]\);
    
    next_reg_H5_cry_16_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[16]\, B => 
        hash_control_st_reg_i(6), C => R5_data(16), D => 
        GND_net_1, FCI => next_reg_H5_cry_15, S => \N5_data[16]\, 
        Y => OPEN, FCO => next_reg_H5_cry_16);
    
    \reg_H7[13]\ : SLE
      port map(D => \N7_data[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[13]\);
    
    \reg_H7[14]\ : SLE
      port map(D => \N7_data[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[14]\);
    
    \reg_H1[13]\ : SLE
      port map(D => \N1_data[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[13]\);
    
    next_reg_H3_cry_12_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[12]\, B => 
        hash_control_st_reg_i(6), C => R3_data(12), D => 
        GND_net_1, FCI => next_reg_H3_cry_11, S => \N3_data[12]\, 
        Y => OPEN, FCO => next_reg_H3_cry_12);
    
    \reg_H1[14]\ : SLE
      port map(D => \N1_data[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[14]\);
    
    next_reg_H7_cry_8_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[8]\, B => 
        hash_control_st_reg_i(6), C => R7_data(8), D => GND_net_1, 
        FCI => next_reg_H7_cry_7, S => \N7_data[8]\, Y => OPEN, 
        FCO => next_reg_H7_cry_8);
    
    next_reg_H5_cry_4_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[4]\, B => 
        hash_control_st_reg_i(6), C => R5_data(4), D => GND_net_1, 
        FCI => next_reg_H5_cry_3, S => \N5_data[4]\, Y => OPEN, 
        FCO => next_reg_H5_cry_4);
    
    next_reg_H4_cry_21_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[21]\, B => 
        hash_control_st_reg_i(6), C => R4_data(21), D => 
        GND_net_1, FCI => next_reg_H4_cry_20, S => \N4_data[21]\, 
        Y => OPEN, FCO => next_reg_H4_cry_21);
    
    \reg_H1[0]\ : SLE
      port map(D => \next_reg_H1_cry_0_0_Y\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[0]\);
    
    next_reg_H3_cry_10_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[10]\, B => 
        hash_control_st_reg_i(6), C => R3_data(10), D => 
        GND_net_1, FCI => next_reg_H3_cry_9, S => \N3_data[10]\, 
        Y => OPEN, FCO => next_reg_H3_cry_10);
    
    next_reg_H1_cry_15_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[15]\, B => 
        hash_control_st_reg_i(6), C => R1_data(15), D => 
        GND_net_1, FCI => next_reg_H1_cry_14, S => \N1_data[15]\, 
        Y => OPEN, FCO => next_reg_H1_cry_15);
    
    \reg_H1[29]\ : SLE
      port map(D => \N1_data[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[29]\);
    
    next_reg_H7_cry_23_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[23]\, B => 
        hash_control_st_reg_i(6), C => R7_data(23), D => 
        GND_net_1, FCI => next_reg_H7_cry_22, S => \N7_data[23]\, 
        Y => OPEN, FCO => next_reg_H7_cry_23);
    
    next_reg_H6_cry_26_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[26]\, B => 
        hash_control_st_reg_i(6), C => R6_data(26), D => 
        GND_net_1, FCI => next_reg_H6_cry_25, S => \N6_data[26]\, 
        Y => OPEN, FCO => next_reg_H6_cry_26);
    
    \reg_H2[7]\ : SLE
      port map(D => \N2_data[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[7]\);
    
    next_reg_H5_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[23]\, B => 
        hash_control_st_reg_i(6), C => R5_data(23), D => 
        GND_net_1, FCI => next_reg_H5_cry_22, S => \N5_data[23]\, 
        Y => OPEN, FCO => next_reg_H5_cry_23);
    
    \reg_H3[16]\ : SLE
      port map(D => \N3_data[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[16]\);
    
    next_reg_H0_cry_3_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[3]\, B => 
        hash_control_st_reg_i(6), C => R0_data(3), D => GND_net_1, 
        FCI => next_reg_H0_cry_2, S => \N0_data[3]\, Y => OPEN, 
        FCO => next_reg_H0_cry_3);
    
    \reg_H6[28]\ : SLE
      port map(D => \N6_data[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[28]\);
    
    \reg_H3[25]\ : SLE
      port map(D => \N3_data[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[25]\);
    
    next_reg_H7_cry_19_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[19]\, B => 
        hash_control_st_reg_i(6), C => R7_data(19), D => 
        GND_net_1, FCI => next_reg_H7_cry_18, S => \N7_data[19]\, 
        Y => OPEN, FCO => next_reg_H7_cry_19);
    
    \reg_H7[2]\ : SLE
      port map(D => \N7_data[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[2]\);
    
    \reg_H2[1]\ : SLE
      port map(D => \N2_data[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[1]\);
    
    next_reg_H7_cry_9_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[9]\, B => 
        hash_control_st_reg_i(6), C => R7_data(9), D => GND_net_1, 
        FCI => next_reg_H7_cry_8, S => \N7_data[9]\, Y => OPEN, 
        FCO => next_reg_H7_cry_9);
    
    next_reg_H0_cry_0_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[0]\, B => 
        hash_control_st_reg_i(6), C => R0_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H0_cry_0_0_Y\, 
        FCO => next_reg_H0_cry_0);
    
    \reg_H2[8]\ : SLE
      port map(D => \N2_data[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[8]\);
    
    next_reg_H7_cry_0_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[0]\, B => 
        hash_control_st_reg_i(6), C => R7_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H7_cry_0_0_Y\, 
        FCO => next_reg_H7_cry_0);
    
    \reg_H5[7]\ : SLE
      port map(D => \N5_data[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[7]\);
    
    next_reg_H4_cry_15_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[15]\, B => 
        hash_control_st_reg_i(6), C => R4_data(15), D => 
        GND_net_1, FCI => next_reg_H4_cry_14, S => \N4_data[15]\, 
        Y => OPEN, FCO => next_reg_H4_cry_15);
    
    \reg_H3[1]\ : SLE
      port map(D => \N3_data[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[1]\);
    
    \reg_H0[28]\ : SLE
      port map(D => \N0_data[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[28]\);
    
    \reg_H2[13]\ : SLE
      port map(D => \N2_data[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[13]\);
    
    next_reg_H6_cry_9_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[9]\, B => 
        hash_control_st_reg_i(6), C => R6_data(9), D => GND_net_1, 
        FCI => next_reg_H6_cry_8, S => \N6_data[9]\, Y => OPEN, 
        FCO => next_reg_H6_cry_9);
    
    \reg_H6[25]\ : SLE
      port map(D => \N6_data[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[25]\);
    
    \reg_H6[13]\ : SLE
      port map(D => \N6_data[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[13]\);
    
    \reg_H2[14]\ : SLE
      port map(D => \N2_data[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[14]\);
    
    \reg_H6[14]\ : SLE
      port map(D => \N6_data[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[14]\);
    
    next_reg_H4_cry_8_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[8]\, B => 
        hash_control_st_reg_i(6), C => R4_data(8), D => GND_net_1, 
        FCI => next_reg_H4_cry_7, S => \N4_data[8]\, Y => OPEN, 
        FCO => next_reg_H4_cry_8);
    
    next_reg_H5_cry_19_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[19]\, B => 
        hash_control_st_reg_i(6), C => R5_data(19), D => 
        GND_net_1, FCI => next_reg_H5_cry_18, S => \N5_data[19]\, 
        Y => OPEN, FCO => next_reg_H5_cry_19);
    
    \reg_H7[3]\ : SLE
      port map(D => \N7_data[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[3]\);
    
    next_reg_H2_cry_13_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[13]\, B => 
        hash_control_st_reg_i(6), C => R2_data(13), D => 
        GND_net_1, FCI => next_reg_H2_cry_12, S => \N2_data[13]\, 
        Y => OPEN, FCO => next_reg_H2_cry_13);
    
    \reg_H4[23]\ : SLE
      port map(D => \N4_data[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[23]\);
    
    \reg_H7[20]\ : SLE
      port map(D => \N7_data[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[20]\);
    
    \reg_H4[24]\ : SLE
      port map(D => \N4_data[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[24]\);
    
    next_reg_H6_cry_12_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[12]\, B => 
        hash_control_st_reg_i(6), C => R6_data(12), D => 
        GND_net_1, FCI => next_reg_H6_cry_11, S => \N6_data[12]\, 
        Y => OPEN, FCO => next_reg_H6_cry_12);
    
    next_reg_H0_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[27]\, B => 
        hash_control_st_reg_i(6), C => R0_data(27), D => 
        GND_net_1, FCI => next_reg_H0_cry_26, S => \N0_data[27]\, 
        Y => OPEN, FCO => next_reg_H0_cry_27);
    
    next_reg_H6_cry_29_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[29]\, B => 
        hash_control_st_reg_i(6), C => R6_data(29), D => 
        GND_net_1, FCI => next_reg_H6_cry_28, S => \N6_data[29]\, 
        Y => OPEN, FCO => next_reg_H6_cry_29);
    
    next_reg_H6_cry_10_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[10]\, B => 
        hash_control_st_reg_i(6), C => R6_data(10), D => 
        GND_net_1, FCI => next_reg_H6_cry_9, S => \N6_data[10]\, 
        Y => OPEN, FCO => next_reg_H6_cry_10);
    
    next_reg_H1_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[23]\, B => 
        hash_control_st_reg_i(6), C => R1_data(23), D => 
        GND_net_1, FCI => next_reg_H1_cry_22, S => \N1_data[23]\, 
        Y => OPEN, FCO => next_reg_H1_cry_23);
    
    \reg_H5[8]\ : SLE
      port map(D => \N5_data[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[8]\);
    
    \reg_H0[3]\ : SLE
      port map(D => \N0_data[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[3]\);
    
    \reg_H0[25]\ : SLE
      port map(D => \N0_data[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[25]\);
    
    next_reg_H3_cry_28_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[28]\, B => 
        hash_control_st_reg_i(6), C => R3_data(28), D => 
        GND_net_1, FCI => next_reg_H3_cry_27, S => \N3_data[28]\, 
        Y => OPEN, FCO => next_reg_H3_cry_28);
    
    next_reg_H1_cry_9_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[9]\, B => 
        hash_control_st_reg_i(6), C => R1_data(9), D => GND_net_1, 
        FCI => next_reg_H1_cry_8, S => \N1_data[9]\, Y => OPEN, 
        FCO => next_reg_H1_cry_9);
    
    \reg_H3[21]\ : SLE
      port map(D => \N3_data[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[21]\);
    
    next_reg_H1_cry_7_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[7]\, B => 
        hash_control_st_reg_i(6), C => R1_data(7), D => GND_net_1, 
        FCI => next_reg_H1_cry_6, S => \N1_data[7]\, Y => OPEN, 
        FCO => next_reg_H1_cry_7);
    
    \reg_H5[2]\ : SLE
      port map(D => \N5_data[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[2]\);
    
    \reg_H0[0]\ : SLE
      port map(D => \next_reg_H0_cry_0_0_Y\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[0]\);
    
    next_reg_H7_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[27]\, B => 
        hash_control_st_reg_i(6), C => R7_data(27), D => 
        GND_net_1, FCI => next_reg_H7_cry_26, S => \N7_data[27]\, 
        Y => OPEN, FCO => next_reg_H7_cry_27);
    
    next_reg_H2_cry_23_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[23]\, B => 
        hash_control_st_reg_i(6), C => R2_data(23), D => 
        GND_net_1, FCI => next_reg_H2_cry_22, S => \N2_data[23]\, 
        Y => OPEN, FCO => next_reg_H2_cry_23);
    
    \reg_H3[31]\ : SLE
      port map(D => \N3_data[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[31]\);
    
    next_reg_H5_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[27]\, B => 
        hash_control_st_reg_i(6), C => R5_data(27), D => 
        GND_net_1, FCI => next_reg_H5_cry_26, S => \N5_data[27]\, 
        Y => OPEN, FCO => next_reg_H5_cry_27);
    
    \reg_H3[12]\ : SLE
      port map(D => \N3_data[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[12]\);
    
    \reg_H0[9]\ : SLE
      port map(D => \N0_data[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[9]\);
    
    \reg_H6[0]\ : SLE
      port map(D => \next_reg_H6_cry_0_0_Y\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[0]\);
    
    \reg_H0[5]\ : SLE
      port map(D => \N0_data[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[5]\);
    
    next_reg_H4_cry_25_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[25]\, B => 
        hash_control_st_reg_i(6), C => R4_data(25), D => 
        GND_net_1, FCI => next_reg_H4_cry_24, S => \N4_data[25]\, 
        Y => OPEN, FCO => next_reg_H4_cry_25);
    
    \reg_H3[17]\ : SLE
      port map(D => \N3_data[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[17]\);
    
    next_reg_H7_cry_12_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[12]\, B => 
        hash_control_st_reg_i(6), C => R7_data(12), D => 
        GND_net_1, FCI => next_reg_H7_cry_11, S => \N7_data[12]\, 
        Y => OPEN, FCO => next_reg_H7_cry_12);
    
    \reg_H7[29]\ : SLE
      port map(D => \N7_data[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[29]\);
    
    next_reg_H0_cry_13_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[13]\, B => 
        hash_control_st_reg_i(6), C => R0_data(13), D => 
        GND_net_1, FCI => next_reg_H0_cry_12, S => \N0_data[13]\, 
        Y => OPEN, FCO => next_reg_H0_cry_13);
    
    \reg_H6[21]\ : SLE
      port map(D => \N6_data[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[21]\);
    
    next_reg_H7_cry_10_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[10]\, B => 
        hash_control_st_reg_i(6), C => R7_data(10), D => 
        GND_net_1, FCI => next_reg_H7_cry_9, S => \N7_data[10]\, 
        Y => OPEN, FCO => next_reg_H7_cry_10);
    
    \reg_H5[3]\ : SLE
      port map(D => \N5_data[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[3]\);
    
    next_reg_H6_cry_6_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[6]\, B => 
        hash_control_st_reg_i(6), C => R6_data(6), D => GND_net_1, 
        FCI => next_reg_H6_cry_5, S => \N6_data[6]\, Y => OPEN, 
        FCO => next_reg_H6_cry_6);
    
    next_reg_H0_cry_24_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[24]\, B => 
        hash_control_st_reg_i(6), C => R0_data(24), D => 
        GND_net_1, FCI => next_reg_H0_cry_23, S => \N0_data[24]\, 
        Y => OPEN, FCO => next_reg_H0_cry_24);
    
    \reg_H3[26]\ : SLE
      port map(D => \N3_data[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[26]\);
    
    next_reg_H4_cry_3_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[3]\, B => 
        hash_control_st_reg_i(6), C => R4_data(3), D => GND_net_1, 
        FCI => next_reg_H4_cry_2, S => \N4_data[3]\, Y => OPEN, 
        FCO => next_reg_H4_cry_3);
    
    next_reg_H1_cry_0_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[0]\, B => 
        hash_control_st_reg_i(6), C => R1_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H1_cry_0_0_Y\, 
        FCO => next_reg_H1_cry_0);
    
    next_reg_H3_s_31 : ARI1
      generic map(INIT => x"47D00")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R3_data(31), D => \SHA256_BLOCK_0_H3_o[31]\, FCI => 
        next_reg_H3_cry_30, S => \N3_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    \reg_H7[10]\ : SLE
      port map(D => \N7_data[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[10]\);
    
    \reg_H1[9]\ : SLE
      port map(D => \N1_data[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[9]\);
    
    next_reg_H3_cry_21_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[21]\, B => 
        hash_control_st_reg_i(6), C => R3_data(21), D => 
        GND_net_1, FCI => next_reg_H3_cry_20, S => \N3_data[21]\, 
        Y => OPEN, FCO => next_reg_H3_cry_21);
    
    next_reg_H2_cry_7_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[7]\, B => 
        hash_control_st_reg_i(6), C => R2_data(7), D => GND_net_1, 
        FCI => next_reg_H2_cry_6, S => \N2_data[7]\, Y => OPEN, 
        FCO => next_reg_H2_cry_7);
    
    next_reg_H0_cry_8_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[8]\, B => 
        hash_control_st_reg_i(6), C => R0_data(8), D => GND_net_1, 
        FCI => next_reg_H0_cry_7, S => \N0_data[8]\, Y => OPEN, 
        FCO => next_reg_H0_cry_8);
    
    next_reg_H3_cry_13_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[13]\, B => 
        hash_control_st_reg_i(6), C => R3_data(13), D => 
        GND_net_1, FCI => next_reg_H3_cry_12, S => \N3_data[13]\, 
        Y => OPEN, FCO => next_reg_H3_cry_13);
    
    \reg_H1[10]\ : SLE
      port map(D => \N1_data[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[10]\);
    
    \reg_H6[30]\ : SLE
      port map(D => \N6_data[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[30]\);
    
    next_reg_H2_cry_17_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[17]\, B => 
        hash_control_st_reg_i(6), C => R2_data(17), D => 
        GND_net_1, FCI => next_reg_H2_cry_16, S => \N2_data[17]\, 
        Y => OPEN, FCO => next_reg_H2_cry_17);
    
    \reg_H0[21]\ : SLE
      port map(D => \N0_data[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[21]\);
    
    next_reg_H1_cry_16_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[16]\, B => 
        hash_control_st_reg_i(6), C => R1_data(16), D => 
        GND_net_1, FCI => next_reg_H1_cry_15, S => \N1_data[16]\, 
        Y => OPEN, FCO => next_reg_H1_cry_16);
    
    \reg_H0[30]\ : SLE
      port map(D => \N0_data[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[30]\);
    
    \reg_H3[9]\ : SLE
      port map(D => \N3_data[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[9]\);
    
    next_reg_H5_cry_12_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[12]\, B => 
        hash_control_st_reg_i(6), C => R5_data(12), D => 
        GND_net_1, FCI => next_reg_H5_cry_11, S => \N5_data[12]\, 
        Y => OPEN, FCO => next_reg_H5_cry_12);
    
    next_reg_H0_s_31 : ARI1
      generic map(INIT => x"42800")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R0_data(31), D => \SHA256_BLOCK_0_H0_o[31]\, FCI => 
        next_reg_H0_cry_30, S => \N0_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_H5_cry_30_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[30]\, B => 
        hash_control_st_reg_i(6), C => R5_data(30), D => 
        GND_net_1, FCI => next_reg_H5_cry_29, S => \N5_data[30]\, 
        Y => OPEN, FCO => next_reg_H5_cry_30);
    
    next_reg_H5_cry_10_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[10]\, B => 
        hash_control_st_reg_i(6), C => R5_data(10), D => 
        GND_net_1, FCI => next_reg_H5_cry_9, S => \N5_data[10]\, 
        Y => OPEN, FCO => next_reg_H5_cry_10);
    
    next_reg_H7_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[24]\, B => 
        hash_control_st_reg_i(6), C => R7_data(24), D => 
        GND_net_1, FCI => next_reg_H7_cry_23, S => \N7_data[24]\, 
        Y => OPEN, FCO => next_reg_H7_cry_24);
    
    next_reg_H2_cry_1_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[1]\, B => 
        hash_control_st_reg_i(6), C => R2_data(1), D => GND_net_1, 
        FCI => next_reg_H2_cry_0, S => \N2_data[1]\, Y => OPEN, 
        FCO => next_reg_H2_cry_1);
    
    next_reg_H1_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[27]\, B => 
        hash_control_st_reg_i(6), C => R1_data(27), D => 
        GND_net_1, FCI => next_reg_H1_cry_26, S => \N1_data[27]\, 
        Y => OPEN, FCO => next_reg_H1_cry_27);
    
    \reg_H6[26]\ : SLE
      port map(D => \N6_data[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[26]\);
    
    \reg_H2[5]\ : SLE
      port map(D => \N2_data[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[5]\);
    
    next_reg_H5_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[24]\, B => 
        hash_control_st_reg_i(6), C => R5_data(24), D => 
        GND_net_1, FCI => next_reg_H5_cry_23, S => \N5_data[24]\, 
        Y => OPEN, FCO => next_reg_H5_cry_24);
    
    \reg_H7[8]\ : SLE
      port map(D => \N7_data[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[8]\);
    
    \reg_H4[18]\ : SLE
      port map(D => \N4_data[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[18]\);
    
    next_reg_H6_cry_22_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[22]\, B => 
        hash_control_st_reg_i(6), C => R6_data(22), D => 
        GND_net_1, FCI => next_reg_H6_cry_21, S => \N6_data[22]\, 
        Y => OPEN, FCO => next_reg_H6_cry_22);
    
    next_reg_H7_cry_1_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[1]\, B => 
        hash_control_st_reg_i(6), C => R7_data(1), D => GND_net_1, 
        FCI => next_reg_H7_cry_0, S => \N7_data[1]\, Y => OPEN, 
        FCO => next_reg_H7_cry_1);
    
    next_reg_H5_cry_6_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[6]\, B => 
        hash_control_st_reg_i(6), C => R5_data(6), D => GND_net_1, 
        FCI => next_reg_H5_cry_5, S => \N5_data[6]\, Y => OPEN, 
        FCO => next_reg_H5_cry_6);
    
    \reg_H5[5]\ : SLE
      port map(D => \N5_data[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[5]\);
    
    next_reg_H6_cry_20_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[20]\, B => 
        hash_control_st_reg_i(6), C => R6_data(20), D => 
        GND_net_1, FCI => next_reg_H6_cry_19, S => \N6_data[20]\, 
        Y => OPEN, FCO => next_reg_H6_cry_20);
    
    \reg_H3[13]\ : SLE
      port map(D => \N3_data[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[13]\);
    
    next_reg_H3_cry_7_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[7]\, B => 
        hash_control_st_reg_i(6), C => R3_data(7), D => GND_net_1, 
        FCI => next_reg_H3_cry_6, S => \N3_data[7]\, Y => OPEN, 
        FCO => next_reg_H3_cry_7);
    
    \reg_H3[14]\ : SLE
      port map(D => \N3_data[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[14]\);
    
    next_reg_H4_cry_16_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[16]\, B => 
        hash_control_st_reg_i(6), C => R4_data(16), D => 
        GND_net_1, FCI => next_reg_H4_cry_15, S => \N4_data[16]\, 
        Y => OPEN, FCO => next_reg_H4_cry_16);
    
    \reg_H5[4]\ : SLE
      port map(D => \N5_data[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[4]\);
    
    next_reg_H4_cry_7_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[7]\, B => 
        hash_control_st_reg_i(6), C => R4_data(7), D => GND_net_1, 
        FCI => next_reg_H4_cry_6, S => \N4_data[7]\, Y => OPEN, 
        FCO => next_reg_H4_cry_7);
    
    \reg_H2[10]\ : SLE
      port map(D => \N2_data[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[10]\);
    
    next_reg_H7_cry_7_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[7]\, B => 
        hash_control_st_reg_i(6), C => R7_data(7), D => GND_net_1, 
        FCI => next_reg_H7_cry_6, S => \N7_data[7]\, Y => OPEN, 
        FCO => next_reg_H7_cry_7);
    
    \reg_H6[10]\ : SLE
      port map(D => \N6_data[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[10]\);
    
    \reg_H0[26]\ : SLE
      port map(D => \N0_data[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[26]\);
    
    next_reg_H6_cry_0_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[0]\, B => 
        hash_control_st_reg_i(6), C => R6_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H6_cry_0_0_Y\, 
        FCO => next_reg_H6_cry_0);
    
    next_reg_H2_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[27]\, B => 
        hash_control_st_reg_i(6), C => R2_data(27), D => 
        GND_net_1, FCI => next_reg_H2_cry_26, S => \N2_data[27]\, 
        Y => OPEN, FCO => next_reg_H2_cry_27);
    
    \reg_H7[19]\ : SLE
      port map(D => \N7_data[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[19]\);
    
    \reg_H1[19]\ : SLE
      port map(D => \N1_data[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[19]\);
    
    \reg_H6[7]\ : SLE
      port map(D => \N6_data[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[7]\);
    
    \reg_H5[18]\ : SLE
      port map(D => \N5_data[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[18]\);
    
    \reg_H4[20]\ : SLE
      port map(D => \N4_data[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[20]\);
    
    \reg_H4[15]\ : SLE
      port map(D => \N4_data[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[15]\);
    
    next_reg_H6_cry_13_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H6_o[13]\, B => 
        hash_control_st_reg_i(6), C => R6_data(13), D => 
        GND_net_1, FCI => next_reg_H6_cry_12, S => \N6_data[13]\, 
        Y => OPEN, FCO => next_reg_H6_cry_13);
    
    \reg_H1[30]\ : SLE
      port map(D => \N1_data[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[30]\);
    
    next_reg_H2_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[14]\, B => 
        hash_control_st_reg_i(6), C => R2_data(14), D => 
        GND_net_1, FCI => next_reg_H2_cry_13, S => \N2_data[14]\, 
        Y => OPEN, FCO => next_reg_H2_cry_14);
    
    next_reg_H1_cry_19_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[19]\, B => 
        hash_control_st_reg_i(6), C => R1_data(19), D => 
        GND_net_1, FCI => next_reg_H1_cry_18, S => \N1_data[19]\, 
        Y => OPEN, FCO => next_reg_H1_cry_19);
    
    next_reg_H0_cry_17_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[17]\, B => 
        hash_control_st_reg_i(6), C => R0_data(17), D => 
        GND_net_1, FCI => next_reg_H0_cry_16, S => \N0_data[17]\, 
        Y => OPEN, FCO => next_reg_H0_cry_17);
    
    \reg_H4[31]\ : SLE
      port map(D => \N4_data[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[31]\);
    
    \reg_H5[28]\ : SLE
      port map(D => \N5_data[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[28]\);
    
    \reg_H3[22]\ : SLE
      port map(D => \N3_data[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[22]\);
    
    next_reg_H5_cry_5_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[5]\, B => 
        hash_control_st_reg_i(6), C => R5_data(5), D => GND_net_1, 
        FCI => next_reg_H5_cry_4, S => \N5_data[5]\, Y => OPEN, 
        FCO => next_reg_H5_cry_5);
    
    next_reg_H4_cry_2_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[2]\, B => 
        hash_control_st_reg_i(6), C => R4_data(2), D => GND_net_1, 
        FCI => next_reg_H4_cry_1, S => \N4_data[2]\, Y => OPEN, 
        FCO => next_reg_H4_cry_2);
    
    next_reg_H3_cry_0_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[0]\, B => 
        hash_control_st_reg_i(6), C => R3_data(0), D => GND_net_1, 
        FCI => GND_net_1, S => OPEN, Y => \next_reg_H3_cry_0_0_Y\, 
        FCO => next_reg_H3_cry_0);
    
    next_reg_H1_cry_24_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[24]\, B => 
        hash_control_st_reg_i(6), C => R1_data(24), D => 
        GND_net_1, FCI => next_reg_H1_cry_23, S => \N1_data[24]\, 
        Y => OPEN, FCO => next_reg_H1_cry_24);
    
    next_reg_H0_cry_28_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[28]\, B => 
        hash_control_st_reg_i(6), C => R0_data(28), D => 
        GND_net_1, FCI => next_reg_H0_cry_27, S => \N0_data[28]\, 
        Y => OPEN, FCO => next_reg_H0_cry_28);
    
    next_reg_H3_cry_3_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[3]\, B => 
        hash_control_st_reg_i(6), C => R3_data(3), D => GND_net_1, 
        FCI => next_reg_H3_cry_2, S => \N3_data[3]\, Y => OPEN, 
        FCO => next_reg_H3_cry_3);
    
    next_reg_H3_cry_17_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[17]\, B => 
        hash_control_st_reg_i(6), C => R3_data(17), D => 
        GND_net_1, FCI => next_reg_H3_cry_16, S => \N3_data[17]\, 
        Y => OPEN, FCO => next_reg_H3_cry_17);
    
    \reg_H3[27]\ : SLE
      port map(D => \N3_data[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[27]\);
    
    \reg_H5[15]\ : SLE
      port map(D => \N5_data[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[15]\);
    
    next_reg_H2_cry_30_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[30]\, B => 
        hash_control_st_reg_i(6), C => R2_data(30), D => 
        GND_net_1, FCI => next_reg_H2_cry_29, S => \N2_data[30]\, 
        Y => OPEN, FCO => next_reg_H2_cry_30);
    
    next_reg_H4_cry_19_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[19]\, B => 
        hash_control_st_reg_i(6), C => R4_data(19), D => 
        GND_net_1, FCI => next_reg_H4_cry_18, S => \N4_data[19]\, 
        Y => OPEN, FCO => next_reg_H4_cry_19);
    
    \reg_H7[6]\ : SLE
      port map(D => \N7_data[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[6]\);
    
    \reg_H2[19]\ : SLE
      port map(D => \N2_data[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[19]\);
    
    next_reg_H3_cry_25_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[25]\, B => 
        hash_control_st_reg_i(6), C => R3_data(25), D => 
        GND_net_1, FCI => next_reg_H3_cry_24, S => \N3_data[25]\, 
        Y => OPEN, FCO => next_reg_H3_cry_25);
    
    \reg_H6[19]\ : SLE
      port map(D => \N6_data[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[19]\);
    
    next_reg_H4_cry_30_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[30]\, B => 
        hash_control_st_reg_i(6), C => R4_data(30), D => 
        GND_net_1, FCI => next_reg_H4_cry_29, S => \N4_data[30]\, 
        Y => OPEN, FCO => next_reg_H4_cry_30);
    
    \reg_H5[25]\ : SLE
      port map(D => \N5_data[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[25]\);
    
    \reg_H2[28]\ : SLE
      port map(D => \N2_data[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[28]\);
    
    \reg_H6[22]\ : SLE
      port map(D => \N6_data[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[22]\);
    
    next_reg_H7_cry_13_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[13]\, B => 
        hash_control_st_reg_i(6), C => R7_data(13), D => 
        GND_net_1, FCI => next_reg_H7_cry_12, S => \N7_data[13]\, 
        Y => OPEN, FCO => next_reg_H7_cry_13);
    
    next_reg_H4_cry_26_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[26]\, B => 
        hash_control_st_reg_i(6), C => R4_data(26), D => 
        GND_net_1, FCI => next_reg_H4_cry_25, S => \N4_data[26]\, 
        Y => OPEN, FCO => next_reg_H4_cry_26);
    
    next_reg_H2_cry_24_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[24]\, B => 
        hash_control_st_reg_i(6), C => R2_data(24), D => 
        GND_net_1, FCI => next_reg_H2_cry_23, S => \N2_data[24]\, 
        Y => OPEN, FCO => next_reg_H2_cry_24);
    
    \reg_H4[29]\ : SLE
      port map(D => \N4_data[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[29]\);
    
    \reg_H3[5]\ : SLE
      port map(D => \N3_data[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[5]\);
    
    next_reg_H7_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[28]\, B => 
        hash_control_st_reg_i(6), C => R7_data(28), D => 
        GND_net_1, FCI => next_reg_H7_cry_27, S => \N7_data[28]\, 
        Y => OPEN, FCO => next_reg_H7_cry_28);
    
    \reg_H6[27]\ : SLE
      port map(D => \N6_data[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[27]\);
    
    next_reg_H5_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[28]\, B => 
        hash_control_st_reg_i(6), C => R5_data(28), D => 
        GND_net_1, FCI => next_reg_H5_cry_27, S => \N5_data[28]\, 
        Y => OPEN, FCO => next_reg_H5_cry_28);
    
    \reg_H7[9]\ : SLE
      port map(D => \N7_data[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[9]\);
    
    \reg_H1[7]\ : SLE
      port map(D => \N1_data[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[7]\);
    
    \reg_H4[11]\ : SLE
      port map(D => \N4_data[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[11]\);
    
    next_reg_H0_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[14]\, B => 
        hash_control_st_reg_i(6), C => R0_data(14), D => 
        GND_net_1, FCI => next_reg_H0_cry_13, S => \N0_data[14]\, 
        Y => OPEN, FCO => next_reg_H0_cry_14);
    
    next_reg_H4_cry_6_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[6]\, B => 
        hash_control_st_reg_i(6), C => R4_data(6), D => GND_net_1, 
        FCI => next_reg_H4_cry_5, S => \N4_data[6]\, Y => OPEN, 
        FCO => next_reg_H4_cry_6);
    
    next_reg_H0_cry_2_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[2]\, B => 
        hash_control_st_reg_i(6), C => R0_data(2), D => GND_net_1, 
        FCI => next_reg_H0_cry_1, S => \N0_data[2]\, Y => OPEN, 
        FCO => next_reg_H0_cry_2);
    
    next_reg_H0_cry_21_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[21]\, B => 
        hash_control_st_reg_i(6), C => R0_data(21), D => 
        GND_net_1, FCI => next_reg_H0_cry_20, S => \N0_data[21]\, 
        Y => OPEN, FCO => next_reg_H0_cry_21);
    
    \reg_H0[22]\ : SLE
      port map(D => \N0_data[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[22]\);
    
    \reg_H2[25]\ : SLE
      port map(D => \N2_data[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[25]\);
    
    next_reg_H2_s_31 : ARI1
      generic map(INIT => x"42800")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R2_data(31), D => \SHA256_BLOCK_0_H2_o[31]\, FCI => 
        next_reg_H2_cry_30, S => \N2_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_H1_cry_3_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[3]\, B => 
        hash_control_st_reg_i(6), C => R1_data(3), D => GND_net_1, 
        FCI => next_reg_H1_cry_2, S => \N1_data[3]\, Y => OPEN, 
        FCO => next_reg_H1_cry_3);
    
    \reg_H0[27]\ : SLE
      port map(D => \N0_data[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[27]\);
    
    \reg_H0[18]\ : SLE
      port map(D => \N0_data[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[18]\);
    
    next_reg_H5_cry_13_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[13]\, B => 
        hash_control_st_reg_i(6), C => R5_data(13), D => 
        GND_net_1, FCI => next_reg_H5_cry_12, S => \N5_data[13]\, 
        Y => OPEN, FCO => next_reg_H5_cry_13);
    
    next_reg_H3_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[14]\, B => 
        hash_control_st_reg_i(6), C => R3_data(14), D => 
        GND_net_1, FCI => next_reg_H3_cry_13, S => \N3_data[14]\, 
        Y => OPEN, FCO => next_reg_H3_cry_14);
    
    \reg_H5[1]\ : SLE
      port map(D => \N5_data[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[1]\);
    
    next_reg_H6_cry_17_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[17]\, B => 
        hash_control_st_reg_i(6), C => R6_data(17), D => 
        GND_net_1, FCI => next_reg_H6_cry_16, S => \N6_data[17]\, 
        Y => OPEN, FCO => next_reg_H6_cry_17);
    
    \reg_H3[23]\ : SLE
      port map(D => \N3_data[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[23]\);
    
    \reg_H3[24]\ : SLE
      port map(D => \N3_data[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[24]\);
    
    \reg_H5[11]\ : SLE
      port map(D => \N5_data[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[11]\);
    
    \reg_H2[3]\ : SLE
      port map(D => \N2_data[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[3]\);
    
    \reg_H2[31]\ : SLE
      port map(D => \N2_data[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[31]\);
    
    next_reg_H6_cry_23_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[23]\, B => 
        hash_control_st_reg_i(6), C => R6_data(23), D => 
        GND_net_1, FCI => next_reg_H6_cry_22, S => \N6_data[23]\, 
        Y => OPEN, FCO => next_reg_H6_cry_23);
    
    next_reg_H2_cry_18_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[18]\, B => 
        hash_control_st_reg_i(6), C => R2_data(18), D => 
        GND_net_1, FCI => next_reg_H2_cry_17, S => \N2_data[18]\, 
        Y => OPEN, FCO => next_reg_H2_cry_18);
    
    next_reg_H1_cry_12_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[12]\, B => 
        hash_control_st_reg_i(6), C => R1_data(12), D => 
        GND_net_1, FCI => next_reg_H1_cry_11, S => \N1_data[12]\, 
        Y => OPEN, FCO => next_reg_H1_cry_12);
    
    next_reg_H7_cry_21_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H7_o[21]\, B => 
        hash_control_st_reg_i(6), C => R7_data(21), D => 
        GND_net_1, FCI => next_reg_H7_cry_20, S => \N7_data[21]\, 
        Y => OPEN, FCO => next_reg_H7_cry_21);
    
    \reg_H2[4]\ : SLE
      port map(D => \N2_data[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[4]\);
    
    \reg_H4[16]\ : SLE
      port map(D => \N4_data[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[16]\);
    
    next_reg_H5_cry_21_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[21]\, B => 
        hash_control_st_reg_i(6), C => R5_data(21), D => 
        GND_net_1, FCI => next_reg_H5_cry_20, S => \N5_data[21]\, 
        Y => OPEN, FCO => next_reg_H5_cry_21);
    
    next_reg_H4_cry_29_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[29]\, B => 
        hash_control_st_reg_i(6), C => R4_data(29), D => 
        GND_net_1, FCI => next_reg_H4_cry_28, S => \N4_data[29]\, 
        Y => OPEN, FCO => next_reg_H4_cry_29);
    
    next_reg_H1_cry_10_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[10]\, B => 
        hash_control_st_reg_i(6), C => R1_data(10), D => 
        GND_net_1, FCI => next_reg_H1_cry_9, S => \N1_data[10]\, 
        Y => OPEN, FCO => next_reg_H1_cry_10);
    
    \reg_H3[10]\ : SLE
      port map(D => \N3_data[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[10]\);
    
    \reg_H5[21]\ : SLE
      port map(D => \N5_data[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[21]\);
    
    \reg_H4[9]\ : SLE
      port map(D => \N4_data[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[9]\);
    
    next_reg_H1_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[28]\, B => 
        hash_control_st_reg_i(6), C => R1_data(28), D => 
        GND_net_1, FCI => next_reg_H1_cry_27, S => \N1_data[28]\, 
        Y => OPEN, FCO => next_reg_H1_cry_28);
    
    \reg_H0[15]\ : SLE
      port map(D => \N0_data[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[15]\);
    
    \reg_H6[23]\ : SLE
      port map(D => \N6_data[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[23]\);
    
    next_reg_H1_cry_4_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[4]\, B => 
        hash_control_st_reg_i(6), C => R1_data(4), D => GND_net_1, 
        FCI => next_reg_H1_cry_3, S => \N1_data[4]\, Y => OPEN, 
        FCO => next_reg_H1_cry_4);
    
    \reg_H7[1]\ : SLE
      port map(D => \N7_data[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H7_o[1]\);
    
    \reg_H6[24]\ : SLE
      port map(D => \N6_data[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H6_o[24]\);
    
    next_reg_H4_cry_12_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[12]\, B => 
        hash_control_st_reg_i(6), C => R4_data(12), D => 
        GND_net_1, FCI => next_reg_H4_cry_11, S => \N4_data[12]\, 
        Y => OPEN, FCO => next_reg_H4_cry_12);
    
    next_reg_H7_cry_17_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[17]\, B => 
        hash_control_st_reg_i(6), C => R7_data(17), D => 
        GND_net_1, FCI => next_reg_H7_cry_16, S => \N7_data[17]\, 
        Y => OPEN, FCO => next_reg_H7_cry_17);
    
    next_reg_H4_s_31 : ARI1
      generic map(INIT => x"42800")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R4_data(31), D => \SHA256_BLOCK_0_H4_o[31]\, FCI => 
        next_reg_H4_cry_30, S => \N4_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_H3_cry_30_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H3_o[30]\, B => 
        hash_control_st_reg_i(6), C => R3_data(30), D => 
        GND_net_1, FCI => next_reg_H3_cry_29, S => \N3_data[30]\, 
        Y => OPEN, FCO => next_reg_H3_cry_30);
    
    \reg_H5[16]\ : SLE
      port map(D => \N5_data[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[16]\);
    
    \reg_H4[6]\ : SLE
      port map(D => \N4_data[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[6]\);
    
    next_reg_H4_cry_10_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H4_o[10]\, B => 
        hash_control_st_reg_i(6), C => R4_data(10), D => 
        GND_net_1, FCI => next_reg_H4_cry_9, S => \N4_data[10]\, 
        Y => OPEN, FCO => next_reg_H4_cry_10);
    
    next_reg_H2_cry_6_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[6]\, B => 
        hash_control_st_reg_i(6), C => R2_data(6), D => GND_net_1, 
        FCI => next_reg_H2_cry_5, S => \N2_data[6]\, Y => OPEN, 
        FCO => next_reg_H2_cry_6);
    
    next_reg_H2_cry_28_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H2_o[28]\, B => 
        hash_control_st_reg_i(6), C => R2_data(28), D => 
        GND_net_1, FCI => next_reg_H2_cry_27, S => \N2_data[28]\, 
        Y => OPEN, FCO => next_reg_H2_cry_28);
    
    \reg_H2[6]\ : SLE
      port map(D => \N2_data[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[6]\);
    
    \reg_H1[28]\ : SLE
      port map(D => \N1_data[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[28]\);
    
    \reg_H2[2]\ : SLE
      port map(D => \N2_data[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[2]\);
    
    \reg_H0[23]\ : SLE
      port map(D => \N0_data[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[23]\);
    
    next_reg_H6_s_31 : ARI1
      generic map(INIT => x"42800")

      port map(A => VCC_net_1, B => hash_control_st_reg_i(6), C
         => R6_data(31), D => \SHA256_BLOCK_0_H6_o[31]\, FCI => 
        next_reg_H6_cry_30, S => \N6_data[31]\, Y => OPEN, FCO
         => OPEN);
    
    next_reg_H1_cry_5_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H1_o[5]\, B => 
        hash_control_st_reg_i(6), C => R1_data(5), D => GND_net_1, 
        FCI => next_reg_H1_cry_4, S => \N1_data[5]\, Y => OPEN, 
        FCO => next_reg_H1_cry_5);
    
    \reg_H2[21]\ : SLE
      port map(D => \N2_data[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[21]\);
    
    \reg_H0[24]\ : SLE
      port map(D => \N0_data[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[24]\);
    
    next_reg_H6_cry_14_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[14]\, B => 
        hash_control_st_reg_i(6), C => R6_data(14), D => 
        GND_net_1, FCI => next_reg_H6_cry_13, S => \N6_data[14]\, 
        Y => OPEN, FCO => next_reg_H6_cry_14);
    
    next_reg_H6_cry_3_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[3]\, B => 
        hash_control_st_reg_i(6), C => R6_data(3), D => GND_net_1, 
        FCI => next_reg_H6_cry_2, S => \N6_data[3]\, Y => OPEN, 
        FCO => next_reg_H6_cry_3);
    
    next_reg_H2_cry_11_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[11]\, B => 
        hash_control_st_reg_i(6), C => R2_data(11), D => 
        GND_net_1, FCI => next_reg_H2_cry_10, S => \N2_data[11]\, 
        Y => OPEN, FCO => next_reg_H2_cry_11);
    
    next_reg_H4_cry_5_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H4_o[5]\, B => 
        hash_control_st_reg_i(6), C => R4_data(5), D => GND_net_1, 
        FCI => next_reg_H4_cry_4, S => \N4_data[5]\, Y => OPEN, 
        FCO => next_reg_H4_cry_5);
    
    \reg_H5[26]\ : SLE
      port map(D => \N5_data[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H5_o[26]\);
    
    next_reg_H7_cry_6_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H7_o[6]\, B => 
        hash_control_st_reg_i(6), C => R7_data(6), D => GND_net_1, 
        FCI => next_reg_H7_cry_5, S => \N7_data[6]\, Y => OPEN, 
        FCO => next_reg_H7_cry_6);
    
    next_reg_H0_cry_18_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H0_o[18]\, B => 
        hash_control_st_reg_i(6), C => R0_data(18), D => 
        GND_net_1, FCI => next_reg_H0_cry_17, S => \N0_data[18]\, 
        Y => OPEN, FCO => next_reg_H0_cry_18);
    
    next_reg_H1_cry_21_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H1_o[21]\, B => 
        hash_control_st_reg_i(6), C => R1_data(21), D => 
        GND_net_1, FCI => next_reg_H1_cry_20, S => \N1_data[21]\, 
        Y => OPEN, FCO => next_reg_H1_cry_21);
    
    \reg_H4[3]\ : SLE
      port map(D => \N4_data[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H4_o[3]\);
    
    \reg_H3[19]\ : SLE
      port map(D => \N3_data[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H3_o[19]\);
    
    next_reg_H0_cry_1_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[1]\, B => 
        hash_control_st_reg_i(6), C => R0_data(1), D => GND_net_1, 
        FCI => next_reg_H0_cry_0, S => \N0_data[1]\, Y => OPEN, 
        FCO => next_reg_H0_cry_1);
    
    next_reg_H5_cry_7_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H5_o[7]\, B => 
        hash_control_st_reg_i(6), C => R5_data(7), D => GND_net_1, 
        FCI => next_reg_H5_cry_6, S => \N5_data[7]\, Y => OPEN, 
        FCO => next_reg_H5_cry_7);
    
    next_reg_H6_cry_5_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[5]\, B => 
        hash_control_st_reg_i(6), C => R6_data(5), D => GND_net_1, 
        FCI => next_reg_H6_cry_4, S => \N6_data[5]\, Y => OPEN, 
        FCO => next_reg_H6_cry_5);
    
    next_reg_H5_cry_17_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H5_o[17]\, B => 
        hash_control_st_reg_i(6), C => R5_data(17), D => 
        GND_net_1, FCI => next_reg_H5_cry_16, S => \N5_data[17]\, 
        Y => OPEN, FCO => next_reg_H5_cry_17);
    
    \reg_H1[25]\ : SLE
      port map(D => \N1_data[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H1_o[25]\);
    
    next_reg_H3_cry_26_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[26]\, B => 
        hash_control_st_reg_i(6), C => R3_data(26), D => 
        GND_net_1, FCI => next_reg_H3_cry_25, S => \N3_data[26]\, 
        Y => OPEN, FCO => next_reg_H3_cry_26);
    
    next_reg_H3_cry_18_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[18]\, B => 
        hash_control_st_reg_i(6), C => R3_data(18), D => 
        GND_net_1, FCI => next_reg_H3_cry_17, S => \N3_data[18]\, 
        Y => OPEN, FCO => next_reg_H3_cry_18);
    
    next_reg_H0_cry_25_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H0_o[25]\, B => 
        hash_control_st_reg_i(6), C => R0_data(25), D => 
        GND_net_1, FCI => next_reg_H0_cry_24, S => \N0_data[25]\, 
        Y => OPEN, FCO => next_reg_H0_cry_25);
    
    next_reg_H6_cry_1_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[1]\, B => 
        hash_control_st_reg_i(6), C => R6_data(1), D => GND_net_1, 
        FCI => next_reg_H6_cry_0, S => \N6_data[1]\, Y => OPEN, 
        FCO => next_reg_H6_cry_1);
    
    next_reg_H3_cry_4_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H3_o[4]\, B => 
        hash_control_st_reg_i(6), C => R3_data(4), D => GND_net_1, 
        FCI => next_reg_H3_cry_3, S => \N3_data[4]\, Y => OPEN, 
        FCO => next_reg_H3_cry_4);
    
    next_reg_H2_cry_3_0 : ARI1
      generic map(INIT => x"52288")

      port map(A => \SHA256_BLOCK_0_H2_o[3]\, B => 
        hash_control_st_reg_i(6), C => R2_data(3), D => GND_net_1, 
        FCI => next_reg_H2_cry_2, S => \N2_data[3]\, Y => OPEN, 
        FCO => next_reg_H2_cry_3);
    
    \reg_H0[7]\ : SLE
      port map(D => \N0_data[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[7]\);
    
    \reg_H0[11]\ : SLE
      port map(D => \N0_data[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H0_o[11]\);
    
    next_reg_H6_cry_27_0 : ARI1
      generic map(INIT => x"577DD")

      port map(A => \SHA256_BLOCK_0_H6_o[27]\, B => 
        hash_control_st_reg_i(6), C => R6_data(27), D => 
        GND_net_1, FCI => next_reg_H6_cry_26, S => \N6_data[27]\, 
        Y => OPEN, FCO => next_reg_H6_cry_27);
    
    \reg_H2[26]\ : SLE
      port map(D => \N2_data[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_168_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \SHA256_BLOCK_0_H2_o[26]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_padding is

    port( di_o_0                                    : out   std_logic_vector(1 to 1);
          reg_17x32_0_valid_bytes_0                 : in    std_logic_vector(1 downto 0);
          Kt_addr_fast                              : in    std_logic_vector(0 to 0);
          hash_control_st_reg                       : in    std_logic_vector(2 to 2);
          W_out_2_0                                 : out   std_logic_vector(5 to 5);
          W_out_i_i_2                               : out   std_logic_vector(31 to 31);
          W_out_i_i_1                               : out   std_logic_vector(31 to 31);
          W_out_i_1                                 : out   std_logic_vector(1 downto 0);
          W_out_i_0                                 : out   std_logic_vector(2 to 2);
          msg_bitlen                                : in    std_logic_vector(63 downto 3);
          state_2                                   : in    std_logic;
          state_0                                   : in    std_logic;
          state_3                                   : in    std_logic;
          Kt_addr_5                                 : in    std_logic;
          Kt_addr_0                                 : in    std_logic;
          W_out_2_0_0_1                             : out   std_logic;
          W_out_2_0_0_0                             : out   std_logic;
          W_out_2_0_0_3                             : out   std_logic;
          W_out_2_0_1_8                             : out   std_logic;
          W_out_2_0_1_0                             : out   std_logic;
          W_out_2_i_0_18                            : out   std_logic;
          W_out_2_i_0_21                            : out   std_logic;
          W_out_2_i_0_17                            : out   std_logic;
          W_out_2_i_0_22                            : out   std_logic;
          W_out_2_i_0_20                            : out   std_logic;
          W_out_2_i_0_16                            : out   std_logic;
          W_out_2_i_0_19                            : out   std_logic;
          W_out_2_0_2_0                             : out   std_logic;
          W_out_2_0_2_8                             : out   std_logic;
          sha256_controller_0_di_o_3                : in    std_logic;
          sha256_controller_0_di_o_5                : in    std_logic;
          sha256_controller_0_di_o_0                : in    std_logic;
          W_out_2_i_1_18                            : out   std_logic;
          W_out_2_i_1_21                            : out   std_logic;
          W_out_2_i_1_17                            : out   std_logic;
          W_out_2_i_1_22                            : out   std_logic;
          W_out_2_i_1_20                            : out   std_logic;
          W_out_2_i_1_16                            : out   std_logic;
          W_out_2_i_1_19                            : out   std_logic;
          W_out_2_i_1_12                            : out   std_logic;
          W_out_2_i_1_8                             : out   std_logic;
          W_out_2_i_1_10                            : out   std_logic;
          W_out_2_i_1_13                            : out   std_logic;
          W_out_2_i_1_14                            : out   std_logic;
          W_out_2_i_1_11                            : out   std_logic;
          W_out_2_i_1_9                             : out   std_logic;
          W_out_2_i_1_1                             : out   std_logic;
          W_out_2_i_1_2                             : out   std_logic;
          W_out_2_i_1_0                             : out   std_logic;
          W_out_2_i_1_4                             : out   std_logic;
          W_out_2_i_1_3                             : out   std_logic;
          W_out_2_i_1_6                             : out   std_logic;
          W_out_2_i_1_5                             : out   std_logic;
          N_223                                     : in    std_logic;
          N_1702                                    : in    std_logic;
          N_1710                                    : in    std_logic;
          SHA256_Module_0_di_req_o                  : in    std_logic;
          N_388                                     : out   std_logic;
          N_112                                     : in    std_logic;
          one_insert                                : in    std_logic;
          Kt_addr_0_rep2                            : in    std_logic;
          sha_last_blk_reg                          : in    std_logic;
          Kt_addr_4_rep1                            : in    std_logic;
          bytes_sel                                 : in    std_logic;
          ren_pos                                   : in    std_logic;
          N_102                                     : in    std_logic;
          sha_last_blk_next_0_o2_2_out_0            : in    std_logic;
          N_361                                     : in    std_logic;
          SHA256_Module_0_data_available_lastbank_8 : in    std_logic;
          N_111                                     : in    std_logic;
          N_1690                                    : in    std_logic;
          N_245                                     : out   std_logic;
          N_1691                                    : in    std_logic;
          N_248                                     : out   std_logic;
          N_1693                                    : in    std_logic;
          N_251                                     : out   std_logic;
          N_1692                                    : in    std_logic;
          N_349                                     : out   std_logic;
          N_1718                                    : in    std_logic;
          N_1694                                    : in    std_logic;
          N_255                                     : out   std_logic;
          N_1698                                    : in    std_logic;
          N_1701                                    : in    std_logic;
          N_98                                      : out   std_logic;
          N_307                                     : out   std_logic;
          N_1696                                    : in    std_logic;
          N_1697                                    : in    std_logic;
          N_1695                                    : in    std_logic;
          N_1699                                    : in    std_logic;
          N_1707                                    : in    std_logic;
          N_1708                                    : in    std_logic;
          N_1709                                    : in    std_logic;
          N_1706                                    : in    std_logic;
          N_1704                                    : in    std_logic;
          N_1688                                    : in    std_logic;
          N_1687                                    : in    std_logic;
          N_1689                                    : in    std_logic;
          N_1713                                    : in    std_logic;
          N_1716                                    : in    std_logic;
          N_1712                                    : in    std_logic;
          N_1717                                    : in    std_logic;
          N_1715                                    : in    std_logic;
          N_1711                                    : in    std_logic;
          N_1714                                    : in    std_logic;
          N_273                                     : out   std_logic;
          N_266                                     : out   std_logic;
          N_263                                     : out   std_logic;
          N_260                                     : out   std_logic;
          N_287                                     : out   std_logic;
          N_290                                     : out   std_logic;
          N_293                                     : out   std_logic;
          N_296                                     : out   std_logic;
          N_299                                     : out   std_logic;
          N_302                                     : out   std_logic;
          N_305                                     : out   std_logic;
          N_268                                     : out   std_logic;
          N_275                                     : out   std_logic;
          N_278                                     : out   std_logic
        );

end sha256_padding;

architecture DEF_ARCH of sha256_padding is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_116, N_211, \W_out_2_0_2_1[15]_net_1\, N_109, 
        \di_o_0[1]\, N_106, \W_out_2_0_1_1[23]_net_1\, 
        \W_out_2_0_1[23]_net_1\, \N_388\, N_390, 
        \W_out_2_0_a4_1[7]_net_1\, N_392, N_384, 
        \W_out_2_0_o2_0_0[15]_net_1\, \W_out_2_0_o2_0[23]_net_1\, 
        W_out_2_0_o2_out_2, N_108, \W_out_2_i_o2_0_0_tz[8]_net_1\, 
        N_954, \W_out_2_i_o2_4_d[8]_net_1\, N_282, N_333, N_314, 
        N_317, N_320, N_323, N_326, N_329, N_332, N_379, N_393, 
        N_256, \W_out_2_i_o2_4_0_0[8]_net_1\, N_281, N_306, N_334, 
        \W_out_2_i_o2_4_c[8]_net_1\, N_267, N_277, N_405, N_335, 
        \W_out_2_i_0[9]_net_1\, \W_out_2_i_0[10]_net_1\, 
        \W_out_2_i_0[8]_net_1\, \W_out_2_i_0[12]_net_1\, 
        \W_out_2_i_0[20]_net_1\, \W_out_2_i_0[21]_net_1\, 
        \W_out_2_i_0[22]_net_1\, \W_out_2_i_0[19]_net_1\, 
        \W_out_2_i_0[17]_net_1\, N_95, N_286, N_292, N_276, 
        GND_net_1, VCC_net_1 : std_logic;

begin 

    di_o_0(1) <= \di_o_0[1]\;
    N_388 <= \N_388\;

    \W_out_2_i_0[25]\ : CFG4
      generic map(INIT => x"BFAA")

      port map(A => N_317, B => \di_o_0[1]\, C => N_1712, D => 
        N_108, Y => W_out_2_i_0_17);
    
    \W_out_2_i_a2[16]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => N_102, B => one_insert, C => N_116, D => 
        sha_last_blk_next_0_o2_2_out_0, Y => N_379);
    
    \W_out_2_0_o2_s_0[15]\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => hash_control_st_reg(2), B => Kt_addr_4_rep1, 
        C => Kt_addr_5, D => N_384, Y => W_out_2_0_o2_out_2);
    
    \W_out_2_0_o2_0[23]\ : CFG3
      generic map(INIT => x"DF")

      port map(A => bytes_sel, B => reg_17x32_0_valid_bytes_0(1), 
        C => reg_17x32_0_valid_bytes_0(0), Y => 
        \W_out_2_0_o2_0[23]_net_1\);
    
    \W_out_2_0_a2_0[15]\ : CFG2
      generic map(INIT => x"4")

      port map(A => Kt_addr_0_rep2, B => one_insert, Y => \N_388\);
    
    \W_out_2_i_a4_1[28]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => one_insert, B => msg_bitlen(60), C => 
        sha_last_blk_next_0_o2_2_out_0, D => N_102, Y => N_326);
    
    \W_out_2_i_1[28]\ : CFG4
      generic map(INIT => x"5073")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(28), 
        C => N_108, D => N_109, Y => W_out_2_i_1_20);
    
    \W_out_2_i_1[8]\ : CFG4
      generic map(INIT => x"FF01")

      port map(A => msg_bitlen(40), B => 
        \W_out_2_i_o2_4_c[8]_net_1\, C => 
        \W_out_2_i_o2_4_0_0[8]_net_1\, D => 
        \W_out_2_i_0[8]_net_1\, Y => W_out_2_i_1_0);
    
    \W_out_2_0_a2[15]\ : CFG2
      generic map(INIT => x"2")

      port map(A => Kt_addr_fast(0), B => sha_last_blk_reg, Y => 
        N_384);
    
    \W_out_2_i_1[13]\ : CFG4
      generic map(INIT => x"CFEF")

      port map(A => N_108, B => N_276, C => N_405, D => 
        sha256_controller_0_di_o_0, Y => W_out_2_i_1_5);
    
    \W_out_2_i_0[17]\ : CFG4
      generic map(INIT => x"B0F0")

      port map(A => N_116, B => \di_o_0[1]\, C => N_108, D => 
        N_1704, Y => \W_out_2_i_0[17]_net_1\);
    
    \W_out_2_0_a4_0[15]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \N_388\, B => N_116, C => \di_o_0[1]\, D => 
        N_1702, Y => N_281);
    
    \W_out_2_0_0[6]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(38), B => msg_bitlen(6), C => 
        N_111, D => N_109, Y => W_out_2_0_0_3);
    
    \W_out_2_i_a4_1[16]\ : CFG4
      generic map(INIT => x"4505")

      port map(A => msg_bitlen(48), B => N_116, C => N_111, D => 
        N_109, Y => N_287);
    
    \W_out_2_i_0[10]\ : CFG4
      generic map(INIT => x"7F33")

      port map(A => N_1697, B => N_405, C => \di_o_0[1]\, D => 
        N_108, Y => \W_out_2_i_0[10]_net_1\);
    
    \W_out_2_0_a2[7]\ : CFG2
      generic map(INIT => x"8")

      port map(A => SHA256_Module_0_di_req_o, B => one_insert, Y
         => N_390);
    
    \W_out_2_i_o2_0[8]\ : CFG3
      generic map(INIT => x"B3")

      port map(A => \W_out_2_i_o2_0_0_tz[8]_net_1\, B => N_109, C
         => N_211, Y => N_95);
    
    \W_out_2_i_1[22]\ : CFG4
      generic map(INIT => x"FF51")

      port map(A => msg_bitlen(22), B => N_109, C => N_379, D => 
        \W_out_2_i_0[22]_net_1\, Y => W_out_2_i_1_14);
    
    \W_out_2_i_0[24]\ : CFG4
      generic map(INIT => x"BFAA")

      port map(A => N_314, B => \di_o_0[1]\, C => N_1711, D => 
        N_108, Y => W_out_2_i_0_16);
    
    \W_out_2_i_a4_1[18]\ : CFG4
      generic map(INIT => x"4505")

      port map(A => msg_bitlen(50), B => N_116, C => N_111, D => 
        N_109, Y => N_293);
    
    \W_out_2_i_0[28]\ : CFG4
      generic map(INIT => x"BFAA")

      port map(A => N_326, B => \di_o_0[1]\, C => N_1715, D => 
        N_108, Y => W_out_2_i_0_20);
    
    \W_out_2_i_0[19]\ : CFG4
      generic map(INIT => x"B0F0")

      port map(A => N_116, B => \di_o_0[1]\, C => N_108, D => 
        N_1706, Y => \W_out_2_i_0[19]_net_1\);
    
    \W_out_i_0[2]\ : CFG4
      generic map(INIT => x"35F5")

      port map(A => msg_bitlen(34), B => \di_o_0[1]\, C => N_111, 
        D => N_1689, Y => W_out_i_0(2));
    
    \W_out_2_0_o2[7]\ : CFG4
      generic map(INIT => x"FFF7")

      port map(A => sha_last_blk_reg, B => Kt_addr_0, C => 
        \W_out_2_0_o2_0_0[15]_net_1\, D => N_102, Y => N_109);
    
    \W_out_2_0_a4[6]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \di_o_0[1]\, B => N_1693, C => N_393, Y => 
        N_251);
    
    \W_out_2_0_1_1[23]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => \di_o_0[1]\, B => SHA256_Module_0_di_req_o, C
         => \N_388\, Y => \W_out_2_0_1_1[23]_net_1\);
    
    \W_out_2_0_o2[15]\ : CFG2
      generic map(INIT => x"E")

      port map(A => W_out_2_0_o2_out_2, B => N_102, Y => N_106);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \W_out_2_i_1[14]\ : CFG4
      generic map(INIT => x"DFDD")

      port map(A => N_405, B => N_277, C => msg_bitlen(14), D => 
        N_95, Y => W_out_2_i_1_6);
    
    \W_out_2_i_0[22]\ : CFG4
      generic map(INIT => x"B0F0")

      port map(A => N_116, B => \di_o_0[1]\, C => N_108, D => 
        N_1709, Y => \W_out_2_i_0[22]_net_1\);
    
    \W_out_2_0_1[15]\ : CFG4
      generic map(INIT => x"EEFE")

      port map(A => N_282, B => N_281, C => msg_bitlen(47), D => 
        N_111, Y => W_out_2_0_1_8);
    
    \W_out_2_0_a4_1[7]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => one_insert, B => msg_bitlen(39), C => 
        sha_last_blk_next_0_o2_2_out_0, D => N_102, Y => N_256);
    
    \W_out_2_0_a4_0[23]\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_390, B => N_116, C => N_109, Y => N_307);
    
    \W_out_2_i_1[18]\ : CFG4
      generic map(INIT => x"FF8A")

      port map(A => N_108, B => N_116, C => 
        sha256_controller_0_di_o_5, D => N_292, Y => 
        W_out_2_i_1_10);
    
    \W_out_2_0_a4_1[15]\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_392, B => N_109, C => N_390, Y => N_282);
    
    \W_out_2_i_o2_0_3[8]\ : CFG4
      generic map(INIT => x"0D05")

      port map(A => N_109, B => N_211, C => msg_bitlen(10), D => 
        \W_out_2_i_o2_0_0_tz[8]_net_1\, Y => N_266);
    
    \W_out_2_i_0[8]\ : CFG4
      generic map(INIT => x"7F33")

      port map(A => N_1695, B => N_405, C => \di_o_0[1]\, D => 
        N_108, Y => \W_out_2_i_0[8]_net_1\);
    
    \W_out_i_1[1]\ : CFG4
      generic map(INIT => x"35F5")

      port map(A => msg_bitlen(33), B => \di_o_0[1]\, C => N_111, 
        D => N_1688, Y => W_out_i_1(1));
    
    \W_out_2_i_a4_1[20]\ : CFG4
      generic map(INIT => x"4505")

      port map(A => msg_bitlen(52), B => N_116, C => N_111, D => 
        N_109, Y => N_299);
    
    \W_out_2_a4[5]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \di_o_0[1]\, B => N_1692, C => N_393, Y => 
        N_349);
    
    \W_out_2_i_o2_4_0_0[8]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \W_out_2_i_o2_4_d[8]_net_1\, B => N_954, C
         => N_390, Y => \W_out_2_i_o2_4_0_0[8]_net_1\);
    
    \W_out_2_i_1[12]\ : CFG4
      generic map(INIT => x"FF01")

      port map(A => msg_bitlen(44), B => 
        \W_out_2_i_o2_4_c[8]_net_1\, C => 
        \W_out_2_i_o2_4_0_0[8]_net_1\, D => 
        \W_out_2_i_0[12]_net_1\, Y => W_out_2_i_1_4);
    
    \W_out_2_0_o2_0_0[15]\ : CFG3
      generic map(INIT => x"FB")

      port map(A => Kt_addr_5, B => hash_control_st_reg(2), C => 
        Kt_addr_4_rep1, Y => \W_out_2_0_o2_0_0[15]_net_1\);
    
    \W_out_2_0_a4[23]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => N_116, B => \di_o_0[1]\, C => N_106, D => 
        N_1710, Y => N_306);
    
    \W_out_2_0_1[23]\ : CFG4
      generic map(INIT => x"50DC")

      port map(A => \W_out_2_0_1_1[23]_net_1\, B => 
        msg_bitlen(23), C => N_1710, D => N_109, Y => 
        \W_out_2_0_1[23]_net_1\);
    
    \W_out_2_i_1[26]\ : CFG4
      generic map(INIT => x"5073")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(26), 
        C => N_108, D => N_109, Y => W_out_2_i_1_18);
    
    \W_out_2_0_o2_2[15]\ : CFG3
      generic map(INIT => x"8F")

      port map(A => reg_17x32_0_valid_bytes_0(1), B => 
        reg_17x32_0_valid_bytes_0(0), C => N_361, Y => N_954);
    
    \W_out_2_0_o2_1[15]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => SHA256_Module_0_di_req_o, B => 
        \W_out_2_0_o2_0[23]_net_1\, C => 
        SHA256_Module_0_data_available_lastbank_8, D => state_0, 
        Y => N_116);
    
    \W_out_2_0_2[15]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \W_out_2_0_2_1[15]_net_1\, B => N_1702, C => 
        msg_bitlen(15), D => N_109, Y => W_out_2_0_2_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \W_out_2_0_0[4]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(36), B => msg_bitlen(4), C => 
        N_111, D => N_109, Y => W_out_2_0_0_1);
    
    \W_out_2_i_a4_1[27]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => one_insert, B => msg_bitlen(59), C => 
        sha_last_blk_next_0_o2_2_out_0, D => N_102, Y => N_323);
    
    \W_out_2_0_a4[4]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \di_o_0[1]\, B => N_1691, C => N_393, Y => 
        N_248);
    
    \W_out_2_0_0[3]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(35), B => msg_bitlen(3), C => 
        N_111, D => N_109, Y => W_out_2_0_0_0);
    
    \W_out_2_i_1[21]\ : CFG4
      generic map(INIT => x"FF51")

      port map(A => msg_bitlen(21), B => N_109, C => N_379, D => 
        \W_out_2_i_0[21]_net_1\, Y => W_out_2_i_1_13);
    
    \W_out_2_i_o2_0_2[8]\ : CFG4
      generic map(INIT => x"0D05")

      port map(A => N_109, B => N_211, C => msg_bitlen(9), D => 
        \W_out_2_i_o2_0_0_tz[8]_net_1\, Y => N_263);
    
    \W_out_2_i_a4[14]\ : CFG3
      generic map(INIT => x"70")

      port map(A => N_1701, B => \di_o_0[1]\, C => N_108, Y => 
        N_277);
    
    \W_out_2_i_1[27]\ : CFG4
      generic map(INIT => x"5073")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(27), 
        C => N_108, D => N_109, Y => W_out_2_i_1_19);
    
    \W_out_2_i_1[20]\ : CFG4
      generic map(INIT => x"FF51")

      port map(A => msg_bitlen(20), B => N_109, C => N_379, D => 
        \W_out_2_i_0[20]_net_1\, Y => W_out_2_i_1_12);
    
    \W_out_2_i_o2[8]\ : CFG4
      generic map(INIT => x"0F1F")

      port map(A => N_102, B => \N_388\, C => N_211, D => 
        W_out_2_0_o2_out_2, Y => N_405);
    
    \W_out_2_i_0[26]\ : CFG4
      generic map(INIT => x"BFAA")

      port map(A => N_320, B => \di_o_0[1]\, C => N_1713, D => 
        N_108, Y => W_out_2_i_0_18);
    
    \W_out_2_i_a4_1[17]\ : CFG4
      generic map(INIT => x"4505")

      port map(A => msg_bitlen(49), B => N_116, C => N_111, D => 
        N_109, Y => N_290);
    
    \W_out_i_i_a4_1[31]\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_1718, B => \N_388\, C => \di_o_0[1]\, Y => 
        N_335);
    
    \W_out_2_0_2[23]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => N_111, B => msg_bitlen(55), C => N_306, D => 
        \W_out_2_0_1[23]_net_1\, Y => W_out_2_0_2_8);
    
    \W_out_i_i_a4_0[31]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \di_o_0[1]\, B => SHA256_Module_0_di_req_o, C
         => N_1718, D => N_106, Y => N_334);
    
    \W_out_2_i_1[9]\ : CFG4
      generic map(INIT => x"FF01")

      port map(A => msg_bitlen(41), B => 
        \W_out_2_i_o2_4_c[8]_net_1\, C => 
        \W_out_2_i_o2_4_0_0[8]_net_1\, D => 
        \W_out_2_i_0[9]_net_1\, Y => W_out_2_i_1_1);
    
    \W_out_i_i_2[31]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => N_334, B => msg_bitlen(31), C => N_109, Y => 
        W_out_i_i_2(31));
    
    \W_out_2_i_1[29]\ : CFG4
      generic map(INIT => x"5073")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(29), 
        C => N_108, D => N_109, Y => W_out_2_i_1_21);
    
    \W_out_2_i_0[21]\ : CFG4
      generic map(INIT => x"B0F0")

      port map(A => N_116, B => \di_o_0[1]\, C => N_108, D => 
        N_1708, Y => \W_out_2_i_0[21]_net_1\);
    
    \W_out_2_0_a2_1[15]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_223, B => reg_17x32_0_valid_bytes_0(0), Y
         => N_392);
    
    \W_out_2_i_a4_0[13]\ : CFG3
      generic map(INIT => x"01")

      port map(A => msg_bitlen(45), B => 
        \W_out_2_i_o2_4_c[8]_net_1\, C => 
        \W_out_2_i_o2_4_0_0[8]_net_1\, Y => N_275);
    
    \W_out_2_i_0[12]\ : CFG4
      generic map(INIT => x"7F33")

      port map(A => N_1699, B => N_405, C => \di_o_0[1]\, D => 
        N_108, Y => \W_out_2_i_0[12]_net_1\);
    
    \W_out_2_0_a4_0[7]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \di_o_0[1]\, B => N_1694, C => N_393, Y => 
        N_255);
    
    \W_out_2_i_0[27]\ : CFG4
      generic map(INIT => x"BFAA")

      port map(A => N_323, B => \di_o_0[1]\, C => N_1714, D => 
        N_108, Y => W_out_2_i_0_19);
    
    \W_out_2_i_o2_0_0_tz[8]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => one_insert, B => N_102, C => 
        sha_last_blk_next_0_o2_2_out_0, Y => 
        \W_out_2_i_o2_0_0_tz[8]_net_1\);
    
    \W_out_2_i_0[20]\ : CFG4
      generic map(INIT => x"B0F0")

      port map(A => N_116, B => \di_o_0[1]\, C => N_108, D => 
        N_1707, Y => \W_out_2_i_0[20]_net_1\);
    
    \W_out_2_i_1[16]\ : CFG4
      generic map(INIT => x"FF8A")

      port map(A => N_108, B => N_116, C => 
        sha256_controller_0_di_o_3, D => N_286, Y => 
        W_out_2_i_1_8);
    
    \W_out_i_1[0]\ : CFG4
      generic map(INIT => x"35F5")

      port map(A => msg_bitlen(32), B => \di_o_0[1]\, C => N_111, 
        D => N_1687, Y => W_out_i_1(0));
    
    \W_out_2_i_a4_0[14]\ : CFG3
      generic map(INIT => x"01")

      port map(A => msg_bitlen(46), B => 
        \W_out_2_i_o2_4_c[8]_net_1\, C => 
        \W_out_2_i_o2_4_0_0[8]_net_1\, Y => N_278);
    
    \W_out_2_i_0[9]\ : CFG4
      generic map(INIT => x"7F33")

      port map(A => N_1696, B => N_405, C => \di_o_0[1]\, D => 
        N_108, Y => \W_out_2_i_0[9]_net_1\);
    
    \W_out_2_0[5]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => msg_bitlen(37), B => msg_bitlen(5), C => 
        N_111, D => N_109, Y => W_out_2_0(5));
    
    \W_out_2_i_a4_1[30]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => one_insert, B => msg_bitlen(62), C => 
        sha_last_blk_next_0_o2_2_out_0, D => N_102, Y => N_332);
    
    \W_out_2_i_1[11]\ : CFG4
      generic map(INIT => x"DFDD")

      port map(A => N_405, B => N_267, C => msg_bitlen(11), D => 
        N_95, Y => W_out_2_i_1_3);
    
    \W_out_2_0_a4[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \di_o_0[1]\, B => N_1690, C => N_393, Y => 
        N_245);
    
    \W_out_2_i_a4_1[22]\ : CFG4
      generic map(INIT => x"4505")

      port map(A => msg_bitlen(54), B => N_116, C => N_111, D => 
        N_109, Y => N_305);
    
    \W_out_2_i_a4[11]\ : CFG3
      generic map(INIT => x"70")

      port map(A => N_1698, B => \di_o_0[1]\, C => N_108, Y => 
        N_267);
    
    \W_out_2_i_0[29]\ : CFG4
      generic map(INIT => x"BFAA")

      port map(A => N_329, B => \di_o_0[1]\, C => N_1716, D => 
        N_108, Y => W_out_2_i_0_21);
    
    \W_out_2_i_a4_1[29]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => one_insert, B => msg_bitlen(61), C => 
        sha_last_blk_next_0_o2_2_out_0, D => N_102, Y => N_329);
    
    \W_out_2_i_1[17]\ : CFG4
      generic map(INIT => x"FF51")

      port map(A => msg_bitlen(17), B => N_109, C => N_379, D => 
        \W_out_2_i_0[17]_net_1\, Y => W_out_2_i_1_9);
    
    \W_out_2_i_a4_2[24]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => one_insert, B => msg_bitlen(56), C => 
        sha_last_blk_next_0_o2_2_out_0, D => N_102, Y => N_314);
    
    \W_out_2_i_1[10]\ : CFG4
      generic map(INIT => x"FF01")

      port map(A => msg_bitlen(42), B => 
        \W_out_2_i_o2_4_c[8]_net_1\, C => 
        \W_out_2_i_o2_4_0_0[8]_net_1\, D => 
        \W_out_2_i_0[10]_net_1\, Y => W_out_2_i_1_2);
    
    \W_out_2_i_a4_0[11]\ : CFG3
      generic map(INIT => x"01")

      port map(A => msg_bitlen(43), B => 
        \W_out_2_i_o2_4_c[8]_net_1\, C => 
        \W_out_2_i_o2_4_0_0[8]_net_1\, Y => N_268);
    
    \W_out_2_0_a4_0_0[3]\ : CFG4
      generic map(INIT => x"AAA8")

      port map(A => ren_pos, B => state_2, C => state_0, D => 
        state_3, Y => \di_o_0[1]\);
    
    \W_out_2_i_o2_5[8]\ : CFG3
      generic map(INIT => x"CD")

      port map(A => N_223, B => N_116, C => 
        reg_17x32_0_valid_bytes_0(0), Y => N_211);
    
    \W_out_2_0_1[7]\ : CFG4
      generic map(INIT => x"FEBA")

      port map(A => N_256, B => N_109, C => msg_bitlen(7), D => 
        \W_out_2_0_a4_1[7]_net_1\, Y => W_out_2_0_1_0);
    
    \W_out_2_i_o2_0_1[8]\ : CFG4
      generic map(INIT => x"0D05")

      port map(A => N_109, B => N_211, C => msg_bitlen(8), D => 
        \W_out_2_i_o2_0_0_tz[8]_net_1\, Y => N_260);
    
    \W_out_2_0_2_1[15]\ : CFG3
      generic map(INIT => x"40")

      port map(A => N_211, B => \di_o_0[1]\, C => N_106, Y => 
        \W_out_2_0_2_1[15]_net_1\);
    
    \W_out_2_i_a4_0[16]\ : CFG4
      generic map(INIT => x"4055")

      port map(A => msg_bitlen(16), B => N_116, C => N_111, D => 
        N_109, Y => N_286);
    
    \W_out_2_i_1[25]\ : CFG4
      generic map(INIT => x"5073")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(25), 
        C => N_108, D => N_109, Y => W_out_2_i_1_17);
    
    \W_out_2_i_a4_1[13]\ : CFG4
      generic map(INIT => x"0D05")

      port map(A => N_109, B => N_211, C => msg_bitlen(13), D => 
        \W_out_2_i_o2_0_0_tz[8]_net_1\, Y => N_276);
    
    \W_out_i_i_a4[31]\ : CFG3
      generic map(INIT => x"40")

      port map(A => SHA256_Module_0_di_req_o, B => N_109, C => 
        one_insert, Y => N_333);
    
    \W_out_2_0_a4_1_0[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_390, B => reg_17x32_0_valid_bytes_0(1), C
         => N_112, Y => \W_out_2_0_a4_1[7]_net_1\);
    
    \W_out_2_i_o2_4_c[8]\ : CFG4
      generic map(INIT => x"000E")

      port map(A => sha_last_blk_next_0_o2_2_out_0, B => N_102, C
         => N_392, D => N_116, Y => \W_out_2_i_o2_4_c[8]_net_1\);
    
    \W_out_2_i_a4_1[25]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => one_insert, B => msg_bitlen(57), C => 
        sha_last_blk_next_0_o2_2_out_0, D => N_102, Y => N_317);
    
    \W_out_2_i_a4_1[19]\ : CFG4
      generic map(INIT => x"4505")

      port map(A => msg_bitlen(51), B => N_116, C => N_111, D => 
        N_109, Y => N_296);
    
    \W_out_2_i_1[19]\ : CFG4
      generic map(INIT => x"FF51")

      port map(A => msg_bitlen(19), B => N_109, C => N_379, D => 
        \W_out_2_i_0[19]_net_1\, Y => W_out_2_i_1_11);
    
    \W_out_2_0_a2[3]\ : CFG3
      generic map(INIT => x"20")

      port map(A => SHA256_Module_0_di_req_o, B => N_361, C => 
        N_108, Y => N_393);
    
    \W_out_2_i_o2[24]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \N_388\, B => N_102, C => W_out_2_0_o2_out_2, 
        Y => N_108);
    
    \W_out_2_i_a4_0[18]\ : CFG4
      generic map(INIT => x"4055")

      port map(A => msg_bitlen(18), B => N_116, C => N_111, D => 
        N_109, Y => N_292);
    
    \W_out_2_i_0[30]\ : CFG4
      generic map(INIT => x"BFAA")

      port map(A => N_332, B => \di_o_0[1]\, C => N_1717, D => 
        N_108, Y => W_out_2_i_0_22);
    
    \W_out_2_i_a4_1[21]\ : CFG4
      generic map(INIT => x"4505")

      port map(A => msg_bitlen(53), B => N_116, C => N_111, D => 
        N_109, Y => N_302);
    
    \W_out_i_o2[0]\ : CFG4
      generic map(INIT => x"2F0F")

      port map(A => SHA256_Module_0_di_req_o, B => N_361, C => 
        N_111, D => N_109, Y => N_98);
    
    \W_out_i_i_1[31]\ : CFG4
      generic map(INIT => x"EEFE")

      port map(A => N_333, B => N_335, C => msg_bitlen(63), D => 
        N_111, Y => W_out_i_i_1(31));
    
    \W_out_2_i_o2_4_d[8]\ : CFG4
      generic map(INIT => x"0040")

      port map(A => N_102, B => sha_last_blk_next_0_o2_2_out_0, C
         => sha_last_blk_reg, D => \W_out_2_0_o2_0_0[15]_net_1\, 
        Y => \W_out_2_i_o2_4_d[8]_net_1\);
    
    \W_out_2_i_o2_0_4[8]\ : CFG4
      generic map(INIT => x"0D05")

      port map(A => N_109, B => N_211, C => msg_bitlen(12), D => 
        \W_out_2_i_o2_0_0_tz[8]_net_1\, Y => N_273);
    
    \W_out_2_i_a4_1[26]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => one_insert, B => msg_bitlen(58), C => 
        sha_last_blk_next_0_o2_2_out_0, D => N_102, Y => N_320);
    
    \W_out_2_i_1[30]\ : CFG4
      generic map(INIT => x"5073")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(30), 
        C => N_108, D => N_109, Y => W_out_2_i_1_22);
    
    \W_out_2_i_1[24]\ : CFG4
      generic map(INIT => x"5073")

      port map(A => SHA256_Module_0_di_req_o, B => msg_bitlen(24), 
        C => N_108, D => N_109, Y => W_out_2_i_1_16);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_msg_sch is

    port( Wt_data                              : out   std_logic_vector(31 downto 0);
          W_out_2_0                            : in    std_logic_vector(5 to 5);
          W_out_i_i_2                          : in    std_logic_vector(31 to 31);
          W_out_i_i_1                          : in    std_logic_vector(31 to 31);
          W_out_2_i_0                          : in    std_logic_vector(30 downto 24);
          W_out_i_0                            : in    std_logic_vector(2 to 2);
          W_out_i_1                            : in    std_logic_vector(1 downto 0);
          W_out_2_0_0_3                        : in    std_logic;
          W_out_2_0_0_1                        : in    std_logic;
          W_out_2_0_0_0                        : in    std_logic;
          W_out_2_0_2_8                        : in    std_logic;
          W_out_2_0_2_0                        : in    std_logic;
          W_out_2_0_1_0                        : in    std_logic;
          W_out_2_0_1_8                        : in    std_logic;
          W_out_2_i_1_22                       : in    std_logic;
          W_out_2_i_1_21                       : in    std_logic;
          W_out_2_i_1_20                       : in    std_logic;
          W_out_2_i_1_19                       : in    std_logic;
          W_out_2_i_1_18                       : in    std_logic;
          W_out_2_i_1_17                       : in    std_logic;
          W_out_2_i_1_16                       : in    std_logic;
          W_out_2_i_1_14                       : in    std_logic;
          W_out_2_i_1_13                       : in    std_logic;
          W_out_2_i_1_12                       : in    std_logic;
          W_out_2_i_1_11                       : in    std_logic;
          W_out_2_i_1_10                       : in    std_logic;
          W_out_2_i_1_9                        : in    std_logic;
          W_out_2_i_1_8                        : in    std_logic;
          W_out_2_i_1_6                        : in    std_logic;
          W_out_2_i_1_5                        : in    std_logic;
          W_out_2_i_1_4                        : in    std_logic;
          W_out_2_i_1_3                        : in    std_logic;
          W_out_2_i_1_2                        : in    std_logic;
          W_out_2_i_1_1                        : in    std_logic;
          W_out_2_i_1_0                        : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          N_244_i_0                            : in    std_logic;
          next_r0_0_cry_0_Y                    : out   std_logic;
          N_251                                : in    std_logic;
          ld_i_i_3                             : in    std_logic;
          N_349                                : in    std_logic;
          N_248                                : in    std_logic;
          N_245                                : in    std_logic;
          N_255                                : in    std_logic;
          N_98                                 : in    std_logic;
          N_307                                : in    std_logic;
          N_305                                : in    std_logic;
          N_302                                : in    std_logic;
          N_299                                : in    std_logic;
          N_296                                : in    std_logic;
          N_293                                : in    std_logic;
          N_290                                : in    std_logic;
          N_287                                : in    std_logic;
          N_278                                : in    std_logic;
          N_275                                : in    std_logic;
          N_273                                : in    std_logic;
          N_268                                : in    std_logic;
          N_266                                : in    std_logic;
          N_263                                : in    std_logic;
          N_260                                : in    std_logic
        );

end sha256_msg_sch;

architecture DEF_ARCH of sha256_msg_sch is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \r13[18]_net_1\, VCC_net_1, \r14[18]_net_1\, 
        GND_net_1, \r13[19]_net_1\, \r14[19]_net_1\, 
        \r13[20]_net_1\, \r14[20]_net_1\, \r13[21]_net_1\, 
        \r14[21]_net_1\, \r13[22]_net_1\, \r14[22]_net_1\, 
        \r13[23]_net_1\, \r14[23]_net_1\, \r13[24]_net_1\, 
        \r14[24]_net_1\, \r13[25]_net_1\, \r14[25]_net_1\, 
        \r13[26]_net_1\, \r14[26]_net_1\, \r13[27]_net_1\, 
        \r14[27]_net_1\, \r13[28]_net_1\, \r14[28]_net_1\, 
        \r13[29]_net_1\, \r14[29]_net_1\, \r13[30]_net_1\, 
        \r14[30]_net_1\, \r13[31]_net_1\, \r14[31]_net_1\, 
        \r13[3]_net_1\, \r14[3]_net_1\, \r13[4]_net_1\, 
        \r14[4]_net_1\, \r13[5]_net_1\, \r14[5]_net_1\, 
        \r13[6]_net_1\, \r14[6]_net_1\, \r13[7]_net_1\, 
        \r14[7]_net_1\, \r13[8]_net_1\, \r14[8]_net_1\, 
        \r13[9]_net_1\, \r14[9]_net_1\, \r13[10]_net_1\, 
        \r14[10]_net_1\, \r13[11]_net_1\, \r14[11]_net_1\, 
        \r13[12]_net_1\, \r14[12]_net_1\, \r13[13]_net_1\, 
        \r14[13]_net_1\, \r13[14]_net_1\, \r14[14]_net_1\, 
        \r13[15]_net_1\, \r14[15]_net_1\, \r13[16]_net_1\, 
        \r14[16]_net_1\, \r13[17]_net_1\, \r14[17]_net_1\, 
        \r15[20]_net_1\, \r15[21]_net_1\, \r15[22]_net_1\, 
        \r15[23]_net_1\, \r15[24]_net_1\, \r15[25]_net_1\, 
        \r15[26]_net_1\, \r15[27]_net_1\, \r15[28]_net_1\, 
        \r15[29]_net_1\, \r15[30]_net_1\, \r15[31]_net_1\, 
        \r13[0]_net_1\, \r14[0]_net_1\, \r13[1]_net_1\, 
        \r14[1]_net_1\, \r13[2]_net_1\, \r14[2]_net_1\, 
        \r15[5]_net_1\, \r15[6]_net_1\, \r15[7]_net_1\, 
        \r15[8]_net_1\, \r15[9]_net_1\, \r15[10]_net_1\, 
        \r15[11]_net_1\, \r15[12]_net_1\, \r15[13]_net_1\, 
        \r15[14]_net_1\, \r15[15]_net_1\, \r15[16]_net_1\, 
        \r15[17]_net_1\, \r15[18]_net_1\, \r15[19]_net_1\, 
        \r6[22]_net_1\, \r7[22]_net_1\, \r6[23]_net_1\, 
        \r7[23]_net_1\, \r6[24]_net_1\, \r7[24]_net_1\, 
        \r6[25]_net_1\, \r7[25]_net_1\, \r6[26]_net_1\, 
        \r7[26]_net_1\, \r6[27]_net_1\, \r7[27]_net_1\, 
        \r6[28]_net_1\, \r7[28]_net_1\, \r6[29]_net_1\, 
        \r7[29]_net_1\, \r6[30]_net_1\, \r7[30]_net_1\, 
        \r6[31]_net_1\, \r7[31]_net_1\, \r15[0]_net_1\, 
        \r15[1]_net_1\, \r15[2]_net_1\, \r15[3]_net_1\, 
        \r15[4]_net_1\, \r6[7]_net_1\, \r7[7]_net_1\, 
        \r6[8]_net_1\, \r7[8]_net_1\, \r6[9]_net_1\, 
        \r7[9]_net_1\, \r6[10]_net_1\, \r7[10]_net_1\, 
        \r6[11]_net_1\, \r7[11]_net_1\, \r6[12]_net_1\, 
        \r7[12]_net_1\, \r6[13]_net_1\, \r7[13]_net_1\, 
        \r6[14]_net_1\, \r7[14]_net_1\, \r6[15]_net_1\, 
        \r7[15]_net_1\, \r6[16]_net_1\, \r7[16]_net_1\, 
        \r6[17]_net_1\, \r7[17]_net_1\, \r6[18]_net_1\, 
        \r7[18]_net_1\, \r6[19]_net_1\, \r7[19]_net_1\, 
        \r6[20]_net_1\, \r7[20]_net_1\, \r6[21]_net_1\, 
        \r7[21]_net_1\, \r5[24]_net_1\, \r5[25]_net_1\, 
        \r5[26]_net_1\, \r5[27]_net_1\, \r5[28]_net_1\, 
        \r5[29]_net_1\, \r5[30]_net_1\, \r5[31]_net_1\, 
        \r6[0]_net_1\, \r7[0]_net_1\, \r6[1]_net_1\, 
        \r7[1]_net_1\, \r6[2]_net_1\, \r7[2]_net_1\, 
        \r6[3]_net_1\, \r7[3]_net_1\, \r6[4]_net_1\, 
        \r7[4]_net_1\, \r6[5]_net_1\, \r7[5]_net_1\, 
        \r6[6]_net_1\, \r7[6]_net_1\, \r5[9]_net_1\, 
        \r5[10]_net_1\, \r5[11]_net_1\, \r5[12]_net_1\, 
        \r5[13]_net_1\, \r5[14]_net_1\, \r5[15]_net_1\, 
        \r5[16]_net_1\, \r5[17]_net_1\, \r5[18]_net_1\, 
        \r5[19]_net_1\, \r5[20]_net_1\, \r5[21]_net_1\, 
        \r5[22]_net_1\, \r5[23]_net_1\, \r4[26]_net_1\, 
        \r4[27]_net_1\, \r4[28]_net_1\, \r4[29]_net_1\, 
        \r4[30]_net_1\, \r4[31]_net_1\, \r5[0]_net_1\, 
        \r5[1]_net_1\, \r5[2]_net_1\, \r5[3]_net_1\, 
        \r5[4]_net_1\, \r5[5]_net_1\, \r5[6]_net_1\, 
        \r5[7]_net_1\, \r5[8]_net_1\, \r4[11]_net_1\, 
        \r4[12]_net_1\, \r4[13]_net_1\, \r4[14]_net_1\, 
        \r4[15]_net_1\, \r4[16]_net_1\, \r4[17]_net_1\, 
        \r4[18]_net_1\, \r4[19]_net_1\, \r4[20]_net_1\, 
        \r4[21]_net_1\, \r4[22]_net_1\, \r4[23]_net_1\, 
        \r4[24]_net_1\, \r4[25]_net_1\, \r3[28]_net_1\, 
        \r3[29]_net_1\, \r3[30]_net_1\, \r3[31]_net_1\, 
        \r4[0]_net_1\, \r4[1]_net_1\, \r4[2]_net_1\, 
        \r4[3]_net_1\, \r4[4]_net_1\, \r4[5]_net_1\, 
        \r4[6]_net_1\, \r4[7]_net_1\, \r4[8]_net_1\, 
        \r4[9]_net_1\, \r4[10]_net_1\, \r3[13]_net_1\, 
        \r3[14]_net_1\, \r3[15]_net_1\, \r3[16]_net_1\, 
        \r3[17]_net_1\, \r3[18]_net_1\, \r3[19]_net_1\, 
        \r3[20]_net_1\, \r3[21]_net_1\, \r3[22]_net_1\, 
        \r3[23]_net_1\, \r3[24]_net_1\, \r3[25]_net_1\, 
        \r3[26]_net_1\, \r3[27]_net_1\, \r2[30]_net_1\, 
        \r2[31]_net_1\, \r3[0]_net_1\, \r3[1]_net_1\, 
        \r3[2]_net_1\, \r3[3]_net_1\, \r3[4]_net_1\, 
        \r3[5]_net_1\, \r3[6]_net_1\, \r3[7]_net_1\, 
        \r3[8]_net_1\, \r3[9]_net_1\, \r3[10]_net_1\, 
        \r3[11]_net_1\, \r3[12]_net_1\, \r2[15]_net_1\, 
        \r2[16]_net_1\, \r2[17]_net_1\, \r2[18]_net_1\, 
        \r2[19]_net_1\, \r2[20]_net_1\, \r2[21]_net_1\, 
        \r2[22]_net_1\, \r2[23]_net_1\, \r2[24]_net_1\, 
        \r2[25]_net_1\, \r2[26]_net_1\, \r2[27]_net_1\, 
        \r2[28]_net_1\, \r2[29]_net_1\, \r2[0]_net_1\, 
        \r2[1]_net_1\, \r2[2]_net_1\, \r2[3]_net_1\, 
        \r2[4]_net_1\, \r2[5]_net_1\, \r2[6]_net_1\, 
        \r2[7]_net_1\, \r2[8]_net_1\, \r2[9]_net_1\, 
        \r2[10]_net_1\, \r2[11]_net_1\, \r2[12]_net_1\, 
        \r2[13]_net_1\, \r2[14]_net_1\, \r1[17]_net_1\, 
        \r1[18]_net_1\, \r1[19]_net_1\, \r1[20]_net_1\, 
        \r1[21]_net_1\, \r1[22]_net_1\, \r1[23]_net_1\, 
        \r1[24]_net_1\, \r1[25]_net_1\, \r1[26]_net_1\, 
        \r1[27]_net_1\, \r1[28]_net_1\, \r1[29]_net_1\, 
        \r1[30]_net_1\, \r1[31]_net_1\, \r1[2]_net_1\, 
        \r1[3]_net_1\, \r1[4]_net_1\, \r1[5]_net_1\, 
        \r1[6]_net_1\, \r1[7]_net_1\, \r1[8]_net_1\, 
        \r1[9]_net_1\, \r1[10]_net_1\, \r1[11]_net_1\, 
        \r1[12]_net_1\, \r1[13]_net_1\, \r1[14]_net_1\, 
        \r1[15]_net_1\, \r1[16]_net_1\, \r0[19]_net_1\, 
        \Wt_data[19]\, \r0[20]_net_1\, \Wt_data[20]\, 
        \r0[21]_net_1\, \Wt_data[21]\, \r0[22]_net_1\, 
        \Wt_data[22]\, \r0[23]_net_1\, \Wt_data[23]\, 
        \r0[24]_net_1\, \Wt_data[24]\, \r0[25]_net_1\, 
        \Wt_data[25]\, \r0[26]_net_1\, \Wt_data[26]\, 
        \r0[27]_net_1\, \Wt_data[27]\, \r0[28]_net_1\, 
        \Wt_data[28]\, \r0[29]_net_1\, \Wt_data[29]\, 
        \r0[30]_net_1\, \Wt_data[30]\, \r0[31]_net_1\, 
        \Wt_data[31]\, \r1[0]_net_1\, \r1[1]_net_1\, 
        \r0[4]_net_1\, \Wt_data[4]\, \r0[5]_net_1\, \Wt_data[5]\, 
        \r0[6]_net_1\, \Wt_data[6]\, \r0[7]_net_1\, \Wt_data[7]\, 
        \r0[8]_net_1\, \Wt_data[8]\, \r0[9]_net_1\, \Wt_data[9]\, 
        \r0[10]_net_1\, \Wt_data[10]\, \r0[11]_net_1\, 
        \Wt_data[11]\, \r0[12]_net_1\, \Wt_data[12]\, 
        \r0[13]_net_1\, \Wt_data[13]\, \r0[14]_net_1\, 
        \Wt_data[14]\, \r0[15]_net_1\, \Wt_data[15]\, 
        \r0[16]_net_1\, \Wt_data[16]\, \r0[17]_net_1\, 
        \Wt_data[17]\, \r0[18]_net_1\, \Wt_data[18]\, 
        \r0[0]_net_1\, \Wt_data[0]\, \r0[1]_net_1\, \Wt_data[1]\, 
        \r0[2]_net_1\, \Wt_data[2]\, \r0[3]_net_1\, \Wt_data[3]\, 
        \r10[23]_net_1\, \r11[23]_net_1\, \r10[24]_net_1\, 
        \r11[24]_net_1\, \r10[25]_net_1\, \r11[25]_net_1\, 
        \r10[26]_net_1\, \r11[26]_net_1\, \r10[27]_net_1\, 
        \r11[27]_net_1\, \r10[28]_net_1\, \r11[28]_net_1\, 
        \r10[29]_net_1\, \r11[29]_net_1\, \r10[30]_net_1\, 
        \r11[30]_net_1\, \r10[31]_net_1\, \r11[31]_net_1\, 
        \r10[8]_net_1\, \r11[8]_net_1\, \r10[9]_net_1\, 
        \r11[9]_net_1\, \r10[10]_net_1\, \r11[10]_net_1\, 
        \r10[11]_net_1\, \r11[11]_net_1\, \r10[12]_net_1\, 
        \r11[12]_net_1\, \r10[13]_net_1\, \r11[13]_net_1\, 
        \r10[14]_net_1\, \r11[14]_net_1\, \r10[15]_net_1\, 
        \r11[15]_net_1\, \r10[16]_net_1\, \r11[16]_net_1\, 
        \r10[17]_net_1\, \r11[17]_net_1\, \r10[18]_net_1\, 
        \r11[18]_net_1\, \r10[19]_net_1\, \r11[19]_net_1\, 
        \r10[20]_net_1\, \r11[20]_net_1\, \r10[21]_net_1\, 
        \r11[21]_net_1\, \r10[22]_net_1\, \r11[22]_net_1\, 
        \r9[25]_net_1\, \r9[26]_net_1\, \r9[27]_net_1\, 
        \r9[28]_net_1\, \r9[29]_net_1\, \r9[30]_net_1\, 
        \r9[31]_net_1\, \r10[0]_net_1\, \r11[0]_net_1\, 
        \r10[1]_net_1\, \r11[1]_net_1\, \r10[2]_net_1\, 
        \r11[2]_net_1\, \r10[3]_net_1\, \r11[3]_net_1\, 
        \r10[4]_net_1\, \r11[4]_net_1\, \r10[5]_net_1\, 
        \r11[5]_net_1\, \r10[6]_net_1\, \r11[6]_net_1\, 
        \r10[7]_net_1\, \r11[7]_net_1\, \r9[10]_net_1\, 
        \r9[11]_net_1\, \r9[12]_net_1\, \r9[13]_net_1\, 
        \r9[14]_net_1\, \r9[15]_net_1\, \r9[16]_net_1\, 
        \r9[17]_net_1\, \r9[18]_net_1\, \r9[19]_net_1\, 
        \r9[20]_net_1\, \r9[21]_net_1\, \r9[22]_net_1\, 
        \r9[23]_net_1\, \r9[24]_net_1\, \r12[27]_net_1\, 
        \r12[28]_net_1\, \r12[29]_net_1\, \r12[30]_net_1\, 
        \r12[31]_net_1\, \r9[0]_net_1\, \r9[1]_net_1\, 
        \r9[2]_net_1\, \r9[3]_net_1\, \r9[4]_net_1\, 
        \r9[5]_net_1\, \r9[6]_net_1\, \r9[7]_net_1\, 
        \r9[8]_net_1\, \r9[9]_net_1\, \r12[12]_net_1\, 
        \r12[13]_net_1\, \r12[14]_net_1\, \r12[15]_net_1\, 
        \r12[16]_net_1\, \r12[17]_net_1\, \r12[18]_net_1\, 
        \r12[19]_net_1\, \r12[20]_net_1\, \r12[21]_net_1\, 
        \r12[22]_net_1\, \r12[23]_net_1\, \r12[24]_net_1\, 
        \r12[25]_net_1\, \r12[26]_net_1\, \r12[0]_net_1\, 
        \r12[1]_net_1\, \r12[2]_net_1\, \r12[3]_net_1\, 
        \r12[4]_net_1\, \r12[5]_net_1\, \r12[6]_net_1\, 
        \r12[7]_net_1\, \r12[8]_net_1\, \r12[9]_net_1\, 
        \r12[10]_net_1\, \r12[11]_net_1\, \r8[31]_net_1\, 
        \r8[16]_net_1\, \r8[17]_net_1\, \r8[18]_net_1\, 
        \r8[19]_net_1\, \r8[20]_net_1\, \r8[21]_net_1\, 
        \r8[22]_net_1\, \r8[23]_net_1\, \r8[24]_net_1\, 
        \r8[25]_net_1\, \r8[26]_net_1\, \r8[27]_net_1\, 
        \r8[28]_net_1\, \r8[29]_net_1\, \r8[30]_net_1\, 
        \r8[1]_net_1\, \r8[2]_net_1\, \r8[3]_net_1\, 
        \r8[4]_net_1\, \r8[5]_net_1\, \r8[6]_net_1\, 
        \r8[7]_net_1\, \r8[8]_net_1\, \r8[9]_net_1\, 
        \r8[10]_net_1\, \r8[11]_net_1\, \r8[12]_net_1\, 
        \r8[13]_net_1\, \r8[14]_net_1\, \r8[15]_net_1\, 
        \r8[0]_net_1\, \next_r0_0_cry_0\, \next_r0_0_cry_0_Y\, 
        sum0_5_cry_0_Y, sum0_4_cry_0_Y, \next_r0_0_cry_1\, 
        next_r0_0_cry_1_S, \sum0_4[1]\, \sum0_5[1]\, 
        \next_r0_0_cry_2\, next_r0_0_cry_2_S, \sum0_4[2]\, 
        \sum0_5[2]\, \next_r0_0_cry_3\, next_r0_0_cry_3_S, 
        \sum0_4[3]\, \sum0_5[3]\, \next_r0_0_cry_4\, 
        next_r0_0_cry_4_S, \sum0_4[4]\, \sum0_5[4]\, 
        \next_r0_0_cry_5\, next_r0_0_cry_5_S, \sum0_4[5]\, 
        \sum0_5[5]\, \next_r0_0_cry_6\, next_r0_0_cry_6_S, 
        \sum0_4[6]\, \sum0_5[6]\, \next_r0_0_cry_7\, 
        next_r0_0_cry_7_S, \sum0_4[7]\, \sum0_5[7]\, 
        \next_r0_0_cry_8\, next_r0_0_cry_8_S, \sum0_4[8]\, 
        \sum0_5[8]\, \next_r0_0_cry_9\, next_r0_0_cry_9_S, 
        \sum0_4[9]\, \sum0_5[9]\, \next_r0_0_cry_10\, 
        next_r0_0_cry_10_S, \sum0_4[10]\, \sum0_5[10]\, 
        \next_r0_0_cry_11\, next_r0_0_cry_11_S, \sum0_4[11]\, 
        \sum0_5[11]\, \next_r0_0_cry_12\, next_r0_0_cry_12_S, 
        \sum0_4[12]\, \sum0_5[12]\, \next_r0_0_cry_13\, 
        next_r0_0_cry_13_S, \sum0_4[13]\, \sum0_5[13]\, 
        \next_r0_0_cry_14\, next_r0_0_cry_14_S, \sum0_4[14]\, 
        \sum0_5[14]\, \next_r0_0_cry_15\, next_r0_0_cry_15_S, 
        \sum0_4[15]\, \sum0_5[15]\, \next_r0_0_cry_16\, 
        next_r0_0_cry_16_S, \sum0_4[16]\, \sum0_5[16]\, 
        \next_r0_0_cry_17\, next_r0_0_cry_17_S, \sum0_4[17]\, 
        \sum0_5[17]\, \next_r0_0_cry_18\, next_r0_0_cry_18_S, 
        \sum0_4[18]\, \sum0_5[18]\, \next_r0_0_cry_19\, 
        next_r0_0_cry_19_S, \sum0_4[19]\, \sum0_5[19]\, 
        \next_r0_0_cry_20\, next_r0_0_cry_20_S, \sum0_4[20]\, 
        \sum0_5[20]\, \next_r0_0_cry_21\, next_r0_0_cry_21_S, 
        \sum0_4[21]\, \sum0_5[21]\, \next_r0_0_cry_22\, 
        next_r0_0_cry_22_S, \sum0_4[22]\, \sum0_5[22]\, 
        \next_r0_0_cry_23\, next_r0_0_cry_23_S, \sum0_4[23]\, 
        \sum0_5[23]\, \next_r0_0_cry_24\, next_r0_0_cry_24_S, 
        \sum0_4[24]\, \sum0_5[24]\, \next_r0_0_cry_25\, 
        next_r0_0_cry_25_S, \sum0_4[25]\, \sum0_5[25]\, 
        \next_r0_0_cry_26\, next_r0_0_cry_26_S, \sum0_4[26]\, 
        \sum0_5[26]\, \next_r0_0_cry_27\, next_r0_0_cry_27_S, 
        \sum0_4[27]\, \sum0_5[27]\, \next_r0_0_cry_28\, 
        next_r0_0_cry_28_S, \sum0_4[28]\, \sum0_5[28]\, 
        \next_r0_0_cry_29\, next_r0_0_cry_29_S, \sum0_4[29]\, 
        \sum0_5[29]\, next_r0_0_s_31_S, \sum0_4[31]\, 
        \sum0_5[31]\, \next_r0_0_cry_30\, next_r0_0_cry_30_S, 
        \sum0_4[30]\, \sum0_5[30]\, \sum0_4_cry_0\, \s0_0[0]\, 
        \sum0_4[0]\, \sum0_4_cry_1\, \s0_0[1]\, \sum0_4_axb_1\, 
        \sum0_4_cry_2\, \s0_0[2]\, \sum0_4_axb_2\, \sum0_4_cry_3\, 
        \s0_0[3]\, \sum0_4_axb_3\, \sum0_4_cry_4\, \s0_0[4]\, 
        \sum0_4_axb_4\, \sum0_4_cry_5\, \s0_0[5]\, \sum0_4_axb_5\, 
        \sum0_4_cry_6\, \s0_0[6]\, \sum0_4_axb_6\, \sum0_4_cry_7\, 
        \s0_0[7]\, \sum0_4_axb_7\, \sum0_4_cry_8\, \s0_0[8]\, 
        \sum0_4_axb_8\, \sum0_4_cry_9\, \s0_0[9]\, \sum0_4_axb_9\, 
        \sum0_4_cry_10\, \s0_0[10]\, \sum0_4_axb_10\, 
        \sum0_4_cry_11\, \s0_0[11]\, \sum0_4_axb_11\, 
        \sum0_4_cry_12\, \s0_0[12]\, \sum0_4_axb_12\, 
        \sum0_4_cry_13\, \s0_0[13]\, \sum0_4_axb_13\, 
        \sum0_4_cry_14\, \s0_0[14]\, \sum0_4_axb_14\, 
        \sum0_4_cry_15\, \s0_0[15]\, \sum0_4_axb_15\, 
        \sum0_4_cry_16\, \s0_0[16]\, \sum0_4_axb_16\, 
        \sum0_4_cry_17\, \s0_0[17]\, \sum0_4_axb_17\, 
        \sum0_4_cry_18\, \s0_0[18]\, \sum0_4_axb_18\, 
        \sum0_4_cry_19\, \s0_0[19]\, \sum0_4_axb_19\, 
        \sum0_4_cry_20\, \s0_0[20]\, \sum0_4_axb_20\, 
        \sum0_4_cry_21\, \s0_0[21]\, \sum0_4_axb_21\, 
        \sum0_4_cry_22\, \s0_0[22]\, \sum0_4_axb_22\, 
        \sum0_4_cry_23\, \s0_0[23]\, \sum0_4_axb_23\, 
        \sum0_4_cry_24\, \s0_0[24]\, \sum0_4_axb_24\, 
        \sum0_4_cry_25\, \s0_0[25]\, \sum0_4_axb_25\, 
        \sum0_4_cry_26\, \s0_0[26]\, \sum0_4_axb_26\, 
        \sum0_4_cry_27\, \s0_0[27]\, \sum0_4_axb_27\, 
        \sum0_4_cry_28\, \s0_0[28]\, \sum0_4_axb_28\, 
        \sum0_4_cry_29\, \s0_0[29]\, \sum0_4_axb_29\, 
        \sum0_4_cry_30\, \s0_0[30]\, \sum0_4_axb_30\, 
        \sum0_5_cry_0\, \sum0_5_cry_1\, \sum0_5_cry_2\, 
        \sum0_5_cry_3\, \sum0_5_cry_4\, \sum0_5_cry_5\, 
        \sum0_5_cry_6\, \sum0_5_cry_7\, \sum0_5_cry_8\, 
        \sum0_5_cry_9\, \sum0_5_cry_10\, \sum0_5_cry_11\, 
        \sum0_5_cry_12\, \sum0_5_cry_13\, \sum0_5_cry_14\, 
        \sum0_5_cry_15\, \sum0_5_cry_16\, \sum0_5_cry_17\, 
        \sum0_5_cry_18\, \sum0_5_cry_19\, \sum0_5_cry_20\, 
        \sum0_5_cry_21\, \sum0_5_cry_22\, \sum0_5_cry_23\, 
        \sum0_5_cry_24\, \sum0_5_cry_25\, \sum0_5_cry_26\, 
        \sum0_5_cry_27\, \sum0_5_cry_28\, \sum0_5_cry_29\, 
        \sum0_5_cry_30\, \s0[29]_net_1\, \s0[30]_net_1\, 
        \s0[5]_net_1\, \s0[4]_net_1\, \s0[3]_net_1\, 
        \s0[2]_net_1\, \s0[1]_net_1\, \s0[0]_net_1\, 
        \s0[20]_net_1\, \s0[19]_net_1\, \s0[18]_net_1\, 
        \s0[17]_net_1\, \s0[16]_net_1\, \s0[15]_net_1\, 
        \s0[14]_net_1\, \s0[13]_net_1\, \s0[12]_net_1\, 
        \s0[11]_net_1\, \s0[10]_net_1\, \s0[9]_net_1\, 
        \s0[8]_net_1\, \s0[7]_net_1\, \s0[6]_net_1\, 
        \s0[28]_net_1\, \s0[27]_net_1\, \s0[26]_net_1\, 
        \s0[25]_net_1\, \s0[24]_net_1\, \s0[23]_net_1\, 
        \s0[22]_net_1\, \s0[21]_net_1\ : std_logic;

begin 

    Wt_data(31) <= \Wt_data[31]\;
    Wt_data(30) <= \Wt_data[30]\;
    Wt_data(29) <= \Wt_data[29]\;
    Wt_data(28) <= \Wt_data[28]\;
    Wt_data(27) <= \Wt_data[27]\;
    Wt_data(26) <= \Wt_data[26]\;
    Wt_data(25) <= \Wt_data[25]\;
    Wt_data(24) <= \Wt_data[24]\;
    Wt_data(23) <= \Wt_data[23]\;
    Wt_data(22) <= \Wt_data[22]\;
    Wt_data(21) <= \Wt_data[21]\;
    Wt_data(20) <= \Wt_data[20]\;
    Wt_data(19) <= \Wt_data[19]\;
    Wt_data(18) <= \Wt_data[18]\;
    Wt_data(17) <= \Wt_data[17]\;
    Wt_data(16) <= \Wt_data[16]\;
    Wt_data(15) <= \Wt_data[15]\;
    Wt_data(14) <= \Wt_data[14]\;
    Wt_data(13) <= \Wt_data[13]\;
    Wt_data(12) <= \Wt_data[12]\;
    Wt_data(11) <= \Wt_data[11]\;
    Wt_data(10) <= \Wt_data[10]\;
    Wt_data(9) <= \Wt_data[9]\;
    Wt_data(8) <= \Wt_data[8]\;
    Wt_data(7) <= \Wt_data[7]\;
    Wt_data(6) <= \Wt_data[6]\;
    Wt_data(5) <= \Wt_data[5]\;
    Wt_data(4) <= \Wt_data[4]\;
    Wt_data(3) <= \Wt_data[3]\;
    Wt_data(2) <= \Wt_data[2]\;
    Wt_data(1) <= \Wt_data[1]\;
    Wt_data(0) <= \Wt_data[0]\;
    next_r0_0_cry_0_Y <= \next_r0_0_cry_0_Y\;

    \r4[9]\ : SLE
      port map(D => \r5[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[9]_net_1\);
    
    \r5[22]\ : SLE
      port map(D => \r6[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[22]_net_1\);
    
    \r12[21]\ : SLE
      port map(D => \r13[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[21]_net_1\);
    
    \r12[0]\ : SLE
      port map(D => \r13[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[0]_net_1\);
    
    \r10[21]\ : SLE
      port map(D => \r11[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[21]_net_1\);
    
    sum0_4_cry_0_1030 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[22]_net_1\, B => \r2[11]_net_1\, C => 
        \r2[7]_net_1\, Y => \s0_0[4]\);
    
    \r1[13]\ : SLE
      port map(D => \r2[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[13]_net_1\);
    
    sum0_4_cry_0 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[0]\, C => \sum0_4[0]\, 
        D => GND_net_1, FCI => GND_net_1, S => OPEN, Y => 
        sum0_4_cry_0_Y, FCO => \sum0_4_cry_0\);
    
    \r9[18]\ : SLE
      port map(D => \r10[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[18]_net_1\);
    
    \r6[0]\ : SLE
      port map(D => \r7[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[0]_net_1\);
    
    \r9[29]\ : SLE
      port map(D => \r10[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[29]_net_1\);
    
    \r6[9]\ : SLE
      port map(D => \r7[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[9]_net_1\);
    
    \r13[28]\ : SLE
      port map(D => \r14[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[28]_net_1\);
    
    \r3[24]\ : SLE
      port map(D => \r4[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[24]_net_1\);
    
    \r15[14]\ : SLE
      port map(D => \r0[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[14]_net_1\);
    
    \r3[18]\ : SLE
      port map(D => \r4[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[18]_net_1\);
    
    \r3[3]\ : SLE
      port map(D => \r4[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[3]_net_1\);
    
    \next_r0[14]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_278, C => next_r0_0_cry_14_S, 
        D => W_out_2_i_1_6, Y => \Wt_data[14]\);
    
    \next_r0[17]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_290, C => next_r0_0_cry_17_S, 
        D => W_out_2_i_1_9, Y => \Wt_data[17]\);
    
    \r15[12]\ : SLE
      port map(D => \r0[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[12]_net_1\);
    
    \r15[24]\ : SLE
      port map(D => \r0[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[24]_net_1\);
    
    \r5[31]\ : SLE
      port map(D => \r6[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[31]_net_1\);
    
    sum0_4_cry_20 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[20]\, C => 
        \sum0_4_axb_20\, D => GND_net_1, FCI => \sum0_4_cry_19\, 
        S => \sum0_4[20]\, Y => OPEN, FCO => \sum0_4_cry_20\);
    
    \r15[22]\ : SLE
      port map(D => \r0[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[22]_net_1\);
    
    \r15[31]\ : SLE
      port map(D => \r0[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[31]_net_1\);
    
    \r13[3]\ : SLE
      port map(D => \r14[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[3]_net_1\);
    
    \r4[17]\ : SLE
      port map(D => \r5[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[17]_net_1\);
    
    \r0[3]\ : SLE
      port map(D => \Wt_data[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[3]_net_1\);
    
    sum0_5_cry_11 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[11]_net_1\, B => \r10[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_10\, S => 
        \sum0_5[11]\, Y => OPEN, FCO => \sum0_5_cry_11\);
    
    sum0_5_cry_4 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[4]_net_1\, B => \r10[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_3\, S => 
        \sum0_5[4]\, Y => OPEN, FCO => \sum0_5_cry_4\);
    
    \r14[13]\ : SLE
      port map(D => \r15[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[13]_net_1\);
    
    \next_r0[18]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_293, C => next_r0_0_cry_18_S, 
        D => W_out_2_i_1_10, Y => \Wt_data[18]\);
    
    \r0[7]\ : SLE
      port map(D => \Wt_data[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[7]_net_1\);
    
    \r10[11]\ : SLE
      port map(D => \r11[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[11]_net_1\);
    
    \r11[0]\ : SLE
      port map(D => \r12[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[0]_net_1\);
    
    \r2[5]\ : SLE
      port map(D => \r3[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[5]_net_1\);
    
    \r5[5]\ : SLE
      port map(D => \r6[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[5]_net_1\);
    
    \r14[25]\ : SLE
      port map(D => \r15[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[25]_net_1\);
    
    next_r0_0_cry_0 : ARI1
      generic map(INIT => x"555AA")

      port map(A => sum0_5_cry_0_Y, B => sum0_4_cry_0_Y, C => 
        GND_net_1, D => GND_net_1, FCI => GND_net_1, S => OPEN, Y
         => \next_r0_0_cry_0_Y\, FCO => \next_r0_0_cry_0\);
    
    sum0_4_cry_23 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[23]\, C => 
        \sum0_4_axb_23\, D => GND_net_1, FCI => \sum0_4_cry_22\, 
        S => \sum0_4[23]\, Y => OPEN, FCO => \sum0_4_cry_23\);
    
    \r14[19]\ : SLE
      port map(D => \r15[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[19]_net_1\);
    
    \next_r0[23]\ : CFG4
      generic map(INIT => x"F5E4")

      port map(A => ld_i_i_3, B => N_307, C => next_r0_0_cry_23_S, 
        D => W_out_2_0_2_8, Y => \Wt_data[23]\);
    
    sum0_4_cry_0_1031 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[10]_net_1\, B => \r2[6]_net_1\, C => 
        \r2[21]_net_1\, Y => \s0_0[3]\);
    
    next_r0_0_cry_11 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[11]\, B => \sum0_5[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_10\, S
         => next_r0_0_cry_11_S, Y => OPEN, FCO => 
        \next_r0_0_cry_11\);
    
    \r12[9]\ : SLE
      port map(D => \r13[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[9]_net_1\);
    
    sum0_4_cry_17 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[17]\, C => 
        \sum0_4_axb_17\, D => GND_net_1, FCI => \sum0_4_cry_16\, 
        S => \sum0_4[17]\, Y => OPEN, FCO => \sum0_4_cry_17\);
    
    sum0_4_cry_0_1020 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[0]_net_1\, B => \r2[17]_net_1\, C => 
        \r2[21]_net_1\, Y => \s0_0[14]\);
    
    next_r0_0_cry_21 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[21]\, B => \sum0_5[21]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_20\, S
         => next_r0_0_cry_21_S, Y => OPEN, FCO => 
        \next_r0_0_cry_21\);
    
    \r7[17]\ : SLE
      port map(D => \r8[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[17]_net_1\);
    
    \r8[9]\ : SLE
      port map(D => \r9[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[9]_net_1\);
    
    \r0[29]\ : SLE
      port map(D => \Wt_data[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[29]_net_1\);
    
    \r13[21]\ : SLE
      port map(D => \r14[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[21]_net_1\);
    
    sum0_4_cry_0_1010 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[27]_net_1\, C => 
        \r2[10]_net_1\, Y => \s0_0[24]\);
    
    \r0[19]\ : SLE
      port map(D => \Wt_data[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[19]_net_1\);
    
    sum0_4_cry_28 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[28]\, C => 
        \sum0_4_axb_28\, D => GND_net_1, FCI => \sum0_4_cry_27\, 
        S => \sum0_4[28]\, Y => OPEN, FCO => \sum0_4_cry_28\);
    
    \s0[4]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[22]_net_1\, B => \r2[11]_net_1\, C => 
        \r2[7]_net_1\, Y => \s0[4]_net_1\);
    
    \r6[2]\ : SLE
      port map(D => \r7[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[2]_net_1\);
    
    \r4[18]\ : SLE
      port map(D => \r5[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[18]_net_1\);
    
    sum0_4_cry_0_1008 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[12]_net_1\, B => \r2[1]_net_1\, C => 
        \r2[29]_net_1\, Y => \s0_0[26]\);
    
    \r1[24]\ : SLE
      port map(D => \r2[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[24]_net_1\);
    
    \r5[14]\ : SLE
      port map(D => \r6[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[14]_net_1\);
    
    \s0[5]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[23]_net_1\, B => \r2[12]_net_1\, C => 
        \r2[8]_net_1\, Y => \s0[5]_net_1\);
    
    \r5[8]\ : SLE
      port map(D => \r6[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[8]_net_1\);
    
    \r7[26]\ : SLE
      port map(D => \r8[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[26]_net_1\);
    
    \r4[24]\ : SLE
      port map(D => \r5[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[24]_net_1\);
    
    \r15[16]\ : SLE
      port map(D => \r0[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[16]_net_1\);
    
    \r14[14]\ : SLE
      port map(D => \r15[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[14]_net_1\);
    
    \s0[6]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[24]_net_1\, B => \r2[13]_net_1\, C => 
        \r2[9]_net_1\, Y => \s0[6]_net_1\);
    
    \r15[3]\ : SLE
      port map(D => \r0[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[3]_net_1\);
    
    \r15[26]\ : SLE
      port map(D => \r0[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[26]_net_1\);
    
    \r14[12]\ : SLE
      port map(D => \r15[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[12]_net_1\);
    
    \s0[25]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[11]_net_1\, B => \r2[0]_net_1\, C => 
        \r2[28]_net_1\, Y => \s0[25]_net_1\);
    
    \r9[15]\ : SLE
      port map(D => \r10[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[15]_net_1\);
    
    \s0[15]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[18]_net_1\, B => \r2[1]_net_1\, C => 
        \r2[22]_net_1\, Y => \s0[15]_net_1\);
    
    \r8[29]\ : SLE
      port map(D => \r9[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[29]_net_1\);
    
    \r1[17]\ : SLE
      port map(D => \r2[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[17]_net_1\);
    
    \r2[14]\ : SLE
      port map(D => \r3[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[14]_net_1\);
    
    \r11[8]\ : SLE
      port map(D => \r12[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[8]_net_1\);
    
    \r11[2]\ : SLE
      port map(D => \r12[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[2]_net_1\);
    
    \r7[21]\ : SLE
      port map(D => \r8[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[21]_net_1\);
    
    \r6[26]\ : SLE
      port map(D => \r7[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[26]_net_1\);
    
    \r3[15]\ : SLE
      port map(D => \r4[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[15]_net_1\);
    
    sum0_5_cry_30 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[30]_net_1\, B => \r10[30]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_29\, S => 
        \sum0_5[30]\, Y => OPEN, FCO => \sum0_5_cry_30\);
    
    \r11[30]\ : SLE
      port map(D => \r12[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[30]_net_1\);
    
    \r7[18]\ : SLE
      port map(D => \r8[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[18]_net_1\);
    
    \r13[30]\ : SLE
      port map(D => \r14[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[30]_net_1\);
    
    \r4[5]\ : SLE
      port map(D => \r5[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[5]_net_1\);
    
    next_r0_0_cry_18 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[18]\, B => \sum0_5[18]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_17\, S
         => next_r0_0_cry_18_S, Y => OPEN, FCO => 
        \next_r0_0_cry_18\);
    
    sum0_4_cry_0_1021 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[20]_net_1\, C => 
        \r2[16]_net_1\, Y => \s0_0[13]\);
    
    \r7[3]\ : SLE
      port map(D => \r8[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[3]_net_1\);
    
    next_r0_0_cry_28 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[28]\, B => \sum0_5[28]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_27\, S
         => next_r0_0_cry_28_S, Y => OPEN, FCO => 
        \next_r0_0_cry_28\);
    
    sum0_4_cry_0_1011 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[30]_net_1\, B => \r2[26]_net_1\, C => 
        \r2[9]_net_1\, Y => \s0_0[23]\);
    
    \r6[21]\ : SLE
      port map(D => \r7[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[21]_net_1\);
    
    \r14[27]\ : SLE
      port map(D => \r15[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[27]_net_1\);
    
    \r8[31]\ : SLE
      port map(D => \r9[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[31]_net_1\);
    
    \r2[1]\ : SLE
      port map(D => \r3[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[1]_net_1\);
    
    sum0_4_axb_28 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[13]_net_1\, B => \s0[28]_net_1\, C => 
        \r15[15]_net_1\, Y => \sum0_4_axb_28\);
    
    \r12[6]\ : SLE
      port map(D => \r13[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[6]_net_1\);
    
    sum0_5_cry_6 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[6]_net_1\, B => \r10[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_5\, S => 
        \sum0_5[6]\, Y => OPEN, FCO => \sum0_5_cry_6\);
    
    sum0_4_cry_14 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[14]\, C => 
        \sum0_4_axb_14\, D => GND_net_1, FCI => \sum0_4_cry_13\, 
        S => \sum0_4[14]\, Y => OPEN, FCO => \sum0_4_cry_14\);
    
    \r9[24]\ : SLE
      port map(D => \r10[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[24]_net_1\);
    
    \r8[10]\ : SLE
      port map(D => \r9[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[10]_net_1\);
    
    \r6[3]\ : SLE
      port map(D => \r7[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[3]_net_1\);
    
    \r8[3]\ : SLE
      port map(D => \r9[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[3]_net_1\);
    
    \s0[8]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[26]_net_1\, B => \r2[15]_net_1\, C => 
        \r2[11]_net_1\, Y => \s0[8]_net_1\);
    
    \r7[23]\ : SLE
      port map(D => \r8[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[23]_net_1\);
    
    \r15[5]\ : SLE
      port map(D => \r0[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[5]_net_1\);
    
    \r9[12]\ : SLE
      port map(D => \r10[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[12]_net_1\);
    
    \r1[18]\ : SLE
      port map(D => \r2[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[18]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    sum0_4_cry_29 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[29]\, C => 
        \sum0_4_axb_29\, D => GND_net_1, FCI => \sum0_4_cry_28\, 
        S => \sum0_4[29]\, Y => OPEN, FCO => \sum0_4_cry_29\);
    
    sum0_5_cry_21 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[21]_net_1\, B => \r10[21]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_20\, S => 
        \sum0_5[21]\, Y => OPEN, FCO => \sum0_5_cry_21\);
    
    \next_r0[13]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_275, C => next_r0_0_cry_13_S, 
        D => W_out_2_i_1_5, Y => \Wt_data[13]\);
    
    \r3[12]\ : SLE
      port map(D => \r4[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[12]_net_1\);
    
    \r6[16]\ : SLE
      port map(D => \r7[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[16]_net_1\);
    
    \r2[2]\ : SLE
      port map(D => \r3[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[2]_net_1\);
    
    \r14[16]\ : SLE
      port map(D => \r15[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[16]_net_1\);
    
    \r2[26]\ : SLE
      port map(D => \r3[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[26]_net_1\);
    
    \r9[0]\ : SLE
      port map(D => \r10[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[0]_net_1\);
    
    \r6[23]\ : SLE
      port map(D => \r7[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[23]_net_1\);
    
    sum0_4_cry_26 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[26]\, C => 
        \sum0_4_axb_26\, D => GND_net_1, FCI => \sum0_4_cry_25\, 
        S => \sum0_4[26]\, Y => OPEN, FCO => \sum0_4_cry_26\);
    
    sum0_5_cry_10 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[10]_net_1\, B => \r10[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_9\, S => 
        \sum0_5[10]\, Y => OPEN, FCO => \sum0_5_cry_10\);
    
    \s0[26]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[12]_net_1\, B => \r2[1]_net_1\, C => 
        \r2[29]_net_1\, Y => \s0[26]_net_1\);
    
    \r4[15]\ : SLE
      port map(D => \r5[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[15]_net_1\);
    
    \r9[30]\ : SLE
      port map(D => \r10[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[30]_net_1\);
    
    \s0[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[18]_net_1\, B => \r2[7]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0[0]_net_1\);
    
    \s0[16]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[19]_net_1\, B => \r2[2]_net_1\, C => 
        \r2[23]_net_1\, Y => \s0[16]_net_1\);
    
    \s0[20]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[23]_net_1\, B => \r2[6]_net_1\, C => 
        \r2[27]_net_1\, Y => \s0[20]_net_1\);
    
    \r7[0]\ : SLE
      port map(D => \r8[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[0]_net_1\);
    
    \r2[6]\ : SLE
      port map(D => \r3[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[6]_net_1\);
    
    \s0[10]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[28]_net_1\, B => \r2[13]_net_1\, C => 
        \r2[17]_net_1\, Y => \s0[10]_net_1\);
    
    \r6[11]\ : SLE
      port map(D => \r7[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[11]_net_1\);
    
    sum0_4_cry_0_1004 : CFG2
      generic map(INIT => x"6")

      port map(A => \r2[5]_net_1\, B => \r2[16]_net_1\, Y => 
        \s0_0[30]\);
    
    sum0_4_axb_6 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[16]_net_1\, B => \s0[6]_net_1\, C => 
        \r15[25]_net_1\, D => \r15[23]_net_1\, Y => 
        \sum0_4_axb_6\);
    
    \r3[26]\ : SLE
      port map(D => \r4[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[26]_net_1\);
    
    \r13[10]\ : SLE
      port map(D => \r14[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[10]_net_1\);
    
    \r12[10]\ : SLE
      port map(D => \r13[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[10]_net_1\);
    
    \r11[28]\ : SLE
      port map(D => \r12[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[28]_net_1\);
    
    \next_r0[8]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_260, C => next_r0_0_cry_8_S, 
        D => W_out_2_i_1_0, Y => \Wt_data[8]\);
    
    \r2[21]\ : SLE
      port map(D => \r3[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[21]_net_1\);
    
    \r3[9]\ : SLE
      port map(D => \r4[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[9]_net_1\);
    
    \r5[20]\ : SLE
      port map(D => \r6[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[20]_net_1\);
    
    \r11[18]\ : SLE
      port map(D => \r12[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[18]_net_1\);
    
    \r0[24]\ : SLE
      port map(D => \Wt_data[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[24]_net_1\);
    
    \r13[5]\ : SLE
      port map(D => \r14[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[5]_net_1\);
    
    \r0[14]\ : SLE
      port map(D => \Wt_data[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[14]_net_1\);
    
    sum0_5_cry_13 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[13]_net_1\, B => \r10[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_12\, S => 
        \sum0_5[13]\, Y => OPEN, FCO => \sum0_5_cry_13\);
    
    \r1[2]\ : SLE
      port map(D => \r2[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[2]_net_1\);
    
    \r3[21]\ : SLE
      port map(D => \r4[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[21]_net_1\);
    
    \r11[5]\ : SLE
      port map(D => \r12[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[5]_net_1\);
    
    \r7[15]\ : SLE
      port map(D => \r8[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[15]_net_1\);
    
    sum0_4_cry_22 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[22]\, C => 
        \sum0_4_axb_22\, D => GND_net_1, FCI => \sum0_4_cry_21\, 
        S => \sum0_4[22]\, Y => OPEN, FCO => \sum0_4_cry_22\);
    
    \r1[0]\ : SLE
      port map(D => \r2[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[0]_net_1\);
    
    \r0[1]\ : SLE
      port map(D => \Wt_data[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[1]_net_1\);
    
    \next_r0[5]\ : CFG4
      generic map(INIT => x"AFAC")

      port map(A => next_r0_0_cry_5_S, B => N_349, C => ld_i_i_3, 
        D => W_out_2_0(5), Y => \Wt_data[5]\);
    
    \r14[23]\ : SLE
      port map(D => \r15[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[23]_net_1\);
    
    sum0_5_cry_18 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[18]_net_1\, B => \r10[18]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_17\, S => 
        \sum0_5[18]\, Y => OPEN, FCO => \sum0_5_cry_18\);
    
    \r6[13]\ : SLE
      port map(D => \r7[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[13]_net_1\);
    
    \r1[5]\ : SLE
      port map(D => \r2[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[5]_net_1\);
    
    \r4[12]\ : SLE
      port map(D => \r5[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[12]_net_1\);
    
    \r2[23]\ : SLE
      port map(D => \r3[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[23]_net_1\);
    
    \next_r0[29]\ : CFG4
      generic map(INIT => x"C0D1")

      port map(A => W_out_2_i_1_21, B => ld_i_i_3, C => 
        next_r0_0_cry_29_S, D => W_out_2_i_0(29), Y => 
        \Wt_data[29]\);
    
    \r8[24]\ : SLE
      port map(D => \r9[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[24]_net_1\);
    
    \r5[0]\ : SLE
      port map(D => \r6[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[0]_net_1\);
    
    \r6[7]\ : SLE
      port map(D => \r7[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[7]_net_1\);
    
    sum0_4_cry_0_1009 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[11]_net_1\, B => \r2[0]_net_1\, C => 
        \r2[28]_net_1\, Y => \s0_0[25]\);
    
    next_r0_0_cry_13 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[13]\, B => \sum0_5[13]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_12\, S
         => next_r0_0_cry_13_S, Y => OPEN, FCO => 
        \next_r0_0_cry_13\);
    
    \r9[7]\ : SLE
      port map(D => \r10[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[7]_net_1\);
    
    next_r0_0_cry_23 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[23]\, B => \sum0_5[23]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_22\, S
         => next_r0_0_cry_23_S, Y => OPEN, FCO => 
        \next_r0_0_cry_23\);
    
    \r14[29]\ : SLE
      port map(D => \r15[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[29]_net_1\);
    
    \next_r0[1]\ : CFG4
      generic map(INIT => x"C0E2")

      port map(A => N_98, B => ld_i_i_3, C => next_r0_0_cry_1_S, 
        D => W_out_i_1(1), Y => \Wt_data[1]\);
    
    sum0_5_s_31 : ARI1
      generic map(INIT => x"46600")

      port map(A => VCC_net_1, B => \r1[31]_net_1\, C => 
        \r10[31]_net_1\, D => GND_net_1, FCI => \sum0_5_cry_30\, 
        S => \sum0_5[31]\, Y => OPEN, FCO => OPEN);
    
    \r3[1]\ : SLE
      port map(D => \r4[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[1]_net_1\);
    
    \next_r0[6]\ : CFG4
      generic map(INIT => x"AFAC")

      port map(A => next_r0_0_cry_6_S, B => N_251, C => ld_i_i_3, 
        D => W_out_2_0_0_3, Y => \Wt_data[6]\);
    
    \r3[23]\ : SLE
      port map(D => \r4[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[23]_net_1\);
    
    \r11[21]\ : SLE
      port map(D => \r12[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[21]_net_1\);
    
    \r7[27]\ : SLE
      port map(D => \r8[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[27]_net_1\);
    
    \next_r0[22]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_305, C => next_r0_0_cry_22_S, 
        D => W_out_2_i_1_14, Y => \Wt_data[22]\);
    
    \r1[15]\ : SLE
      port map(D => \r2[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[15]_net_1\);
    
    \r11[11]\ : SLE
      port map(D => \r12[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[11]_net_1\);
    
    \r9[4]\ : SLE
      port map(D => \r10[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[4]_net_1\);
    
    \r1[26]\ : SLE
      port map(D => \r2[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[26]_net_1\);
    
    \r5[16]\ : SLE
      port map(D => \r6[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[16]_net_1\);
    
    \r3[31]\ : SLE
      port map(D => \r4[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[31]_net_1\);
    
    \r4[26]\ : SLE
      port map(D => \r5[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[26]_net_1\);
    
    \r7[12]\ : SLE
      port map(D => \r8[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[12]_net_1\);
    
    \next_r0[30]\ : CFG4
      generic map(INIT => x"C0D1")

      port map(A => W_out_2_i_1_22, B => ld_i_i_3, C => 
        next_r0_0_cry_30_S, D => W_out_2_i_0(30), Y => 
        \Wt_data[30]\);
    
    \r10[6]\ : SLE
      port map(D => \r11[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[6]_net_1\);
    
    next_r0_0_cry_4 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[4]\, B => \sum0_5[4]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_3\, S => 
        next_r0_0_cry_4_S, Y => OPEN, FCO => \next_r0_0_cry_4\);
    
    \r13[15]\ : SLE
      port map(D => \r14[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[15]_net_1\);
    
    \r12[15]\ : SLE
      port map(D => \r13[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[15]_net_1\);
    
    \r9[5]\ : SLE
      port map(D => \r10[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[5]_net_1\);
    
    \r8[19]\ : SLE
      port map(D => \r9[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[19]_net_1\);
    
    \r6[27]\ : SLE
      port map(D => \r7[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[27]_net_1\);
    
    \r14[24]\ : SLE
      port map(D => \r15[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[24]_net_1\);
    
    \r2[30]\ : SLE
      port map(D => \r3[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[30]_net_1\);
    
    \r14[22]\ : SLE
      port map(D => \r15[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[22]_net_1\);
    
    \r2[4]\ : SLE
      port map(D => \r3[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[4]_net_1\);
    
    \r2[16]\ : SLE
      port map(D => \r3[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[16]_net_1\);
    
    \r1[21]\ : SLE
      port map(D => \r2[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[21]_net_1\);
    
    \r5[11]\ : SLE
      port map(D => \r6[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[11]_net_1\);
    
    \r12[5]\ : SLE
      port map(D => \r13[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[5]_net_1\);
    
    \r15[18]\ : SLE
      port map(D => \r0[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[18]_net_1\);
    
    \r4[21]\ : SLE
      port map(D => \r5[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[21]_net_1\);
    
    \r11[9]\ : SLE
      port map(D => \r12[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[9]_net_1\);
    
    \r15[28]\ : SLE
      port map(D => \r0[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[28]_net_1\);
    
    \r7[5]\ : SLE
      port map(D => \r8[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[5]_net_1\);
    
    \r9[2]\ : SLE
      port map(D => \r10[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[2]_net_1\);
    
    \r4[7]\ : SLE
      port map(D => \r5[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[7]_net_1\);
    
    sum0_4_cry_1 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[1]\, C => 
        \sum0_4_axb_1\, D => GND_net_1, FCI => \sum0_4_cry_0\, S
         => \sum0_4[1]\, Y => OPEN, FCO => \sum0_4_cry_1\);
    
    sum0_4_cry_15 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[15]\, C => 
        \sum0_4_axb_15\, D => GND_net_1, FCI => \sum0_4_cry_14\, 
        S => \sum0_4[15]\, Y => OPEN, FCO => \sum0_4_cry_15\);
    
    \r7[28]\ : SLE
      port map(D => \r8[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[28]_net_1\);
    
    sum0_5_cry_20 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[20]_net_1\, B => \r10[20]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_19\, S => 
        \sum0_5[20]\, Y => OPEN, FCO => \sum0_5_cry_20\);
    
    \r1[12]\ : SLE
      port map(D => \r2[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[12]_net_1\);
    
    \next_r0[3]\ : CFG4
      generic map(INIT => x"AFAC")

      port map(A => next_r0_0_cry_3_S, B => N_245, C => ld_i_i_3, 
        D => W_out_2_0_0_0, Y => \Wt_data[3]\);
    
    \r8[4]\ : SLE
      port map(D => \r9[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[4]_net_1\);
    
    \r2[11]\ : SLE
      port map(D => \r3[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[11]_net_1\);
    
    sum0_5_cry_19 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[19]_net_1\, B => \r10[19]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_18\, S => 
        \sum0_5[19]\, Y => OPEN, FCO => \sum0_5_cry_19\);
    
    \r7[4]\ : SLE
      port map(D => \r8[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[4]_net_1\);
    
    \r6[6]\ : SLE
      port map(D => \r7[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[6]_net_1\);
    
    \r9[26]\ : SLE
      port map(D => \r10[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[26]_net_1\);
    
    \r10[9]\ : SLE
      port map(D => \r11[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[9]_net_1\);
    
    sum0_4_cry_7 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[7]\, C => 
        \sum0_4_axb_7\, D => GND_net_1, FCI => \sum0_4_cry_6\, S
         => \sum0_4[7]\, Y => OPEN, FCO => \sum0_4_cry_7\);
    
    \r4[3]\ : SLE
      port map(D => \r5[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[3]_net_1\);
    
    \r1[23]\ : SLE
      port map(D => \r2[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[23]_net_1\);
    
    sum0_5_cry_16 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[16]_net_1\, B => \r10[16]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_15\, S => 
        \sum0_5[16]\, Y => OPEN, FCO => \sum0_5_cry_16\);
    
    \r5[13]\ : SLE
      port map(D => \r6[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[13]_net_1\);
    
    \s0[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[27]_net_1\, B => \r2[16]_net_1\, C => 
        \r2[12]_net_1\, Y => \s0[9]_net_1\);
    
    \r4[23]\ : SLE
      port map(D => \r5[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[23]_net_1\);
    
    \r14[3]\ : SLE
      port map(D => \r15[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[3]_net_1\);
    
    next_r0_0_cry_5 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[5]\, B => \sum0_5[5]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_4\, S => 
        next_r0_0_cry_5_S, Y => OPEN, FCO => \next_r0_0_cry_5\);
    
    \s0[21]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[28]_net_1\, B => \r2[24]_net_1\, C => 
        \r2[7]_net_1\, Y => \s0[21]_net_1\);
    
    \r6[28]\ : SLE
      port map(D => \r7[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[28]_net_1\);
    
    sum0_4_cry_0_1007 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[13]_net_1\, B => \r2[2]_net_1\, C => 
        \r2[30]_net_1\, Y => \s0_0[27]\);
    
    \r6[17]\ : SLE
      port map(D => \r7[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[17]_net_1\);
    
    \r5[29]\ : SLE
      port map(D => \r6[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[29]_net_1\);
    
    \next_r0[19]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_296, C => next_r0_0_cry_19_S, 
        D => W_out_2_i_1_11, Y => \Wt_data[19]\);
    
    \s0[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[29]_net_1\, B => \r2[18]_net_1\, C => 
        \r2[14]_net_1\, Y => \s0[11]_net_1\);
    
    sum0_4_axb_18 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[3]_net_1\, B => \r15[5]_net_1\, C => 
        \s0[18]_net_1\, D => \r15[28]_net_1\, Y => 
        \sum0_4_axb_18\);
    
    \r5[7]\ : SLE
      port map(D => \r6[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[7]_net_1\);
    
    \r2[27]\ : SLE
      port map(D => \r3[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[27]_net_1\);
    
    sum0_5_cry_23 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[23]_net_1\, B => \r10[23]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_22\, S => 
        \sum0_5[23]\, Y => OPEN, FCO => \sum0_5_cry_23\);
    
    \r4[31]\ : SLE
      port map(D => \r5[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[31]_net_1\);
    
    \r2[8]\ : SLE
      port map(D => \r3[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[8]_net_1\);
    
    \r2[3]\ : SLE
      port map(D => \r3[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[3]_net_1\);
    
    \r9[21]\ : SLE
      port map(D => \r10[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[21]_net_1\);
    
    \r2[13]\ : SLE
      port map(D => \r3[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[13]_net_1\);
    
    \r13[17]\ : SLE
      port map(D => \r14[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[17]_net_1\);
    
    \r12[17]\ : SLE
      port map(D => \r13[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[17]_net_1\);
    
    \r15[11]\ : SLE
      port map(D => \r0[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[11]_net_1\);
    
    \r9[10]\ : SLE
      port map(D => \r10[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[10]_net_1\);
    
    \r14[26]\ : SLE
      port map(D => \r15[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[26]_net_1\);
    
    \s0[23]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[30]_net_1\, B => \r2[26]_net_1\, C => 
        \r2[9]_net_1\, Y => \s0[23]_net_1\);
    
    sum0_4_s_31 : ARI1
      generic map(INIT => x"46996")

      port map(A => \r15[18]_net_1\, B => \r2[6]_net_1\, C => 
        \r2[17]_net_1\, D => \r15[16]_net_1\, FCI => 
        \sum0_4_cry_30\, S => \sum0_4[31]\, Y => OPEN, FCO => 
        OPEN);
    
    \r13[2]\ : SLE
      port map(D => \r14[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[2]_net_1\);
    
    sum0_5_cry_28 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[28]_net_1\, B => \r10[28]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_27\, S => 
        \sum0_5[28]\, Y => OPEN, FCO => \sum0_5_cry_28\);
    
    \r14[9]\ : SLE
      port map(D => \r15[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[9]_net_1\);
    
    \s0[13]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[20]_net_1\, C => 
        \r2[16]_net_1\, Y => \s0[13]_net_1\);
    
    \r3[27]\ : SLE
      port map(D => \r4[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[27]_net_1\);
    
    \next_r0[12]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_273, C => next_r0_0_cry_12_S, 
        D => W_out_2_i_1_4, Y => \Wt_data[12]\);
    
    \r15[21]\ : SLE
      port map(D => \r0[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[21]_net_1\);
    
    sum0_4_cry_6 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[6]\, C => 
        \sum0_4_axb_6\, D => GND_net_1, FCI => \sum0_4_cry_5\, S
         => \sum0_4[6]\, Y => OPEN, FCO => \sum0_4_cry_6\);
    
    \r13[6]\ : SLE
      port map(D => \r14[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[6]_net_1\);
    
    \r6[5]\ : SLE
      port map(D => \r7[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[5]_net_1\);
    
    \r3[10]\ : SLE
      port map(D => \r4[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[10]_net_1\);
    
    \r3[7]\ : SLE
      port map(D => \r4[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[7]_net_1\);
    
    \r11[3]\ : SLE
      port map(D => \r12[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[3]_net_1\);
    
    sum0_5_cry_12 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[12]_net_1\, B => \r10[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_11\, S => 
        \sum0_5[12]\, Y => OPEN, FCO => \sum0_5_cry_12\);
    
    \r14[18]\ : SLE
      port map(D => \r15[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[18]_net_1\);
    
    \r9[3]\ : SLE
      port map(D => \r10[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[3]_net_1\);
    
    \r14[5]\ : SLE
      port map(D => \r15[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[5]_net_1\);
    
    \r12[20]\ : SLE
      port map(D => \r13[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[20]_net_1\);
    
    \r10[20]\ : SLE
      port map(D => \r11[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[20]_net_1\);
    
    \r9[23]\ : SLE
      port map(D => \r10[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[23]_net_1\);
    
    \r0[26]\ : SLE
      port map(D => \Wt_data[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[26]_net_1\);
    
    \r15[2]\ : SLE
      port map(D => \r0[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[2]_net_1\);
    
    \r6[18]\ : SLE
      port map(D => \r7[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[18]_net_1\);
    
    \r0[16]\ : SLE
      port map(D => \Wt_data[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[16]_net_1\);
    
    \r2[28]\ : SLE
      port map(D => \r3[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[28]_net_1\);
    
    \r6[30]\ : SLE
      port map(D => \r7[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[30]_net_1\);
    
    \r12[8]\ : SLE
      port map(D => \r13[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[8]_net_1\);
    
    sum0_4_cry_27 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[27]\, C => 
        \sum0_4_axb_27\, D => GND_net_1, FCI => \sum0_4_cry_26\, 
        S => \sum0_4[27]\, Y => OPEN, FCO => \sum0_4_cry_27\);
    
    sum0_4_cry_0_1025 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[27]_net_1\, B => \r2[16]_net_1\, C => 
        \r2[12]_net_1\, Y => \s0_0[9]\);
    
    sum0_4_axb_26 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[11]_net_1\, B => \s0[26]_net_1\, C => 
        \r15[13]_net_1\, Y => \sum0_4_axb_26\);
    
    \r1[1]\ : SLE
      port map(D => \r2[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[1]_net_1\);
    
    sum0_4_cry_4 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[4]\, C => 
        \sum0_4_axb_4\, D => GND_net_1, FCI => \sum0_4_cry_3\, S
         => \sum0_4[4]\, Y => OPEN, FCO => \sum0_4_cry_4\);
    
    \r7[25]\ : SLE
      port map(D => \r8[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[25]_net_1\);
    
    \r0[21]\ : SLE
      port map(D => \Wt_data[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[21]_net_1\);
    
    \r1[4]\ : SLE
      port map(D => \r2[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[4]_net_1\);
    
    \r15[30]\ : SLE
      port map(D => \r0[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[30]_net_1\);
    
    sum0_4_axb_29 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[14]_net_1\, B => \s0[29]_net_1\, C => 
        \r15[16]_net_1\, Y => \sum0_4_axb_29\);
    
    \r13[4]\ : SLE
      port map(D => \r14[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[4]_net_1\);
    
    sum0_4_cry_0_1015 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[26]_net_1\, B => \r2[22]_net_1\, C => 
        \r2[5]_net_1\, Y => \s0_0[19]\);
    
    \r8[14]\ : SLE
      port map(D => \r9[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[14]_net_1\);
    
    \r0[11]\ : SLE
      port map(D => \Wt_data[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[11]_net_1\);
    
    \r3[28]\ : SLE
      port map(D => \r4[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[28]_net_1\);
    
    \r8[26]\ : SLE
      port map(D => \r9[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[26]_net_1\);
    
    sum0_4_cry_8 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[8]\, C => 
        \sum0_4_axb_8\, D => GND_net_1, FCI => \sum0_4_cry_7\, S
         => \sum0_4[8]\, Y => OPEN, FCO => \sum0_4_cry_8\);
    
    \r12[2]\ : SLE
      port map(D => \r13[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[2]_net_1\);
    
    \r10[2]\ : SLE
      port map(D => \r11[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[2]_net_1\);
    
    sum0_4_cry_3 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[3]\, C => 
        \sum0_4_axb_3\, D => GND_net_1, FCI => \sum0_4_cry_2\, S
         => \sum0_4[3]\, Y => OPEN, FCO => \sum0_4_cry_3\);
    
    \r7[9]\ : SLE
      port map(D => \r8[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[9]_net_1\);
    
    \r10[10]\ : SLE
      port map(D => \r11[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[10]_net_1\);
    
    \r10[8]\ : SLE
      port map(D => \r11[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[8]_net_1\);
    
    \r6[25]\ : SLE
      port map(D => \r7[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[25]_net_1\);
    
    \r4[10]\ : SLE
      port map(D => \r5[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[10]_net_1\);
    
    \r1[27]\ : SLE
      port map(D => \r2[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[27]_net_1\);
    
    \r14[31]\ : SLE
      port map(D => \r15[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[31]_net_1\);
    
    \r14[11]\ : SLE
      port map(D => \r15[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[11]_net_1\);
    
    \r5[17]\ : SLE
      port map(D => \r6[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[17]_net_1\);
    
    \r4[27]\ : SLE
      port map(D => \r5[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[27]_net_1\);
    
    \r13[13]\ : SLE
      port map(D => \r14[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[13]_net_1\);
    
    \r12[13]\ : SLE
      port map(D => \r13[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[13]_net_1\);
    
    next_r0_0_cry_14 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[14]\, B => \sum0_5[14]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_13\, S
         => next_r0_0_cry_14_S, Y => OPEN, FCO => 
        \next_r0_0_cry_14\);
    
    sum0_4_axb_21 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[6]_net_1\, B => \r15[8]_net_1\, C => 
        \s0[21]_net_1\, D => \r15[31]_net_1\, Y => 
        \sum0_4_axb_21\);
    
    \r8[21]\ : SLE
      port map(D => \r9[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[21]_net_1\);
    
    \r0[23]\ : SLE
      port map(D => \Wt_data[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[23]_net_1\);
    
    next_r0_0_cry_24 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[24]\, B => \sum0_5[24]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_23\, S
         => next_r0_0_cry_24_S, Y => OPEN, FCO => 
        \next_r0_0_cry_24\);
    
    \r14[4]\ : SLE
      port map(D => \r15[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[4]_net_1\);
    
    sum0_5_cry_29 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[29]_net_1\, B => \r10[29]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_28\, S => 
        \sum0_5[29]\, Y => OPEN, FCO => \sum0_5_cry_29\);
    
    \r0[13]\ : SLE
      port map(D => \Wt_data[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[13]_net_1\);
    
    \r13[20]\ : SLE
      port map(D => \r14[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[20]_net_1\);
    
    \r13[1]\ : SLE
      port map(D => \r14[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[1]_net_1\);
    
    \r12[25]\ : SLE
      port map(D => \r13[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[25]_net_1\);
    
    \r10[25]\ : SLE
      port map(D => \r11[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[25]_net_1\);
    
    \r2[17]\ : SLE
      port map(D => \r3[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[17]_net_1\);
    
    sum0_5_cry_26 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[26]_net_1\, B => \r10[26]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_25\, S => 
        \sum0_5[26]\, Y => OPEN, FCO => \sum0_5_cry_26\);
    
    \r7[22]\ : SLE
      port map(D => \r8[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[22]_net_1\);
    
    \r14[1]\ : SLE
      port map(D => \r15[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[1]_net_1\);
    
    \r8[6]\ : SLE
      port map(D => \r9[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[6]_net_1\);
    
    \r1[30]\ : SLE
      port map(D => \r2[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[30]_net_1\);
    
    \r15[9]\ : SLE
      port map(D => \r0[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[9]_net_1\);
    
    \r13[19]\ : SLE
      port map(D => \r14[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[19]_net_1\);
    
    \r12[19]\ : SLE
      port map(D => \r13[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[19]_net_1\);
    
    sum0_4_axb_30 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[15]_net_1\, B => \s0[30]_net_1\, C => 
        \r15[17]_net_1\, Y => \sum0_4_axb_30\);
    
    \r2[0]\ : SLE
      port map(D => \r3[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[0]_net_1\);
    
    \r5[24]\ : SLE
      port map(D => \r6[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[24]_net_1\);
    
    \r7[31]\ : SLE
      port map(D => \r8[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[31]_net_1\);
    
    sum0_5_cry_7 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[7]_net_1\, B => \r10[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_6\, S => 
        \sum0_5[7]\, Y => OPEN, FCO => \sum0_5_cry_7\);
    
    \r7[10]\ : SLE
      port map(D => \r8[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[10]_net_1\);
    
    \s0[3]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[10]_net_1\, B => \r2[6]_net_1\, C => 
        \r2[21]_net_1\, Y => \s0[3]_net_1\);
    
    \next_r0[31]\ : CFG4
      generic map(INIT => x"AFAC")

      port map(A => next_r0_0_s_31_S, B => W_out_i_i_2(31), C => 
        ld_i_i_3, D => W_out_i_i_1(31), Y => \Wt_data[31]\);
    
    sum0_4_cry_24 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[24]\, C => 
        \sum0_4_axb_24\, D => GND_net_1, FCI => \sum0_4_cry_23\, 
        S => \sum0_4[24]\, Y => OPEN, FCO => \sum0_4_cry_24\);
    
    \r4[0]\ : SLE
      port map(D => \r5[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[0]_net_1\);
    
    \r15[8]\ : SLE
      port map(D => \r0[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[8]_net_1\);
    
    \r8[23]\ : SLE
      port map(D => \r9[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[23]_net_1\);
    
    sum0_4_axb_22 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[7]_net_1\, B => \s0[22]_net_1\, C => 
        \r15[9]_net_1\, Y => \sum0_4_axb_22\);
    
    \r10[31]\ : SLE
      port map(D => \r11[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[31]_net_1\);
    
    \r6[22]\ : SLE
      port map(D => \r7[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[22]_net_1\);
    
    \r10[5]\ : SLE
      port map(D => \r11[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[5]_net_1\);
    
    \r1[28]\ : SLE
      port map(D => \r2[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[28]_net_1\);
    
    \r6[15]\ : SLE
      port map(D => \r7[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[15]_net_1\);
    
    \r5[18]\ : SLE
      port map(D => \r6[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[18]_net_1\);
    
    \s0[7]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[25]_net_1\, B => \r2[14]_net_1\, C => 
        \r2[10]_net_1\, Y => \s0[7]_net_1\);
    
    \r0[2]\ : SLE
      port map(D => \Wt_data[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[2]_net_1\);
    
    \r4[28]\ : SLE
      port map(D => \r5[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[28]_net_1\);
    
    \r2[25]\ : SLE
      port map(D => \r3[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[25]_net_1\);
    
    \r11[6]\ : SLE
      port map(D => \r12[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[6]_net_1\);
    
    \r9[27]\ : SLE
      port map(D => \r10[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[27]_net_1\);
    
    sum0_4_axb_25 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[10]_net_1\, B => \s0[25]_net_1\, C => 
        \r15[12]_net_1\, Y => \sum0_4_axb_25\);
    
    \r9[19]\ : SLE
      port map(D => \r10[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[19]_net_1\);
    
    \r12[31]\ : SLE
      port map(D => \r13[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[31]_net_1\);
    
    \r13[14]\ : SLE
      port map(D => \r14[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[14]_net_1\);
    
    \r12[14]\ : SLE
      port map(D => \r13[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[14]_net_1\);
    
    next_r0_0_cry_1 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[1]\, B => \sum0_5[1]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_0\, S => 
        next_r0_0_cry_1_S, Y => OPEN, FCO => \next_r0_0_cry_1\);
    
    next_r0_0_cry_19 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[19]\, B => \sum0_5[19]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_18\, S
         => next_r0_0_cry_19_S, Y => OPEN, FCO => 
        \next_r0_0_cry_19\);
    
    \r13[12]\ : SLE
      port map(D => \r14[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[12]_net_1\);
    
    \r12[12]\ : SLE
      port map(D => \r13[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[12]_net_1\);
    
    next_r0_0_cry_2 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[2]\, B => \sum0_5[2]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_1\, S => 
        next_r0_0_cry_2_S, Y => OPEN, FCO => \next_r0_0_cry_2\);
    
    sum0_5_cry_22 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[22]_net_1\, B => \r10[22]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_21\, S => 
        \sum0_5[22]\, Y => OPEN, FCO => \sum0_5_cry_22\);
    
    \r3[19]\ : SLE
      port map(D => \r4[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[19]_net_1\);
    
    next_r0_0_cry_29 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[29]\, B => \sum0_5[29]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_28\, S
         => next_r0_0_cry_29_S, Y => OPEN, FCO => 
        \next_r0_0_cry_29\);
    
    \r10[15]\ : SLE
      port map(D => \r11[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[15]_net_1\);
    
    \r2[18]\ : SLE
      port map(D => \r3[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[18]_net_1\);
    
    \r3[25]\ : SLE
      port map(D => \r4[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[25]_net_1\);
    
    \r1[10]\ : SLE
      port map(D => \r2[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[10]_net_1\);
    
    sum0_5_cry_0 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[0]_net_1\, B => \r10[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => GND_net_1, S => OPEN, Y
         => sum0_5_cry_0_Y, FCO => \sum0_5_cry_0\);
    
    \s0[27]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[13]_net_1\, B => \r2[2]_net_1\, C => 
        \r2[30]_net_1\, Y => \s0[27]_net_1\);
    
    \r14[0]\ : SLE
      port map(D => \r15[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[0]_net_1\);
    
    \next_r0[20]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_299, C => next_r0_0_cry_20_S, 
        D => W_out_2_i_1_12, Y => \Wt_data[20]\);
    
    sum0_4_cry_0_1026 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[26]_net_1\, B => \r2[15]_net_1\, C => 
        \r2[11]_net_1\, Y => \s0_0[8]\);
    
    \s0[17]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[24]_net_1\, B => \r2[20]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0[17]_net_1\);
    
    sum0_4_cry_0_1016 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[25]_net_1\, B => \r2[21]_net_1\, C => 
        \r2[4]_net_1\, Y => \s0_0[18]\);
    
    \r13[25]\ : SLE
      port map(D => \r14[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[25]_net_1\);
    
    \r8[0]\ : SLE
      port map(D => \r9[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[0]_net_1\);
    
    \r12[27]\ : SLE
      port map(D => \r13[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[27]_net_1\);
    
    \r10[27]\ : SLE
      port map(D => \r11[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[27]_net_1\);
    
    \r6[12]\ : SLE
      port map(D => \r7[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[12]_net_1\);
    
    \r3[5]\ : SLE
      port map(D => \r4[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[5]_net_1\);
    
    \r0[30]\ : SLE
      port map(D => \Wt_data[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[30]_net_1\);
    
    \r2[22]\ : SLE
      port map(D => \r3[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[22]_net_1\);
    
    \r9[28]\ : SLE
      port map(D => \r10[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[28]_net_1\);
    
    \r11[1]\ : SLE
      port map(D => \r12[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[1]_net_1\);
    
    sum0_5_cry_17 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[17]_net_1\, B => \r10[17]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_16\, S => 
        \sum0_5[17]\, Y => OPEN, FCO => \sum0_5_cry_17\);
    
    next_r0_0_cry_8 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[8]\, B => \sum0_5[8]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_7\, S => 
        next_r0_0_cry_8_S, Y => OPEN, FCO => \next_r0_0_cry_8\);
    
    \r0[27]\ : SLE
      port map(D => \Wt_data[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[27]_net_1\);
    
    next_r0_0_cry_6 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[6]\, B => \sum0_5[6]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_5\, S => 
        next_r0_0_cry_6_S, Y => OPEN, FCO => \next_r0_0_cry_6\);
    
    \r0[17]\ : SLE
      port map(D => \Wt_data[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[17]_net_1\);
    
    \r15[4]\ : SLE
      port map(D => \r0[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[4]_net_1\);
    
    \r14[8]\ : SLE
      port map(D => \r15[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[8]_net_1\);
    
    \r14[28]\ : SLE
      port map(D => \r15[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[28]_net_1\);
    
    \r12[7]\ : SLE
      port map(D => \r13[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[7]_net_1\);
    
    next_r0_0_cry_3 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[3]\, B => \sum0_5[3]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_2\, S => 
        next_r0_0_cry_3_S, Y => OPEN, FCO => \next_r0_0_cry_3\);
    
    \r3[22]\ : SLE
      port map(D => \r4[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[22]_net_1\);
    
    \r8[2]\ : SLE
      port map(D => \r9[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[2]_net_1\);
    
    \s0[28]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[14]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0[28]_net_1\);
    
    \s0[18]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[25]_net_1\, B => \r2[21]_net_1\, C => 
        \r2[4]_net_1\, Y => \s0[18]_net_1\);
    
    \r4[19]\ : SLE
      port map(D => \r5[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[19]_net_1\);
    
    sum0_4_cry_11 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[11]\, C => 
        \sum0_4_axb_11\, D => GND_net_1, FCI => \sum0_4_cry_10\, 
        S => \sum0_4[11]\, Y => OPEN, FCO => \sum0_4_cry_11\);
    
    \r13[16]\ : SLE
      port map(D => \r14[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[16]_net_1\);
    
    \r12[16]\ : SLE
      port map(D => \r13[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[16]_net_1\);
    
    \r5[30]\ : SLE
      port map(D => \r6[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[30]_net_1\);
    
    \r7[7]\ : SLE
      port map(D => \r8[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[7]_net_1\);
    
    sum0_4_axb_3 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[13]_net_1\, B => \s0[3]_net_1\, C => 
        \r15[22]_net_1\, D => \r15[20]_net_1\, Y => 
        \sum0_4_axb_3\);
    
    \r1[25]\ : SLE
      port map(D => \r2[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[25]_net_1\);
    
    \r5[15]\ : SLE
      port map(D => \r6[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[15]_net_1\);
    
    sum0_4_cry_0_1033 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[19]_net_1\, B => \r2[8]_net_1\, C => 
        \r2[4]_net_1\, Y => \s0_0[1]\);
    
    \r8[27]\ : SLE
      port map(D => \r9[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[27]_net_1\);
    
    \r10[17]\ : SLE
      port map(D => \r11[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[17]_net_1\);
    
    next_r0_0_cry_9 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[9]\, B => \sum0_5[9]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_8\, S => 
        next_r0_0_cry_9_S, Y => OPEN, FCO => \next_r0_0_cry_9\);
    
    \r4[25]\ : SLE
      port map(D => \r5[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[25]_net_1\);
    
    \r1[9]\ : SLE
      port map(D => \r2[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[9]_net_1\);
    
    \r8[16]\ : SLE
      port map(D => \r9[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[16]_net_1\);
    
    sum0_4_axb_16 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[1]_net_1\, B => \r15[3]_net_1\, C => 
        \s0[16]_net_1\, D => \r15[26]_net_1\, Y => 
        \sum0_4_axb_16\);
    
    \r10[1]\ : SLE
      port map(D => \r11[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[1]_net_1\);
    
    \s0[29]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \r2[4]_net_1\, B => \r2[15]_net_1\, Y => 
        \s0[29]_net_1\);
    
    \r0[28]\ : SLE
      port map(D => \Wt_data[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[28]_net_1\);
    
    \r9[6]\ : SLE
      port map(D => \r10[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[6]_net_1\);
    
    \s0[19]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[26]_net_1\, B => \r2[22]_net_1\, C => 
        \r2[5]_net_1\, Y => \s0[19]_net_1\);
    
    sum0_4_axb_19 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[4]_net_1\, B => \r15[6]_net_1\, C => 
        \s0[19]_net_1\, D => \r15[29]_net_1\, Y => 
        \sum0_4_axb_19\);
    
    \r0[18]\ : SLE
      port map(D => \Wt_data[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[18]_net_1\);
    
    \r2[15]\ : SLE
      port map(D => \r3[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[15]_net_1\);
    
    \r7[19]\ : SLE
      port map(D => \r8[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[19]_net_1\);
    
    \r13[27]\ : SLE
      port map(D => \r14[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[27]_net_1\);
    
    \r9[8]\ : SLE
      port map(D => \r10[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[8]_net_1\);
    
    \r8[11]\ : SLE
      port map(D => \r9[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[11]_net_1\);
    
    \r14[21]\ : SLE
      port map(D => \r15[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[21]_net_1\);
    
    \r12[23]\ : SLE
      port map(D => \r13[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[23]_net_1\);
    
    \r10[23]\ : SLE
      port map(D => \r11[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[23]_net_1\);
    
    \r9[14]\ : SLE
      port map(D => \r10[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[14]_net_1\);
    
    sum0_5_cry_14 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[14]_net_1\, B => \r10[14]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_13\, S => 
        \sum0_5[14]\, Y => OPEN, FCO => \sum0_5_cry_14\);
    
    \next_r0[10]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_266, C => next_r0_0_cry_10_S, 
        D => W_out_2_i_1_2, Y => \Wt_data[10]\);
    
    sum0_4_cry_0_1032 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[20]_net_1\, B => \r2[9]_net_1\, C => 
        \r2[5]_net_1\, Y => \s0_0[2]\);
    
    sum0_4_axb_8 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[18]_net_1\, B => \s0[8]_net_1\, C => 
        \r15[27]_net_1\, D => \r15[25]_net_1\, Y => 
        \sum0_4_axb_8\);
    
    \r1[22]\ : SLE
      port map(D => \r2[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[22]_net_1\);
    
    \r11[20]\ : SLE
      port map(D => \r12[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[20]_net_1\);
    
    \r5[12]\ : SLE
      port map(D => \r6[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[12]_net_1\);
    
    \r3[14]\ : SLE
      port map(D => \r4[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[14]_net_1\);
    
    \r8[28]\ : SLE
      port map(D => \r9[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[28]_net_1\);
    
    \r5[6]\ : SLE
      port map(D => \r6[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[6]_net_1\);
    
    sum0_4_axb_11 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[21]_net_1\, B => \s0[11]_net_1\, C => 
        \r15[30]_net_1\, D => \r15[28]_net_1\, Y => 
        \sum0_4_axb_11\);
    
    sum0_4_cry_2 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[2]\, C => 
        \sum0_4_axb_2\, D => GND_net_1, FCI => \sum0_4_cry_1\, S
         => \sum0_4[2]\, Y => OPEN, FCO => \sum0_4_cry_2\);
    
    \r11[10]\ : SLE
      port map(D => \r12[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[10]_net_1\);
    
    sum0_4_cry_25 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[25]\, C => 
        \sum0_4_axb_25\, D => GND_net_1, FCI => \sum0_4_cry_24\, 
        S => \sum0_4[25]\, Y => OPEN, FCO => \sum0_4_cry_25\);
    
    \r4[22]\ : SLE
      port map(D => \r5[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[22]_net_1\);
    
    \r9[25]\ : SLE
      port map(D => \r10[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[25]_net_1\);
    
    \next_r0[26]\ : CFG4
      generic map(INIT => x"C0D1")

      port map(A => W_out_2_i_1_18, B => ld_i_i_3, C => 
        next_r0_0_cry_26_S, D => W_out_2_i_0(26), Y => 
        \Wt_data[26]\);
    
    \r12[29]\ : SLE
      port map(D => \r13[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[29]_net_1\);
    
    \r10[29]\ : SLE
      port map(D => \r11[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[29]_net_1\);
    
    \r5[26]\ : SLE
      port map(D => \r6[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[26]_net_1\);
    
    \r1[19]\ : SLE
      port map(D => \r2[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[19]_net_1\);
    
    sum0_4_axb_23 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[8]_net_1\, B => \r15[10]_net_1\, C => 
        \s0[23]_net_1\, Y => \sum0_4_axb_23\);
    
    \r8[5]\ : SLE
      port map(D => \r9[5]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[5]_net_1\);
    
    sum0_4_axb_5 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[15]_net_1\, B => \s0[5]_net_1\, C => 
        \r15[24]_net_1\, D => \r15[22]_net_1\, Y => 
        \sum0_4_axb_5\);
    
    \r8[13]\ : SLE
      port map(D => \r9[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[13]_net_1\);
    
    sum0_4_cry_0_1023 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[29]_net_1\, B => \r2[18]_net_1\, C => 
        \r2[14]_net_1\, Y => \s0_0[11]\);
    
    \r9[31]\ : SLE
      port map(D => \r10[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[31]_net_1\);
    
    \r0[4]\ : SLE
      port map(D => \Wt_data[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[4]_net_1\);
    
    sum0_4_cry_0_1013 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[28]_net_1\, B => \r2[24]_net_1\, C => 
        \r2[7]_net_1\, Y => \s0_0[21]\);
    
    sum0_4_axb_20 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[5]_net_1\, B => \r15[7]_net_1\, C => 
        \s0[20]_net_1\, D => \r15[30]_net_1\, Y => 
        \sum0_4_axb_20\);
    
    \r7[20]\ : SLE
      port map(D => \r8[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[20]_net_1\);
    
    \r2[12]\ : SLE
      port map(D => \r3[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[12]_net_1\);
    
    \r15[0]\ : SLE
      port map(D => \r0[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[0]_net_1\);
    
    \r1[6]\ : SLE
      port map(D => \r2[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[6]_net_1\);
    
    \s0[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[19]_net_1\, B => \r2[8]_net_1\, C => 
        \r2[4]_net_1\, Y => \s0[1]_net_1\);
    
    \r0[5]\ : SLE
      port map(D => \Wt_data[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[5]_net_1\);
    
    \r15[6]\ : SLE
      port map(D => \r0[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[6]_net_1\);
    
    \r6[4]\ : SLE
      port map(D => \r7[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[4]_net_1\);
    
    \r5[21]\ : SLE
      port map(D => \r6[21]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[21]_net_1\);
    
    \r10[13]\ : SLE
      port map(D => \r11[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[13]_net_1\);
    
    \r0[6]\ : SLE
      port map(D => \Wt_data[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[6]_net_1\);
    
    sum0_4_cry_0_1028 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[24]_net_1\, B => \r2[13]_net_1\, C => 
        \r2[9]_net_1\, Y => \s0_0[6]\);
    
    sum0_4_axb_12 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[22]_net_1\, B => \s0[12]_net_1\, C => 
        \r15[31]_net_1\, D => \r15[29]_net_1\, Y => 
        \sum0_4_axb_12\);
    
    \r4[2]\ : SLE
      port map(D => \r5[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[2]_net_1\);
    
    \r12[24]\ : SLE
      port map(D => \r13[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[24]_net_1\);
    
    \r10[24]\ : SLE
      port map(D => \r11[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[24]_net_1\);
    
    sum0_4_cry_0_1018 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[19]_net_1\, B => \r2[2]_net_1\, C => 
        \r2[23]_net_1\, Y => \s0_0[16]\);
    
    sum0_5_cry_27 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[27]_net_1\, B => \r10[27]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_26\, S => 
        \sum0_5[27]\, Y => OPEN, FCO => \sum0_5_cry_27\);
    
    \r6[20]\ : SLE
      port map(D => \r7[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[20]_net_1\);
    
    \r12[22]\ : SLE
      port map(D => \r13[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[22]_net_1\);
    
    \r10[22]\ : SLE
      port map(D => \r11[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[22]_net_1\);
    
    \r8[30]\ : SLE
      port map(D => \r9[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[30]_net_1\);
    
    \r3[6]\ : SLE
      port map(D => \r4[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[6]_net_1\);
    
    sum0_4_axb_15 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[0]_net_1\, B => \r15[2]_net_1\, C => 
        \s0[15]_net_1\, D => \r15[25]_net_1\, Y => 
        \sum0_4_axb_15\);
    
    sum0_4_axb_9 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[19]_net_1\, B => \s0[9]_net_1\, C => 
        \r15[28]_net_1\, D => \r15[26]_net_1\, Y => 
        \sum0_4_axb_9\);
    
    \r9[22]\ : SLE
      port map(D => \r10[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[22]_net_1\);
    
    \r13[23]\ : SLE
      port map(D => \r14[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[23]_net_1\);
    
    \r10[19]\ : SLE
      port map(D => \r11[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[19]_net_1\);
    
    sum0_4_cry_0_1022 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[30]_net_1\, B => \r2[19]_net_1\, C => 
        \r2[15]_net_1\, Y => \s0_0[12]\);
    
    \r0[25]\ : SLE
      port map(D => \Wt_data[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[25]_net_1\);
    
    sum0_4_cry_5 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[5]\, C => 
        \sum0_4_axb_5\, D => GND_net_1, FCI => \sum0_4_cry_4\, S
         => \sum0_4[5]\, Y => OPEN, FCO => \sum0_4_cry_5\);
    
    \r4[14]\ : SLE
      port map(D => \r5[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[14]_net_1\);
    
    sum0_4_cry_0_1012 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[29]_net_1\, B => \r2[25]_net_1\, C => 
        \r2[8]_net_1\, Y => \s0_0[22]\);
    
    \r0[15]\ : SLE
      port map(D => \Wt_data[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[15]_net_1\);
    
    \r5[23]\ : SLE
      port map(D => \r6[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[23]_net_1\);
    
    \r13[9]\ : SLE
      port map(D => \r14[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[9]_net_1\);
    
    \r11[25]\ : SLE
      port map(D => \r12[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[25]_net_1\);
    
    sum0_4_cry_10 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[10]\, C => 
        \sum0_4_axb_10\, D => GND_net_1, FCI => \sum0_4_cry_9\, S
         => \sum0_4[10]\, Y => OPEN, FCO => \sum0_4_cry_10\);
    
    sum0_4_cry_0_1034 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[18]_net_1\, B => \r2[7]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0_0[0]\);
    
    next_r0_0_cry_7 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[7]\, B => \sum0_5[7]\, C => GND_net_1, 
        D => GND_net_1, FCI => \next_r0_0_cry_6\, S => 
        next_r0_0_cry_7_S, Y => OPEN, FCO => \next_r0_0_cry_7\);
    
    \r11[15]\ : SLE
      port map(D => \r12[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[15]_net_1\);
    
    \r13[29]\ : SLE
      port map(D => \r14[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[29]_net_1\);
    
    sum0_5_cry_3 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[3]_net_1\, B => \r10[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_2\, S => 
        \sum0_5[3]\, Y => OPEN, FCO => \sum0_5_cry_3\);
    
    \r0[8]\ : SLE
      port map(D => \Wt_data[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[8]_net_1\);
    
    next_r0_0_cry_10 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[10]\, B => \sum0_5[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_9\, S
         => next_r0_0_cry_10_S, Y => OPEN, FCO => 
        \next_r0_0_cry_10\);
    
    \r13[7]\ : SLE
      port map(D => \r14[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[7]_net_1\);
    
    \r14[2]\ : SLE
      port map(D => \r15[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[2]_net_1\);
    
    \next_r0[21]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_302, C => next_r0_0_cry_21_S, 
        D => W_out_2_i_1_13, Y => \Wt_data[21]\);
    
    \r10[14]\ : SLE
      port map(D => \r11[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[14]_net_1\);
    
    next_r0_0_cry_20 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[20]\, B => \sum0_5[20]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_19\, S
         => next_r0_0_cry_20_S, Y => OPEN, FCO => 
        \next_r0_0_cry_20\);
    
    \r15[10]\ : SLE
      port map(D => \r0[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[10]_net_1\);
    
    \r10[12]\ : SLE
      port map(D => \r11[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[12]_net_1\);
    
    \r8[25]\ : SLE
      port map(D => \r9[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[25]_net_1\);
    
    \r6[10]\ : SLE
      port map(D => \r7[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[10]_net_1\);
    
    \r7[14]\ : SLE
      port map(D => \r8[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[14]_net_1\);
    
    sum0_4_axb_0 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[10]_net_1\, B => \s0[0]_net_1\, C => 
        \r15[19]_net_1\, D => \r15[17]_net_1\, Y => \sum0_4[0]\);
    
    \r15[20]\ : SLE
      port map(D => \r0[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[20]_net_1\);
    
    \r2[20]\ : SLE
      port map(D => \r3[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[20]_net_1\);
    
    \next_r0[16]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_287, C => next_r0_0_cry_16_S, 
        D => W_out_2_i_1_8, Y => \Wt_data[16]\);
    
    sum0_4_cry_13 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[13]\, C => 
        \sum0_4_axb_13\, D => GND_net_1, FCI => \sum0_4_cry_12\, 
        S => \sum0_4[13]\, Y => OPEN, FCO => \sum0_4_cry_13\);
    
    sum0_4_axb_4 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[14]_net_1\, B => \s0[4]_net_1\, C => 
        \r15[23]_net_1\, D => \r15[21]_net_1\, Y => 
        \sum0_4_axb_4\);
    
    \r0[22]\ : SLE
      port map(D => \Wt_data[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[22]_net_1\);
    
    \r13[24]\ : SLE
      port map(D => \r14[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[24]_net_1\);
    
    \r12[26]\ : SLE
      port map(D => \r13[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[26]_net_1\);
    
    \r10[26]\ : SLE
      port map(D => \r11[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[26]_net_1\);
    
    \r2[31]\ : SLE
      port map(D => \r3[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[31]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \r0[12]\ : SLE
      port map(D => \Wt_data[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[12]_net_1\);
    
    sum0_5_cry_24 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[24]_net_1\, B => \r10[24]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_23\, S => 
        \sum0_5[24]\, Y => OPEN, FCO => \sum0_5_cry_24\);
    
    \r13[22]\ : SLE
      port map(D => \r14[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[22]_net_1\);
    
    \r8[17]\ : SLE
      port map(D => \r9[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[17]_net_1\);
    
    \r11[31]\ : SLE
      port map(D => \r12[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[31]_net_1\);
    
    \r0[0]\ : SLE
      port map(D => \Wt_data[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[0]_net_1\);
    
    \r5[2]\ : SLE
      port map(D => \r6[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[2]_net_1\);
    
    \r13[31]\ : SLE
      port map(D => \r14[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[31]_net_1\);
    
    sum0_4_cry_18 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[18]\, C => 
        \sum0_4_axb_18\, D => GND_net_1, FCI => \sum0_4_cry_17\, 
        S => \sum0_4[18]\, Y => OPEN, FCO => \sum0_4_cry_18\);
    
    \r3[20]\ : SLE
      port map(D => \r4[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[20]_net_1\);
    
    \r12[3]\ : SLE
      port map(D => \r13[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[3]_net_1\);
    
    sum0_4_axb_2 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[12]_net_1\, B => \s0[2]_net_1\, C => 
        \r15[21]_net_1\, D => \r15[19]_net_1\, Y => 
        \sum0_4_axb_2\);
    
    sum0_4_axb_7 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[17]_net_1\, B => \s0[7]_net_1\, C => 
        \r15[26]_net_1\, D => \r15[24]_net_1\, Y => 
        \sum0_4_axb_7\);
    
    \r13[18]\ : SLE
      port map(D => \r14[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[18]_net_1\);
    
    \r12[18]\ : SLE
      port map(D => \r13[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[18]_net_1\);
    
    \r1[14]\ : SLE
      port map(D => \r2[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[14]_net_1\);
    
    sum0_4_cry_0_1024 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[28]_net_1\, B => \r2[13]_net_1\, C => 
        \r2[17]_net_1\, Y => \s0_0[10]\);
    
    \r8[22]\ : SLE
      port map(D => \r9[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[22]_net_1\);
    
    \r5[4]\ : SLE
      port map(D => \r6[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[4]_net_1\);
    
    sum0_4_cry_0_1014 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[23]_net_1\, B => \r2[6]_net_1\, C => 
        \r2[27]_net_1\, Y => \s0_0[20]\);
    
    \r3[2]\ : SLE
      port map(D => \r4[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[2]_net_1\);
    
    sum0_5_cry_1 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[1]_net_1\, B => \r10[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_0\, S => 
        \sum0_5[1]\, Y => OPEN, FCO => \sum0_5_cry_1\);
    
    sum0_5_cry_15 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[15]_net_1\, B => \r10[15]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_14\, S => 
        \sum0_5[15]\, Y => OPEN, FCO => \sum0_5_cry_15\);
    
    \s0[30]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \r2[5]_net_1\, B => \r2[16]_net_1\, Y => 
        \s0[30]_net_1\);
    
    next_r0_0_cry_30 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[30]\, B => \sum0_5[30]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_29\, S
         => next_r0_0_cry_30_S, Y => OPEN, FCO => 
        \next_r0_0_cry_30\);
    
    \r9[1]\ : SLE
      port map(D => \r10[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[1]_net_1\);
    
    \r7[6]\ : SLE
      port map(D => \r8[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[6]_net_1\);
    
    sum0_4_axb_24 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[9]_net_1\, B => \r15[11]_net_1\, C => 
        \s0[24]_net_1\, Y => \sum0_4_axb_24\);
    
    \r11[27]\ : SLE
      port map(D => \r12[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[27]_net_1\);
    
    \r7[29]\ : SLE
      port map(D => \r8[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[29]_net_1\);
    
    \r1[7]\ : SLE
      port map(D => \r2[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[7]_net_1\);
    
    \r11[17]\ : SLE
      port map(D => \r12[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[17]_net_1\);
    
    \r7[8]\ : SLE
      port map(D => \r8[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[8]_net_1\);
    
    \next_r0[4]\ : CFG4
      generic map(INIT => x"AFAC")

      port map(A => next_r0_0_cry_4_S, B => N_248, C => ld_i_i_3, 
        D => W_out_2_0_0_1, Y => \Wt_data[4]\);
    
    \r6[8]\ : SLE
      port map(D => \r7[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[8]_net_1\);
    
    \r13[0]\ : SLE
      port map(D => \r14[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[0]_net_1\);
    
    \r12[4]\ : SLE
      port map(D => \r13[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[4]_net_1\);
    
    \r10[0]\ : SLE
      port map(D => \r11[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[0]_net_1\);
    
    \r9[16]\ : SLE
      port map(D => \r10[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[16]_net_1\);
    
    \r10[16]\ : SLE
      port map(D => \r11[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[16]_net_1\);
    
    \r8[8]\ : SLE
      port map(D => \r9[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[8]_net_1\);
    
    \r8[18]\ : SLE
      port map(D => \r9[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[18]_net_1\);
    
    \r15[15]\ : SLE
      port map(D => \r0[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[15]_net_1\);
    
    \r14[30]\ : SLE
      port map(D => \r15[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[30]_net_1\);
    
    \r14[10]\ : SLE
      port map(D => \r15[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[10]_net_1\);
    
    \r3[30]\ : SLE
      port map(D => \r4[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[30]_net_1\);
    
    sum0_4_axb_27 : CFG3
      generic map(INIT => x"96")

      port map(A => \r15[12]_net_1\, B => \s0[27]_net_1\, C => 
        \r15[14]_net_1\, Y => \sum0_4_axb_27\);
    
    \r5[27]\ : SLE
      port map(D => \r6[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[27]_net_1\);
    
    \r3[16]\ : SLE
      port map(D => \r4[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[16]_net_1\);
    
    \r6[29]\ : SLE
      port map(D => \r7[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[29]_net_1\);
    
    \r15[25]\ : SLE
      port map(D => \r0[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[25]_net_1\);
    
    \next_r0[2]\ : CFG4
      generic map(INIT => x"C0E2")

      port map(A => N_98, B => ld_i_i_3, C => next_r0_0_cry_2_S, 
        D => W_out_i_0(2), Y => \Wt_data[2]\);
    
    \r3[8]\ : SLE
      port map(D => \r4[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[8]_net_1\);
    
    \r13[26]\ : SLE
      port map(D => \r14[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[26]_net_1\);
    
    \r9[11]\ : SLE
      port map(D => \r10[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[11]_net_1\);
    
    \next_r0[11]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_268, C => next_r0_0_cry_11_S, 
        D => W_out_2_i_1_3, Y => \Wt_data[11]\);
    
    sum0_4_cry_0_1029 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[23]_net_1\, B => \r2[12]_net_1\, C => 
        \r2[8]_net_1\, Y => \s0_0[5]\);
    
    sum0_4_cry_0_1005 : CFG2
      generic map(INIT => x"6")

      port map(A => \r2[4]_net_1\, B => \r2[15]_net_1\, Y => 
        \s0_0[29]\);
    
    sum0_4_cry_30 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[30]\, C => 
        \sum0_4_axb_30\, D => GND_net_1, FCI => \sum0_4_cry_29\, 
        S => \sum0_4[30]\, Y => OPEN, FCO => \sum0_4_cry_30\);
    
    \r1[20]\ : SLE
      port map(D => \r2[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[20]_net_1\);
    
    \r13[11]\ : SLE
      port map(D => \r14[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[11]_net_1\);
    
    \r12[11]\ : SLE
      port map(D => \r13[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[11]_net_1\);
    
    \r10[7]\ : SLE
      port map(D => \r11[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[7]_net_1\);
    
    \r5[10]\ : SLE
      port map(D => \r6[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[10]_net_1\);
    
    sum0_4_cry_0_1019 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[18]_net_1\, B => \r2[1]_net_1\, C => 
        \r2[22]_net_1\, Y => \s0_0[15]\);
    
    \r9[9]\ : SLE
      port map(D => \r10[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[9]_net_1\);
    
    \r4[20]\ : SLE
      port map(D => \r5[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[20]_net_1\);
    
    \r3[11]\ : SLE
      port map(D => \r4[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[11]_net_1\);
    
    sum0_4_axb_13 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[0]_net_1\, B => \r15[30]_net_1\, C => 
        \r15[23]_net_1\, D => \s0[13]_net_1\, Y => 
        \sum0_4_axb_13\);
    
    sum0_4_cry_19 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[19]\, C => 
        \sum0_4_axb_19\, D => GND_net_1, FCI => \sum0_4_cry_18\, 
        S => \sum0_4[19]\, Y => OPEN, FCO => \sum0_4_cry_19\);
    
    \r10[4]\ : SLE
      port map(D => \r11[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[4]_net_1\);
    
    sum0_4_axb_10 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[20]_net_1\, B => \s0[10]_net_1\, C => 
        \r15[29]_net_1\, D => \r15[27]_net_1\, Y => 
        \sum0_4_axb_10\);
    
    \r5[9]\ : SLE
      port map(D => \r6[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[9]_net_1\);
    
    \r2[7]\ : SLE
      port map(D => \r3[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[7]_net_1\);
    
    \r2[10]\ : SLE
      port map(D => \r3[10]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[10]_net_1\);
    
    \r10[30]\ : SLE
      port map(D => \r11[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[30]_net_1\);
    
    sum0_5_cry_5 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[5]_net_1\, B => \r10[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_4\, S => 
        \sum0_5[5]\, Y => OPEN, FCO => \sum0_5_cry_5\);
    
    sum0_4_cry_16 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[16]\, C => 
        \sum0_4_axb_16\, D => GND_net_1, FCI => \sum0_4_cry_15\, 
        S => \sum0_4[16]\, Y => OPEN, FCO => \sum0_4_cry_16\);
    
    \r9[13]\ : SLE
      port map(D => \r10[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[13]_net_1\);
    
    \r3[4]\ : SLE
      port map(D => \r4[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[4]_net_1\);
    
    \r5[28]\ : SLE
      port map(D => \r6[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[28]_net_1\);
    
    \r6[31]\ : SLE
      port map(D => \r7[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[31]_net_1\);
    
    \r6[19]\ : SLE
      port map(D => \r7[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[19]_net_1\);
    
    \r12[30]\ : SLE
      port map(D => \r13[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[30]_net_1\);
    
    \r3[13]\ : SLE
      port map(D => \r4[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[13]_net_1\);
    
    \next_r0[9]\ : CFG4
      generic map(INIT => x"A0B1")

      port map(A => ld_i_i_3, B => N_263, C => next_r0_0_cry_9_S, 
        D => W_out_2_i_1_1, Y => \Wt_data[9]\);
    
    \r2[29]\ : SLE
      port map(D => \r3[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[29]_net_1\);
    
    \r11[23]\ : SLE
      port map(D => \r12[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[23]_net_1\);
    
    \r10[3]\ : SLE
      port map(D => \r11[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[3]_net_1\);
    
    \r4[16]\ : SLE
      port map(D => \r5[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[16]_net_1\);
    
    \r4[8]\ : SLE
      port map(D => \r5[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[8]_net_1\);
    
    \r11[13]\ : SLE
      port map(D => \r12[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[13]_net_1\);
    
    next_r0_0_cry_16 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[16]\, B => \sum0_5[16]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_15\, S
         => next_r0_0_cry_16_S, Y => OPEN, FCO => 
        \next_r0_0_cry_16\);
    
    \r4[30]\ : SLE
      port map(D => \r5[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[30]_net_1\);
    
    \r14[6]\ : SLE
      port map(D => \r15[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[6]_net_1\);
    
    \r14[15]\ : SLE
      port map(D => \r15[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[15]_net_1\);
    
    next_r0_0_cry_26 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[26]\, B => \sum0_5[26]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_25\, S
         => next_r0_0_cry_26_S, Y => OPEN, FCO => 
        \next_r0_0_cry_26\);
    
    \r15[17]\ : SLE
      port map(D => \r0[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[17]_net_1\);
    
    \r9[20]\ : SLE
      port map(D => \r10[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[20]_net_1\);
    
    \r15[27]\ : SLE
      port map(D => \r0[27]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[27]_net_1\);
    
    \r3[29]\ : SLE
      port map(D => \r4[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[29]_net_1\);
    
    \r7[2]\ : SLE
      port map(D => \r8[2]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[2]_net_1\);
    
    \r3[0]\ : SLE
      port map(D => \r4[0]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[0]_net_1\);
    
    \r11[29]\ : SLE
      port map(D => \r12[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[29]_net_1\);
    
    sum0_4_cry_21 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[21]\, C => 
        \sum0_4_axb_21\, D => GND_net_1, FCI => \sum0_4_cry_20\, 
        S => \sum0_4[21]\, Y => OPEN, FCO => \sum0_4_cry_21\);
    
    sum0_4_cry_12 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[12]\, C => 
        \sum0_4_axb_12\, D => GND_net_1, FCI => \sum0_4_cry_11\, 
        S => \sum0_4[12]\, Y => OPEN, FCO => \sum0_4_cry_12\);
    
    \r4[11]\ : SLE
      port map(D => \r5[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[11]_net_1\);
    
    \r1[8]\ : SLE
      port map(D => \r2[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[8]_net_1\);
    
    \r11[19]\ : SLE
      port map(D => \r12[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[19]_net_1\);
    
    \r0[9]\ : SLE
      port map(D => \Wt_data[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[9]_net_1\);
    
    \next_r0[25]\ : CFG4
      generic map(INIT => x"C0D1")

      port map(A => W_out_2_i_1_17, B => ld_i_i_3, C => 
        next_r0_0_cry_25_S, D => W_out_2_i_0(25), Y => 
        \Wt_data[25]\);
    
    \r5[1]\ : SLE
      port map(D => \r6[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[1]_net_1\);
    
    next_r0_0_cry_12 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[12]\, B => \sum0_5[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_11\, S
         => next_r0_0_cry_12_S, Y => OPEN, FCO => 
        \next_r0_0_cry_12\);
    
    sum0_4_cry_9 : ARI1
      generic map(INIT => x"5CCAA")

      port map(A => VCC_net_1, B => \s0_0[9]\, C => 
        \sum0_4_axb_9\, D => GND_net_1, FCI => \sum0_4_cry_8\, S
         => \sum0_4[9]\, Y => OPEN, FCO => \sum0_4_cry_9\);
    
    \r8[15]\ : SLE
      port map(D => \r9[15]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[15]_net_1\);
    
    next_r0_0_cry_22 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[22]\, B => \sum0_5[22]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_21\, S
         => next_r0_0_cry_22_S, Y => OPEN, FCO => 
        \next_r0_0_cry_22\);
    
    sum0_5_cry_2 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[2]_net_1\, B => \r10[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_1\, S => 
        \sum0_5[2]\, Y => OPEN, FCO => \sum0_5_cry_2\);
    
    sum0_5_cry_25 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[25]_net_1\, B => \r10[25]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_24\, S => 
        \sum0_5[25]\, Y => OPEN, FCO => \sum0_5_cry_25\);
    
    \r7[16]\ : SLE
      port map(D => \r8[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[16]_net_1\);
    
    \r8[7]\ : SLE
      port map(D => \r9[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[7]_net_1\);
    
    sum0_4_cry_0_1027 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[25]_net_1\, B => \r2[14]_net_1\, C => 
        \r2[10]_net_1\, Y => \s0_0[7]\);
    
    sum0_5_cry_9 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[9]_net_1\, B => \r10[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_8\, S => 
        \sum0_5[9]\, Y => OPEN, FCO => \sum0_5_cry_9\);
    
    sum0_5_cry_8 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \r1[8]_net_1\, B => \r10[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \sum0_5_cry_7\, S => 
        \sum0_5[8]\, Y => OPEN, FCO => \sum0_5_cry_8\);
    
    \r7[24]\ : SLE
      port map(D => \r8[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[24]_net_1\);
    
    \r1[3]\ : SLE
      port map(D => \r2[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[3]_net_1\);
    
    sum0_4_cry_0_1017 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[24]_net_1\, B => \r2[20]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0_0[17]\);
    
    \s0[2]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[20]_net_1\, B => \r2[9]_net_1\, C => 
        \r2[5]_net_1\, Y => \s0[2]_net_1\);
    
    \s0[24]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[27]_net_1\, C => 
        \r2[10]_net_1\, Y => \s0[24]_net_1\);
    
    next_r0_0_cry_17 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[17]\, B => \sum0_5[17]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_16\, S
         => next_r0_0_cry_17_S, Y => OPEN, FCO => 
        \next_r0_0_cry_17\);
    
    \s0[14]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[0]_net_1\, B => \r2[17]_net_1\, C => 
        \r2[21]_net_1\, Y => \s0[14]_net_1\);
    
    \r7[1]\ : SLE
      port map(D => \r8[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[1]_net_1\);
    
    next_r0_0_cry_27 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[27]\, B => \sum0_5[27]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_26\, S
         => next_r0_0_cry_27_S, Y => OPEN, FCO => 
        \next_r0_0_cry_27\);
    
    \next_r0[24]\ : CFG4
      generic map(INIT => x"C0D1")

      port map(A => W_out_2_i_1_16, B => ld_i_i_3, C => 
        next_r0_0_cry_24_S, D => W_out_2_i_0(24), Y => 
        \Wt_data[24]\);
    
    \r1[31]\ : SLE
      port map(D => \r2[31]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[31]_net_1\);
    
    \r11[24]\ : SLE
      port map(D => \r12[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[24]_net_1\);
    
    \next_r0[27]\ : CFG4
      generic map(INIT => x"C0D1")

      port map(A => W_out_2_i_1_19, B => ld_i_i_3, C => 
        next_r0_0_cry_27_S, D => W_out_2_i_0(27), Y => 
        \Wt_data[27]\);
    
    next_r0_0_cry_15 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[15]\, B => \sum0_5[15]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_14\, S
         => next_r0_0_cry_15_S, Y => OPEN, FCO => 
        \next_r0_0_cry_15\);
    
    \r13[8]\ : SLE
      port map(D => \r14[8]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r13[8]_net_1\);
    
    \r11[22]\ : SLE
      port map(D => \r12[22]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[22]_net_1\);
    
    \r11[14]\ : SLE
      port map(D => \r12[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[14]_net_1\);
    
    \r4[13]\ : SLE
      port map(D => \r5[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[13]_net_1\);
    
    next_r0_0_cry_25 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \sum0_4[25]\, B => \sum0_5[25]\, C => 
        GND_net_1, D => GND_net_1, FCI => \next_r0_0_cry_24\, S
         => next_r0_0_cry_25_S, Y => OPEN, FCO => 
        \next_r0_0_cry_25\);
    
    \r7[11]\ : SLE
      port map(D => \r8[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[11]_net_1\);
    
    \r11[12]\ : SLE
      port map(D => \r12[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[12]_net_1\);
    
    \r5[3]\ : SLE
      port map(D => \r6[3]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[3]_net_1\);
    
    \r6[24]\ : SLE
      port map(D => \r7[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[24]_net_1\);
    
    \s0[22]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[29]_net_1\, B => \r2[25]_net_1\, C => 
        \r2[8]_net_1\, Y => \s0[22]_net_1\);
    
    \next_r0[0]\ : CFG4
      generic map(INIT => x"A3A0")

      port map(A => \next_r0_0_cry_0_Y\, B => W_out_i_1(0), C => 
        ld_i_i_3, D => N_98, Y => \Wt_data[0]\);
    
    \r0[20]\ : SLE
      port map(D => \Wt_data[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[20]_net_1\);
    
    sum0_4_cry_0_1006 : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[31]_net_1\, B => \r2[14]_net_1\, C => 
        \r2[3]_net_1\, Y => \s0_0[28]\);
    
    \r4[4]\ : SLE
      port map(D => \r5[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[4]_net_1\);
    
    \s0[12]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \r2[30]_net_1\, B => \r2[19]_net_1\, C => 
        \r2[15]_net_1\, Y => \s0[12]_net_1\);
    
    \r15[1]\ : SLE
      port map(D => \r0[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[1]_net_1\);
    
    \r8[1]\ : SLE
      port map(D => \r9[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[1]_net_1\);
    
    \r12[28]\ : SLE
      port map(D => \r13[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[28]_net_1\);
    
    \r10[28]\ : SLE
      port map(D => \r11[28]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[28]_net_1\);
    
    \r0[10]\ : SLE
      port map(D => \Wt_data[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[10]_net_1\);
    
    \r1[16]\ : SLE
      port map(D => \r2[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[16]_net_1\);
    
    \next_r0[28]\ : CFG4
      generic map(INIT => x"C0D1")

      port map(A => W_out_2_i_1_20, B => ld_i_i_3, C => 
        next_r0_0_cry_28_S, D => W_out_2_i_0(28), Y => 
        \Wt_data[28]\);
    
    \r8[12]\ : SLE
      port map(D => \r9[12]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[12]_net_1\);
    
    \r12[1]\ : SLE
      port map(D => \r13[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r12[1]_net_1\);
    
    \r5[25]\ : SLE
      port map(D => \r6[25]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[25]_net_1\);
    
    sum0_4_axb_1 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[11]_net_1\, B => \s0[1]_net_1\, C => 
        \r15[20]_net_1\, D => \r15[18]_net_1\, Y => 
        \sum0_4_axb_1\);
    
    \r14[17]\ : SLE
      port map(D => \r15[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[17]_net_1\);
    
    \r1[29]\ : SLE
      port map(D => \r2[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[29]_net_1\);
    
    \r9[17]\ : SLE
      port map(D => \r10[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r9[17]_net_1\);
    
    \r5[19]\ : SLE
      port map(D => \r6[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r5[19]_net_1\);
    
    \r11[7]\ : SLE
      port map(D => \r12[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[7]_net_1\);
    
    \r4[29]\ : SLE
      port map(D => \r5[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[29]_net_1\);
    
    \r4[6]\ : SLE
      port map(D => \r5[6]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[6]_net_1\);
    
    \r15[13]\ : SLE
      port map(D => \r0[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[13]_net_1\);
    
    \r11[4]\ : SLE
      port map(D => \r12[4]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[4]_net_1\);
    
    \r7[13]\ : SLE
      port map(D => \r8[13]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[13]_net_1\);
    
    \r3[17]\ : SLE
      port map(D => \r4[17]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r3[17]_net_1\);
    
    \r1[11]\ : SLE
      port map(D => \r2[11]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r1[11]_net_1\);
    
    \r15[23]\ : SLE
      port map(D => \r0[23]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[23]_net_1\);
    
    sum0_4_axb_14 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[1]_net_1\, B => \r15[31]_net_1\, C => 
        \r15[24]_net_1\, D => \s0[14]_net_1\, Y => 
        \sum0_4_axb_14\);
    
    \r4[1]\ : SLE
      port map(D => \r5[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r4[1]_net_1\);
    
    \r8[20]\ : SLE
      port map(D => \r9[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r8[20]_net_1\);
    
    \r15[7]\ : SLE
      port map(D => \r0[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[7]_net_1\);
    
    \r2[9]\ : SLE
      port map(D => \r3[9]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[9]_net_1\);
    
    next_r0_0_s_31 : ARI1
      generic map(INIT => x"46600")

      port map(A => VCC_net_1, B => \sum0_4[31]\, C => 
        \sum0_5[31]\, D => GND_net_1, FCI => \next_r0_0_cry_30\, 
        S => next_r0_0_s_31_S, Y => OPEN, FCO => OPEN);
    
    \r2[19]\ : SLE
      port map(D => \r3[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[19]_net_1\);
    
    \r14[20]\ : SLE
      port map(D => \r15[20]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[20]_net_1\);
    
    \r15[19]\ : SLE
      port map(D => \r0[19]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[19]_net_1\);
    
    \r14[7]\ : SLE
      port map(D => \r15[7]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r14[7]_net_1\);
    
    \r6[14]\ : SLE
      port map(D => \r7[14]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[14]_net_1\);
    
    \r6[1]\ : SLE
      port map(D => \r7[1]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r6[1]_net_1\);
    
    \r10[18]\ : SLE
      port map(D => \r11[18]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r10[18]_net_1\);
    
    \r15[29]\ : SLE
      port map(D => \r0[29]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r15[29]_net_1\);
    
    sum0_4_axb_17 : CFG4
      generic map(INIT => x"6996")

      port map(A => \r15[2]_net_1\, B => \r15[4]_net_1\, C => 
        \s0[17]_net_1\, D => \r15[27]_net_1\, Y => 
        \sum0_4_axb_17\);
    
    \next_r0[15]\ : CFG4
      generic map(INIT => x"F5E4")

      port map(A => ld_i_i_3, B => W_out_2_0_2_0, C => 
        next_r0_0_cry_15_S, D => W_out_2_0_1_8, Y => 
        \Wt_data[15]\);
    
    \r2[24]\ : SLE
      port map(D => \r3[24]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r2[24]_net_1\);
    
    \r11[26]\ : SLE
      port map(D => \r12[26]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[26]_net_1\);
    
    \r0[31]\ : SLE
      port map(D => \Wt_data[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r0[31]_net_1\);
    
    \r7[30]\ : SLE
      port map(D => \r8[30]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r7[30]_net_1\);
    
    \next_r0[7]\ : CFG4
      generic map(INIT => x"AFAC")

      port map(A => next_r0_0_cry_7_S, B => N_255, C => ld_i_i_3, 
        D => W_out_2_0_1_0, Y => \Wt_data[7]\);
    
    \r11[16]\ : SLE
      port map(D => \r12[16]_net_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_244_i_0, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \r11[16]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sha256_kt_rom is

    port( hash_control_st_reg_ns_i_0_a2_0 : in    std_logic_vector(4 to 4);
          Kt_addr_fast                    : in    std_logic_vector(4 downto 0);
          hash_control_st_reg_ns_i_0_a2_2 : out   std_logic_vector(4 to 4);
          Kt_addr                         : in    std_logic_vector(5 downto 0);
          Kt_data_9                       : out   std_logic;
          Kt_data_0                       : out   std_logic;
          Kt_addr_3_rep1                  : in    std_logic;
          m62_am                          : out   std_logic;
          Kt_addr_0_rep1                  : in    std_logic;
          m104_bm                         : out   std_logic;
          Kt_addr_2_rep1                  : in    std_logic;
          Kt_addr_0_rep2                  : in    std_logic;
          m49_am                          : out   std_logic;
          Kt_addr_1_rep1                  : in    std_logic;
          m49_bm                          : out   std_logic;
          m137_am                         : out   std_logic;
          Kt_addr_3_rep2                  : in    std_logic;
          m137_bm                         : out   std_logic;
          Kt_addr_4_rep2                  : in    std_logic;
          m215_am                         : out   std_logic;
          Kt_addr_4_rep1                  : in    std_logic;
          m215_bm                         : out   std_logic;
          Kt_addr_2_rep2                  : in    std_logic;
          m250_am                         : out   std_logic;
          Kt_addr_1_rep2                  : in    std_logic;
          m250_bm                         : out   std_logic;
          m207_1_1                        : out   std_logic;
          m207_1_0                        : out   std_logic;
          m157                            : out   std_logic;
          m197_1_1                        : out   std_logic;
          m197_1_0                        : out   std_logic;
          m95_1_1                         : out   std_logic;
          m95_1_0                         : out   std_logic;
          m325                            : out   std_logic;
          m168_1_1                        : out   std_logic;
          m168_1_0                        : out   std_logic;
          m316                            : out   std_logic;
          m34                             : out   std_logic;
          m114                            : out   std_logic;
          m285                            : out   std_logic;
          m289                            : out   std_logic;
          m254                            : out   std_logic;
          m239                            : out   std_logic;
          m124                            : out   std_logic;
          m141                            : out   std_logic;
          m304                            : out   std_logic;
          m19                             : out   std_logic;
          pad_one_reg_0_0_a2_0            : in    std_logic;
          m296                            : out   std_logic;
          m78                             : out   std_logic;
          m219                            : out   std_logic;
          m230                            : out   std_logic;
          m177                            : out   std_logic;
          m73_0                           : out   std_logic;
          i3_mux_1                        : out   std_logic;
          m10_ns                          : out   std_logic;
          m67_ns                          : out   std_logic;
          m83_ns                          : out   std_logic;
          m110_ns                         : out   std_logic;
          m119_ns                         : out   std_logic;
          m144_ns                         : out   std_logic;
          m172_ns                         : out   std_logic;
          m222_ns                         : out   std_logic;
          m226_ns                         : out   std_logic;
          m235_ns                         : out   std_logic;
          m258_ns                         : out   std_logic;
          m276_ns                         : out   std_logic;
          m281_ns                         : out   std_logic;
          m292_ns                         : out   std_logic;
          m300_ns                         : out   std_logic;
          sha_last_blk_next_0_a4_0        : out   std_logic;
          m273                            : out   std_logic;
          m104_am                         : out   std_logic;
          m62_bm                          : out   std_logic
        );

end sha256_kt_rom;

architecture DEF_ARCH of sha256_kt_rom is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal m62_am_1_0, m62_am_1, m54, m53, m51, m304_2, 
        m104_bm_1, m103_1, m79, m78_1, m49_am_1_0, m35, m48_2, 
        m49_bm_1, m48_1, m43, m137_am_1_0, m129, m126, m127, 
        m137_bm_1_0, m137_bm_1, m17, m133, m132, m215_am_1_0, 
        m211_0, m209, m92, m215_bm_1_0, m215_bm_1, m90, m22, m164, 
        m273_2, m250_am_1, m194, m85, m250_bm_1_0_1, m250_bm_1_0, 
        m205, m202, m207_1_0_1, m155, m157_1_2, m153, m151, m148, 
        m195, m193, m185, m191, m93, m91, m46, m87, m270_2, 
        m270_1_1, m266, m263, m261, 
        \hash_control_st_reg_ns_i_0_a2_2[4]\, m325_1_1, m325_1_0, 
        m323, m318, m325_1_0_1, m166, m163, m168_1_0_1, m316_2, 
        m316_1_1, m313, m311, m310, m186, m188_1_2, m184, m181, 
        m180, m32, m34_1_2, m30, i2_mux, m23, m230_0, m296_2, 
        m114_1_0, m63, m285_1_1_1, m285_1_1, m28, m289_1_1, 
        m289_1_0, m37, m1, m237, m254_1_1, m254_1_0, m252, m232, 
        m105, m239_1_2, m81, m227, m124_1_2, m16, m120, m122, 
        m141_1, m177_1, m138, m304_1_0, m304_1, m216, m19_1_1, 
        m19_1_0, m13, m296_1_1, m78_2, m78_1_0, m219_1_2, m68, 
        m230_1_1, m177_2, m177_1_0, m174, m73_1, m73_1_0, m73, 
        m71, m117, m308_ns_1, m10_bm, m10_am, m67_bm, m67_am, 
        m83_bm, m83_am, m110_bm, m110_am, m119_bm, m119_am, 
        m144_bm, m144_am, m172_bm, m172_am, m222_bm, m222_am, 
        m226_bm, m226_am, m235_bm, m235_am, m258_bm, m258_am, 
        m276_bm, m276_am, m281_bm, m281_am, m292_bm, m292_am, 
        m300_bm, m300_am, m2, \sha_last_blk_next_0_a4_0\, m15, 
        m108, m267, m242, m146, m111, m76, m70, m45, m29, m273_0, 
        m273_1, m98, m60, GND_net_1, VCC_net_1 : std_logic;

begin 

    hash_control_st_reg_ns_i_0_a2_2(4) <= 
        \hash_control_st_reg_ns_i_0_a2_2[4]\;
    sha_last_blk_next_0_a4_0 <= \sha_last_blk_next_0_a4_0\;

    \next_rout_31_0_.m313\ : CFG4
      generic map(INIT => x"5A2F")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m313);
    
    \next_rout_31_0_.m71\ : CFG3
      generic map(INIT => x"71")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m71);
    
    \next_rout_31_0_.m227\ : CFG3
      generic map(INIT => x"4E")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep1, Y => m227);
    
    \next_rout_31_0_.m13\ : CFG3
      generic map(INIT => x"35")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m13);
    
    \next_rout_31_0_.m285_1_1\ : CFG4
      generic map(INIT => x"A2BD")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(2), C => 
        Kt_addr(1), D => m285_1_1_1, Y => m285_1_1);
    
    \next_rout_31_0_.m216\ : CFG3
      generic map(INIT => x"4A")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep1, Y => m216);
    
    \next_rout_31_0_.m2\ : CFG3
      generic map(INIT => x"09")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m2);
    
    \next_rout_31_0_.m137_am\ : CFG4
      generic map(INIT => x"EBAB")

      port map(A => m304_2, B => m137_am_1_0, C => Kt_addr_3_rep1, 
        D => m129, Y => m137_am);
    
    \next_rout_31_0_.m10_am\ : CFG4
      generic map(INIT => x"BA89")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m10_am);
    
    \next_rout_31_0_.m289\ : CFG3
      generic map(INIT => x"47")

      port map(A => m289_1_1, B => Kt_addr(3), C => m289_1_0, Y
         => m289);
    
    \next_rout_31_0_.m177_1_0\ : CFG4
      generic map(INIT => x"0A1B")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => m174, D
         => pad_one_reg_0_0_a2_0, Y => m177_1_0);
    
    \next_rout_31_0_.m98\ : CFG4
      generic map(INIT => x"3479")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m98);
    
    \next_rout_31_0_.m119_am\ : CFG4
      generic map(INIT => x"DD8D")

      port map(A => Kt_addr_4_rep2, B => m108, C => 
        Kt_addr_0_rep2, D => Kt_addr(1), Y => m119_am);
    
    \next_rout_31_0_.m250_am\ : CFG4
      generic map(INIT => x"0051")

      port map(A => m273_2, B => m250_am_1, C => Kt_addr_3_rep2, 
        D => m48_1, Y => m250_am);
    
    \next_rout_31_0_.m157_1_2\ : CFG4
      generic map(INIT => x"4657")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(5), C => m151, D
         => m148, Y => m157_1_2);
    
    \next_rout_31_0_.m141\ : CFG3
      generic map(INIT => x"FD")

      port map(A => m141_1, B => m211_0, C => m177_1, Y => m141);
    
    \next_rout_31_0_.m235_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m235_bm, C => m235_am, Y => 
        m235_ns);
    
    \next_rout_31_0_.m104_bm_1\ : CFG4
      generic map(INIT => x"41EB")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_0_rep1, D => m79, Y => m104_bm_1);
    
    \next_rout_31_0_.m144_am\ : CFG4
      generic map(INIT => x"0216")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m144_am);
    
    \next_rout_31_0_.m270_1_1\ : CFG4
      generic map(INIT => x"4657")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(5), C => m263, D
         => m261, Y => m270_1_1);
    
    \next_rout_31_0_.m289_1_0\ : CFG3
      generic map(INIT => x"74")

      port map(A => m237, B => Kt_addr(4), C => m46, Y => 
        m289_1_0);
    
    \next_rout_31_0_.m51\ : CFG3
      generic map(INIT => x"15")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m51);
    
    \next_rout_31_0_.m108\ : CFG3
      generic map(INIT => x"10")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m108);
    
    \next_rout_31_0_.m67_am\ : CFG4
      generic map(INIT => x"80D5")

      port map(A => Kt_addr_4_rep1, B => Kt_addr(2), C => 
        Kt_addr(1), D => m63, Y => m67_am);
    
    \next_rout_31_0_.m207_1_1\ : CFG3
      generic map(INIT => x"74")

      port map(A => m205, B => Kt_addr_3_rep2, C => m202, Y => 
        m207_1_1);
    
    \next_rout_31_0_.m168_1_0\ : CFG4
      generic map(INIT => x"2C5A")

      port map(A => Kt_addr_4_rep2, B => Kt_addr_3_rep2, C => 
        m168_1_0_1, D => Kt_addr(0), Y => m168_1_0);
    
    \next_rout_31_0_.m92\ : CFG3
      generic map(INIT => x"6B")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m92);
    
    \next_rout_31_0_.m62_am_1\ : CFG4
      generic map(INIT => x"0A1B")

      port map(A => Kt_addr_fast(4), B => Kt_addr_0_rep1, C => 
        m51, D => hash_control_st_reg_ns_i_0_a2_0(4), Y => 
        m62_am_1);
    
    \next_rout_31_0_.m43\ : CFG3
      generic map(INIT => x"4D")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m43);
    
    \next_rout_31_0_.m73_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => Kt_addr_4_rep1, B => m68, C => Kt_addr_3_rep1, 
        Y => m73);
    
    \next_rout_31_0_.m62_am\ : CFG3
      generic map(INIT => x"72")

      port map(A => Kt_addr_3_rep1, B => m62_am_1_0, C => 
        m62_am_1, Y => m62_am);
    
    \next_rout_31_0_.m316_3\ : CFG4
      generic map(INIT => x"8020")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(4), C => 
        Kt_addr(5), D => m126, Y => m316_2);
    
    \next_rout_31_0_.m40_2\ : CFG3
      generic map(INIT => x"40")

      port map(A => Kt_addr_fast(4), B => m37, C => 
        Kt_addr_fast(3), Y => m78_1);
    
    \next_rout_31_0_.m292_am\ : CFG4
      generic map(INIT => x"E4EE")

      port map(A => Kt_addr(4), B => m54, C => Kt_addr(2), D => 
        Kt_addr(1), Y => m292_am);
    
    \next_rout_31_0_.m114_1_0\ : CFG3
      generic map(INIT => x"47")

      port map(A => m63, B => Kt_addr_3_rep1, C => m35, Y => 
        m114_1_0);
    
    \next_rout_31_0_.m34\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => m32, B => Kt_addr(5), C => m34_1_2, D => m30, 
        Y => m34);
    
    \next_rout_31_0_.m23\ : CFG4
      generic map(INIT => x"75C3")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m23);
    
    \next_rout_31_0_.m166\ : CFG4
      generic map(INIT => x"5214")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_fast(4), C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m166);
    
    \next_rout_31_0_.m202\ : CFG4
      generic map(INIT => x"38BA")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m202);
    
    \next_rout_31_0_.m67_bm\ : CFG4
      generic map(INIT => x"6173")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_0_rep2, C => 
        Kt_addr(2), D => Kt_addr(1), Y => m67_bm);
    
    \next_rout_31_0_.m226_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m226_bm, B => Kt_addr(3), C => m226_am, Y => 
        m226_ns);
    
    \next_rout_31_0_.m137_bm_1_0\ : CFG4
      generic map(INIT => x"5D08")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => m17, Y => m137_bm_1_0);
    
    \next_rout_31_0_.m83_am\ : CFG4
      generic map(INIT => x"52A7")

      port map(A => Kt_addr_4_rep2, B => 
        \sha_last_blk_next_0_a4_0\, C => Kt_addr_0_rep2, D => 
        Kt_addr(1), Y => m83_am);
    
    \next_rout_31_0_.m70\ : CFG3
      generic map(INIT => x"79")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m70);
    
    \next_rout_31_0_.m104_am\ : CFG4
      generic map(INIT => x"1D0C")

      port map(A => Kt_addr_0_rep2, B => Kt_addr_3_rep1, C => m98, 
        D => \sha_last_blk_next_0_a4_0\, Y => m104_am);
    
    \next_rout_31_0_.m308_ns\ : CFG4
      generic map(INIT => x"B964")

      port map(A => Kt_addr(3), B => Kt_addr(4), C => m117, D => 
        m308_ns_1, Y => i3_mux_1);
    
    \next_rout_31_0_.m83_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m83_bm, C => m83_am, Y => 
        m83_ns);
    
    \next_rout_31_0_.m281_am\ : CFG4
      generic map(INIT => x"CD45")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => m15, D => 
        \sha_last_blk_next_0_a4_0\, Y => m281_am);
    
    \next_rout_31_0_.m230\ : CFG4
      generic map(INIT => x"F0F7")

      port map(A => Kt_addr(4), B => Kt_addr(2), C => m230_0, D
         => m230_1_1, Y => m230);
    
    \next_rout_31_0_.m137_bm_1\ : CFG3
      generic map(INIT => x"47")

      port map(A => m133, B => Kt_addr_fast(4), C => m132, Y => 
        m137_bm_1);
    
    \next_rout_31_0_.m310\ : CFG4
      generic map(INIT => x"607C")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m310);
    
    \next_rout_31_0_.m188_1_2\ : CFG4
      generic map(INIT => x"5746")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(5), C => m181, D
         => m180, Y => m188_1_2);
    
    \next_rout_31_0_.m133\ : CFG3
      generic map(INIT => x"29")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m133);
    
    \next_rout_31_0_.m110_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m110_bm, B => Kt_addr(3), C => m110_am, Y => 
        m110_ns);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \next_rout_31_0_.m325_1_0\ : CFG4
      generic map(INIT => x"8F85")

      port map(A => Kt_addr_3_rep1, B => m318, C => m325_1_0_1, D
         => hash_control_st_reg_ns_i_0_a2_0(4), Y => m325_1_0);
    
    \next_rout_31_0_.m250_bm_1_0\ : CFG3
      generic map(INIT => x"CB")

      port map(A => Kt_addr_fast(3), B => Kt_addr_1_rep2, C => 
        m250_bm_1_0_1, Y => m250_bm_1_0);
    
    \next_rout_31_0_.m49_am\ : CFG4
      generic map(INIT => x"0A0D")

      port map(A => Kt_addr_3_rep1, B => Kt_addr_0_rep2, C => 
        m78_1, D => m49_am_1_0, Y => m49_am);
    
    \next_rout_31_0_.m292_bm\ : CFG4
      generic map(INIT => x"280C")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m292_bm);
    
    \next_rout_31_0_.m186\ : CFG4
      generic map(INIT => x"6133")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m186);
    
    \next_rout_31_0_.m60\ : CFG4
      generic map(INIT => x"2B0E")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m60);
    
    \next_rout_31_0_.m49_bm\ : CFG4
      generic map(INIT => x"FFAB")

      port map(A => m48_2, B => m49_bm_1, C => Kt_addr_3_rep1, D
         => m48_1, Y => m49_bm);
    
    \next_rout_31_0_.m177_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_4_rep2, B => m22, C => Kt_addr_3_rep2, 
        Y => m177_2);
    
    \next_rout_31_0_.m15\ : CFG2
      generic map(INIT => x"2")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, Y => m15);
    
    \next_rout_31_0_.m132\ : CFG3
      generic map(INIT => x"3B")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m132);
    
    \next_rout_31_0_.m48_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_fast(4), B => m46, C => 
        Kt_addr_fast(3), Y => m48_2);
    
    \next_rout_31_0_.m114_1\ : CFG3
      generic map(INIT => x"02")

      port map(A => Kt_addr_4_rep1, B => m111, C => 
        Kt_addr_3_rep1, Y => m230_0);
    
    \next_rout_31_0_.m258_bm\ : CFG4
      generic map(INIT => x"72FA")

      port map(A => Kt_addr(4), B => Kt_addr(2), C => m120, D => 
        Kt_addr(0), Y => m258_bm);
    
    \next_rout_31_0_.m237\ : CFG3
      generic map(INIT => x"3E")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m237);
    
    \next_rout_31_0_.m157\ : CFG4
      generic map(INIT => x"38F8")

      port map(A => m155, B => Kt_addr(5), C => m157_1_2, D => 
        m153, Y => m157);
    
    \next_rout_31_0_.m126\ : CFG3
      generic map(INIT => x"6E")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m126);
    
    \next_rout_31_0_.m318\ : CFG3
      generic map(INIT => x"36")

      port map(A => Kt_addr_fast(0), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, Y => m318);
    
    \next_rout_31_0_.m151\ : CFG4
      generic map(INIT => x"7B06")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_fast(4), C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m151);
    
    \next_rout_31_0_.m117\ : CFG3
      generic map(INIT => x"19")

      port map(A => Kt_addr(2), B => Kt_addr(1), C => Kt_addr(0), 
        Y => m117);
    
    \next_rout_31_0_.m111\ : CFG3
      generic map(INIT => x"7A")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m111);
    
    \next_rout_31_0_.m219_1_2\ : CFG4
      generic map(INIT => x"2367")

      port map(A => Kt_addr_3_rep2, B => Kt_addr_4_rep2, C => m68, 
        D => m216, Y => m219_1_2);
    
    \next_rout_31_0_.m155\ : CFG4
      generic map(INIT => x"69DF")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m155);
    
    \next_rout_31_0_.m45\ : CFG3
      generic map(INIT => x"28")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m45);
    
    \next_rout_31_0_.m137_bm\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m137_bm_1_0, B => Kt_addr_3_rep2, C => 
        m137_bm_1, Y => m137_bm);
    
    \next_rout_31_0_.m304_2\ : CFG4
      generic map(INIT => x"0002")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(4), C => 
        Kt_addr(0), D => m1, Y => m304_1);
    
    \next_rout_31_0_.m35\ : CFG3
      generic map(INIT => x"5E")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m35);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \next_rout_31_0_.m103_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_fast(4), B => m29, C => 
        Kt_addr_fast(3), Y => m304_2);
    
    \next_rout_31_0_.m239\ : CFG4
      generic map(INIT => x"3E32")

      port map(A => m237, B => m239_1_2, C => Kt_addr(4), D => 
        m81, Y => m239);
    
    \next_rout_31_0_.m172_bm\ : CFG4
      generic map(INIT => x"6C1E")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m172_bm);
    
    \next_rout_31_0_.m93\ : CFG4
      generic map(INIT => x"3465")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m93);
    
    \next_rout_31_0_.m76\ : CFG3
      generic map(INIT => x"6D")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m76);
    
    \next_rout_31_0_.m197_1_0\ : CFG4
      generic map(INIT => x"41EB")

      port map(A => Kt_addr_3_rep2, B => Kt_addr_4_rep2, C => 
        m185, D => m191, Y => m197_1_0);
    
    \next_rout_31_0_.m17\ : CFG3
      generic map(INIT => x"38")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m17);
    
    \next_rout_31_0_.m10_bm\ : CFG4
      generic map(INIT => x"4427")

      port map(A => Kt_addr(4), B => Kt_addr(2), C => 
        hash_control_st_reg_ns_i_0_a2_0(4), D => Kt_addr(0), Y
         => m10_bm);
    
    \next_rout_31_0_.m215_bm_1_0\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr_4_rep1, B => m90, C => m22, Y => 
        m215_bm_1_0);
    
    \next_rout_31_0_.m266\ : CFG4
      generic map(INIT => x"3733")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m266);
    
    \next_rout_31_0_.m119_bm\ : CFG4
      generic map(INIT => x"3A2D")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m119_bm);
    
    \next_rout_31_0_.m235_bm\ : CFG4
      generic map(INIT => x"7E45")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m235_bm);
    
    \next_rout_31_0_.m292_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m292_bm, C => m292_am, Y => 
        m292_ns);
    
    \next_rout_31_0_.m244_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_fast(3), B => Kt_addr_4_rep1, C => 
        m242, Y => m273_2);
    
    \next_rout_31_0_.m215_bm\ : CFG3
      generic map(INIT => x"74")

      port map(A => m215_bm_1_0, B => Kt_addr_3_rep2, C => 
        m215_bm_1, Y => m215_bm);
    
    \next_rout_31_0_.m276_am\ : CFG4
      generic map(INIT => x"8827")

      port map(A => Kt_addr(4), B => Kt_addr(1), C => 
        pad_one_reg_0_0_a2_0, D => Kt_addr(0), Y => m276_am);
    
    \next_rout_31_0_.m188\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => m186, B => Kt_addr(5), C => m188_1_2, D => 
        m184, Y => Kt_data_0);
    
    \next_rout_31_0_.m177\ : CFG4
      generic map(INIT => x"FFAB")

      port map(A => m177_2, B => Kt_addr(3), C => m177_1_0, D => 
        m177_1, Y => m177);
    
    \next_rout_31_0_.m141_1_0\ : CFG4
      generic map(INIT => x"6E7F")

      port map(A => Kt_addr_4_rep2, B => Kt_addr_3_rep2, C => m79, 
        D => m138, Y => m141_1);
    
    \next_rout_31_0_.m197_1_1\ : CFG3
      generic map(INIT => x"74")

      port map(A => m195, B => Kt_addr_3_rep2, C => m193, Y => 
        m197_1_1);
    
    \next_rout_31_0_.m300_bm\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(4), B => m146, C => Kt_addr(2), Y => 
        m300_bm);
    
    \next_rout_31_0_.m261\ : CFG4
      generic map(INIT => x"573C")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m261);
    
    \next_rout_31_0_.m258_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m258_bm, C => m258_am, Y => 
        m258_ns);
    
    \next_rout_31_0_.m168_1_1\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr_3_rep2, B => m166, C => m163, Y => 
        m168_1_1);
    
    \next_rout_31_0_.m153\ : CFG4
      generic map(INIT => x"0A10")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m153);
    
    \next_rout_31_0_.m79\ : CFG3
      generic map(INIT => x"3D")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m79);
    
    \next_rout_31_0_.m273\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => m273_1, B => m273_0, C => m273_2, D => m73, Y
         => m273);
    
    \next_rout_31_0_.m141_1\ : CFG4
      generic map(INIT => x"0040")

      port map(A => Kt_addr_fast(3), B => Kt_addr_4_rep1, C => 
        Kt_addr_0_rep1, D => hash_control_st_reg_ns_i_0_a2_0(4), 
        Y => m211_0);
    
    \next_rout_31_0_.m34_1_2\ : CFG4
      generic map(INIT => x"4657")

      port map(A => Kt_addr_3_rep1, B => Kt_addr(5), C => i2_mux, 
        D => m23, Y => m34_1_2);
    
    \next_rout_31_0_.m119_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m119_bm, C => m119_am, Y => 
        m119_ns);
    
    \next_rout_31_0_.m110_am\ : CFG4
      generic map(INIT => x"E710")

      port map(A => Kt_addr(1), B => Kt_addr_4_rep2, C => 
        Kt_addr_0_rep2, D => Kt_addr(2), Y => m110_am);
    
    \next_rout_31_0_.m296\ : CFG4
      generic map(INIT => x"AEEE")

      port map(A => m296_2, B => m296_1_1, C => Kt_addr(3), D => 
        m16, Y => m296);
    
    \next_rout_31_0_.m321\ : CFG2
      generic map(INIT => x"2")

      port map(A => hash_control_st_reg_ns_i_0_a2_0(4), B => 
        Kt_addr(4), Y => \hash_control_st_reg_ns_i_0_a2_2[4]\);
    
    \next_rout_31_0_.m114\ : CFG4
      generic map(INIT => x"FAFB")

      port map(A => m230_0, B => Kt_addr(4), C => m296_2, D => 
        m114_1_0, Y => m114);
    
    \next_rout_31_0_.m103_2\ : CFG3
      generic map(INIT => x"10")

      port map(A => Kt_addr_fast(4), B => m22, C => 
        Kt_addr_fast(3), Y => m103_1);
    
    \next_rout_31_0_.m67_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m67_bm, C => m67_am, Y => 
        m67_ns);
    
    \next_rout_31_0_.m95_1_0\ : CFG4
      generic map(INIT => x"7520")

      port map(A => Kt_addr_3_rep1, B => Kt_addr_4_rep2, C => m46, 
        D => m87, Y => m95_1_0);
    
    \next_rout_31_0_.m78\ : CFG4
      generic map(INIT => x"FFAB")

      port map(A => m78_2, B => Kt_addr(3), C => m78_1_0, D => 
        m78_1, Y => m78);
    
    \next_rout_31_0_.m37\ : CFG3
      generic map(INIT => x"51")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m37);
    
    \next_rout_31_0_.m207_1_0\ : CFG4
      generic map(INIT => x"67C2")

      port map(A => Kt_addr_4_rep2, B => m207_1_0_1, C => 
        Kt_addr(2), D => Kt_addr(1), Y => m207_1_0);
    
    \next_rout_31_0_.m105\ : CFG3
      generic map(INIT => x"65")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m105);
    
    \next_rout_31_0_.m19_1_0\ : CFG4
      generic map(INIT => x"1B4E")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => m13, D => 
        pad_one_reg_0_0_a2_0, Y => m19_1_0);
    
    \next_rout_31_0_.m250_am_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => Kt_addr_4_rep1, B => m194, C => m85, Y => 
        m250_am_1);
    
    \next_rout_31_0_.m30\ : CFG4
      generic map(INIT => x"4B1D")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_0_rep2, C => 
        Kt_addr(2), D => Kt_addr(1), Y => m30);
    
    \next_rout_31_0_.m276_bm\ : CFG4
      generic map(INIT => x"5ABE")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m276_bm);
    
    \next_rout_31_0_.m83_bm\ : CFG4
      generic map(INIT => x"0398")

      port map(A => Kt_addr(1), B => Kt_addr_4_rep2, C => 
        Kt_addr_0_rep2, D => Kt_addr(2), Y => m83_bm);
    
    \next_rout_31_0_.m323\ : CFG4
      generic map(INIT => x"4202")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m323);
    
    \next_rout_31_0_.m95_1_1\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr_3_rep1, B => m93, C => m91, Y => 
        m95_1_1);
    
    \next_rout_31_0_.m270\ : CFG4
      generic map(INIT => x"EBAB")

      port map(A => m270_2, B => m270_1_1, C => Kt_addr(5), D => 
        m266, Y => Kt_data_9);
    
    \next_rout_31_0_.m174\ : CFG3
      generic map(INIT => x"64")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep1, Y => m174);
    
    \next_rout_31_0_.m146\ : CFG3
      generic map(INIT => x"1B")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m146);
    
    \next_rout_31_0_.m273_1\ : CFG4
      generic map(INIT => x"0440")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(4), C => 
        Kt_addr(0), D => m15, Y => m273_0);
    
    \next_rout_31_0_.m68\ : CFG3
      generic map(INIT => x"3E")

      port map(A => Kt_addr_fast(0), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, Y => m68);
    
    \next_rout_31_0_.m114_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_4_rep1, B => m81, C => Kt_addr_3_rep1, 
        Y => m296_2);
    
    \next_rout_31_0_.m62_am_1_0\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr_fast(4), B => m54, C => m53, Y => 
        m62_am_1_0);
    
    \next_rout_31_0_.m144_bm\ : CFG4
      generic map(INIT => x"F5E4")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => m85, D
         => hash_control_st_reg_ns_i_0_a2_0(4), Y => m144_bm);
    
    \next_rout_31_0_.m316_1_1\ : CFG4
      generic map(INIT => x"3726")

      port map(A => Kt_addr(5), B => Kt_addr_3_rep2, C => m311, D
         => m310, Y => m316_1_1);
    
    \next_rout_31_0_.m304\ : CFG4
      generic map(INIT => x"FFDC")

      port map(A => Kt_addr(3), B => m304_2, C => m304_1_0, D => 
        m304_1, Y => m304);
    
    \next_rout_31_0_.m215_bm_1\ : CFG4
      generic map(INIT => x"01AB")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep2, D => m164, Y => m215_bm_1);
    
    \next_rout_31_0_.m325\ : CFG4
      generic map(INIT => x"04BF")

      port map(A => Kt_addr(3), B => Kt_addr(5), C => 
        \hash_control_st_reg_ns_i_0_a2_2[4]\, D => m325_1_1, Y
         => m325);
    
    \next_rout_31_0_.m254_1_1\ : CFG3
      generic map(INIT => x"72")

      port map(A => Kt_addr_4_rep2, B => m252, C => m232, Y => 
        m254_1_1);
    
    \next_rout_31_0_.m219\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => m127, B => Kt_addr(3), C => m219_1_2, D => 
        m51, Y => m219);
    
    \next_rout_31_0_.m91\ : CFG4
      generic map(INIT => x"774B")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m91);
    
    \next_rout_31_0_.m273_2\ : CFG3
      generic map(INIT => x"20")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(4), C => m81, Y
         => m273_1);
    
    \next_rout_31_0_.m16\ : CFG3
      generic map(INIT => x"5B")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m16);
    
    \next_rout_31_0_.m78_3\ : CFG3
      generic map(INIT => x"80")

      port map(A => Kt_addr_4_rep2, B => m76, C => Kt_addr_3_rep1, 
        Y => m78_2);
    
    \next_rout_31_0_.m110_bm\ : CFG3
      generic map(INIT => x"64")

      port map(A => Kt_addr_4_rep2, B => m2, C => 
        pad_one_reg_0_0_a2_0, Y => m110_bm);
    
    \next_rout_31_0_.m48_2\ : CFG3
      generic map(INIT => x"40")

      port map(A => Kt_addr_fast(4), B => m45, C => 
        Kt_addr_fast(3), Y => m48_1);
    
    \next_rout_31_0_.m85\ : CFG3
      generic map(INIT => x"59")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m85);
    
    \next_rout_31_0_.m325_1_0_1\ : CFG4
      generic map(INIT => x"5456")

      port map(A => Kt_addr_fast(4), B => Kt_addr_fast(3), C => 
        Kt_addr_1_rep1, D => Kt_addr_2_rep1, Y => m325_1_0_1);
    
    \next_rout_31_0_.m250_bm_1_0_1\ : CFG4
      generic map(INIT => x"523F")

      port map(A => Kt_addr_fast(4), B => Kt_addr_fast(0), C => 
        Kt_addr_fast(2), D => Kt_addr_fast(1), Y => m250_bm_1_0_1);
    
    \next_rout_31_0_.m81\ : CFG3
      generic map(INIT => x"46")

      port map(A => Kt_addr_fast(0), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, Y => m81);
    
    \next_rout_31_0_.m276_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m276_bm, C => m276_am, Y => 
        m276_ns);
    
    \next_rout_31_0_.m172_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m172_bm, C => m172_am, Y => 
        m172_ns);
    
    \next_rout_31_0_.m285_1_1_1\ : CFG4
      generic map(INIT => x"100E")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_3_rep1, C => 
        Kt_addr_0_rep2, D => Kt_addr_1_rep2, Y => m285_1_1_1);
    
    \next_rout_31_0_.m19\ : CFG3
      generic map(INIT => x"72")

      port map(A => Kt_addr(3), B => m19_1_1, C => m19_1_0, Y => 
        m19);
    
    \next_rout_31_0_.m104_bm\ : CFG4
      generic map(INIT => x"FFAB")

      port map(A => m304_2, B => Kt_addr_3_rep1, C => m104_bm_1, 
        D => m103_1, Y => m104_bm);
    
    \next_rout_31_0_.m168_1_0_1\ : CFG4
      generic map(INIT => x"083D")

      port map(A => Kt_addr_fast(4), B => Kt_addr_fast(3), C => 
        Kt_addr_1_rep2, D => Kt_addr_2_rep2, Y => m168_1_0_1);
    
    \next_rout_31_0_.m263\ : CFG4
      generic map(INIT => x"7840")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m263);
    
    \next_rout_31_0_.m300_am\ : CFG4
      generic map(INIT => x"6C6A")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => Kt_addr(2), 
        D => Kt_addr(1), Y => m300_am);
    
    \next_rout_31_0_.m205\ : CFG4
      generic map(INIT => x"615F")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m205);
    
    \next_rout_31_0_.m46\ : CFG3
      generic map(INIT => x"1D")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m46);
    
    \next_rout_31_0_.m207_1_0_1\ : CFG4
      generic map(INIT => x"15AC")

      port map(A => Kt_addr_fast(3), B => Kt_addr_4_rep1, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m207_1_0_1);
    
    \next_rout_31_0_.m26\ : CFG4
      generic map(INIT => x"43A5")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => i2_mux);
    
    \next_rout_31_0_.m235_am\ : CFG4
      generic map(INIT => x"E4B1")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => m232, D
         => hash_control_st_reg_ns_i_0_a2_0(4), Y => m235_am);
    
    \next_rout_31_0_.m230_1_0\ : CFG4
      generic map(INIT => x"0B5B")

      port map(A => Kt_addr_4_rep2, B => m227, C => 
        Kt_addr_3_rep2, D => Kt_addr(1), Y => m230_1_1);
    
    \next_rout_31_0_.m316\ : CFG4
      generic map(INIT => x"EEAE")

      port map(A => m316_2, B => m316_1_1, C => Kt_addr(5), D => 
        m313, Y => m316);
    
    \next_rout_31_0_.m222_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m222_bm, B => Kt_addr(3), C => m222_am, Y => 
        m222_ns);
    
    \next_rout_31_0_.m191\ : CFG4
      generic map(INIT => x"14CE")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m191);
    
    \next_rout_31_0_.m10_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m10_bm, B => Kt_addr(3), C => m10_am, Y => 
        m10_ns);
    
    \next_rout_31_0_.m148\ : CFG4
      generic map(INIT => x"3250")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_fast(4), C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m148);
    
    \next_rout_31_0_.m144_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m144_bm, B => Kt_addr(3), C => m144_am, Y => 
        m144_ns);
    
    \next_rout_31_0_.m296_1_1\ : CFG4
      generic map(INIT => x"2367")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(4), C => m237, D
         => hash_control_st_reg_ns_i_0_a2_0(4), Y => m296_1_1);
    
    \next_rout_31_0_.m215_am\ : CFG4
      generic map(INIT => x"DDCD")

      port map(A => m215_am_1_0, B => m211_0, C => Kt_addr_4_rep2, 
        D => m209, Y => m215_am);
    
    \next_rout_31_0_.m138\ : CFG3
      generic map(INIT => x"3A")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m138);
    
    \next_rout_31_0_.m49_am_1_0\ : CFG4
      generic map(INIT => x"4657")

      port map(A => Kt_addr_fast(4), B => Kt_addr_fast(3), C => 
        m35, D => Kt_addr_1_rep1, Y => m49_am_1_0);
    
    \next_rout_31_0_.m222_am\ : CFG4
      generic map(INIT => x"A7F4")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m222_am);
    
    \next_rout_31_0_.m209\ : CFG3
      generic map(INIT => x"21")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m209);
    
    \next_rout_31_0_.m325_1_1\ : CFG3
      generic map(INIT => x"1D")

      port map(A => m325_1_0, B => Kt_addr(5), C => m323, Y => 
        m325_1_1);
    
    \next_rout_31_0_.m90\ : CFG3
      generic map(INIT => x"53")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m90);
    
    \next_rout_31_0_.m195\ : CFG4
      generic map(INIT => x"596C")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m195);
    
    \next_rout_31_0_.m87\ : CFG4
      generic map(INIT => x"1B41")

      port map(A => Kt_addr_fast(4), B => Kt_addr_2_rep1, C => 
        Kt_addr_1_rep1, D => Kt_addr_0_rep1, Y => m87);
    
    \next_rout_31_0_.m254_1_0\ : CFG4
      generic map(INIT => x"058D")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => m105, D
         => m1, Y => m254_1_0);
    
    \next_rout_31_0_.m250_bm\ : CFG4
      generic map(INIT => x"20FD")

      port map(A => Kt_addr_3_rep2, B => Kt_addr_4_rep2, C => 
        m132, D => m250_bm_1_0, Y => m250_bm);
    
    \next_rout_31_0_.m181\ : CFG4
      generic map(INIT => x"2E11")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_4_rep1, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m181);
    
    \next_rout_31_0_.m129\ : CFG3
      generic map(INIT => x"4E")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m129);
    
    \next_rout_31_0_.m29\ : CFG3
      generic map(INIT => x"54")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m29);
    
    \next_rout_31_0_.m242\ : CFG3
      generic map(INIT => x"4A")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m242);
    
    \next_rout_31_0_.m232\ : CFG3
      generic map(INIT => x"45")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m232);
    
    \next_rout_31_0_.m172_am\ : CFG4
      generic map(INIT => x"111B")

      port map(A => Kt_addr_4_rep2, B => m133, C => Kt_addr(2), D
         => Kt_addr(1), Y => m172_am);
    
    \next_rout_31_0_.m163\ : CFG4
      generic map(INIT => x"12AD")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_fast(4), C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m163);
    
    \next_rout_31_0_.m73\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => m73_1, B => Kt_addr(4), C => m73_1_0, D => 
        m73, Y => m73_0);
    
    \next_rout_31_0_.m215_am_1_0\ : CFG4
      generic map(INIT => x"5746")

      port map(A => Kt_addr_fast(3), B => Kt_addr_4_rep1, C => 
        m92, D => m53, Y => m215_am_1_0);
    
    \next_rout_31_0_.m185\ : CFG3
      generic map(INIT => x"87")

      port map(A => Kt_addr_1_rep2, B => Kt_addr_2_rep2, C => 
        Kt_addr_0_rep1, Y => m185);
    
    \next_rout_31_0_.m164\ : CFG3
      generic map(INIT => x"64")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m164);
    
    \next_rout_31_0_.m300_ns\ : CFG3
      generic map(INIT => x"B8")

      port map(A => m300_bm, B => Kt_addr(3), C => m300_am, Y => 
        m300_ns);
    
    \next_rout_31_0_.m78_1_0\ : CFG4
      generic map(INIT => x"5D08")

      port map(A => Kt_addr_4_rep1, B => Kt_addr(2), C => 
        Kt_addr(1), D => m28, Y => m78_1_0);
    
    \next_rout_31_0_.m127\ : CFG3
      generic map(INIT => x"36")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m127);
    
    \next_rout_31_0_.m270_3\ : CFG4
      generic map(INIT => x"2000")

      port map(A => Kt_addr_3_rep2, B => Kt_addr(4), C => 
        Kt_addr(5), D => m267, Y => m270_2);
    
    \next_rout_31_0_.m226_am\ : CFG4
      generic map(INIT => x"F4DE")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m226_am);
    
    \next_rout_31_0_.m28\ : CFG3
      generic map(INIT => x"68")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m28);
    
    \next_rout_31_0_.m304_1_0\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr(4), B => m216, C => m133, Y => 
        m304_1_0);
    
    \next_rout_31_0_.m137_am_1_0\ : CFG4
      generic map(INIT => x"3276")

      port map(A => Kt_addr_fast(3), B => Kt_addr_fast(4), C => 
        m126, D => m127, Y => m137_am_1_0);
    
    \next_rout_31_0_.m254\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr(3), B => m254_1_1, C => m254_1_0, Y
         => m254);
    
    \next_rout_31_0_.m62_bm\ : CFG4
      generic map(INIT => x"BE14")

      port map(A => Kt_addr_3_rep1, B => Kt_addr_0_rep2, C => 
        Kt_addr(1), D => m60, Y => m62_bm);
    
    \next_rout_31_0_.m258_am\ : CFG3
      generic map(INIT => x"38")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => m1, Y
         => m258_am);
    
    \next_rout_31_0_.m222_bm\ : CFG3
      generic map(INIT => x"67")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        \sha_last_blk_next_0_a4_0\, Y => m222_bm);
    
    \next_rout_31_0_.m193\ : CFG4
      generic map(INIT => x"0301")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m193);
    
    \next_rout_31_0_.m141_2\ : CFG3
      generic map(INIT => x"10")

      port map(A => Kt_addr_4_rep2, B => m90, C => Kt_addr_3_rep1, 
        Y => m177_1);
    
    \next_rout_31_0_.m42\ : CFG2
      generic map(INIT => x"4")

      port map(A => Kt_addr_1_rep1, B => Kt_addr_2_rep1, Y => 
        \sha_last_blk_next_0_a4_0\);
    
    \next_rout_31_0_.m194\ : CFG3
      generic map(INIT => x"26")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m194);
    
    \next_rout_31_0_.m54\ : CFG3
      generic map(INIT => x"14")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m54);
    
    \next_rout_31_0_.m53\ : CFG3
      generic map(INIT => x"25")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m53);
    
    \next_rout_31_0_.m281_bm\ : CFG3
      generic map(INIT => x"8B")

      port map(A => m51, B => Kt_addr(4), C => m15, Y => m281_bm);
    
    \next_rout_31_0_.m239_1_2\ : CFG4
      generic map(INIT => x"193B")

      port map(A => Kt_addr_4_rep2, B => Kt_addr_3_rep2, C => 
        m105, D => m227, Y => m239_1_2);
    
    \next_rout_31_0_.m267\ : CFG3
      generic map(INIT => x"42")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m267);
    
    \next_rout_31_0_.m63\ : CFG3
      generic map(INIT => x"4C")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m63);
    
    \next_rout_31_0_.m22\ : CFG3
      generic map(INIT => x"49")

      port map(A => Kt_addr_fast(2), B => Kt_addr_fast(1), C => 
        Kt_addr_fast(0), Y => m22);
    
    \next_rout_31_0_.m32\ : CFG4
      generic map(INIT => x"5B51")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_0_rep2, C => 
        Kt_addr(2), D => Kt_addr(1), Y => m32);
    
    \next_rout_31_0_.m73_2\ : CFG3
      generic map(INIT => x"40")

      port map(A => Kt_addr_4_rep1, B => m70, C => Kt_addr_3_rep1, 
        Y => m73_1);
    
    \next_rout_31_0_.m184\ : CFG4
      generic map(INIT => x"3882")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(0), C => 
        Kt_addr(2), D => Kt_addr(1), Y => m184);
    
    \next_rout_31_0_.m226_bm\ : CFG4
      generic map(INIT => x"66A5")

      port map(A => Kt_addr_4_rep2, B => Kt_addr(2), C => 
        pad_one_reg_0_0_a2_0, D => Kt_addr(0), Y => m226_bm);
    
    \next_rout_31_0_.m124_1_2\ : CFG4
      generic map(INIT => x"2367")

      port map(A => Kt_addr_4_rep2, B => Kt_addr_3_rep1, C => 
        m120, D => m122, Y => m124_1_2);
    
    \next_rout_31_0_.m180\ : CFG4
      generic map(INIT => x"270D")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_4_rep1, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep1, Y => m180);
    
    \next_rout_31_0_.m289_1_1\ : CFG4
      generic map(INIT => x"4E5F")

      port map(A => Kt_addr(4), B => Kt_addr(0), C => m37, D => 
        m1, Y => m289_1_1);
    
    \next_rout_31_0_.m308_ns_1\ : CFG4
      generic map(INIT => x"33B1")

      port map(A => Kt_addr(4), B => Kt_addr(1), C => m1, D => 
        Kt_addr(0), Y => m308_ns_1);
    
    \next_rout_31_0_.m1\ : CFG2
      generic map(INIT => x"9")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep1, Y => m1);
    
    \next_rout_31_0_.m311\ : CFG4
      generic map(INIT => x"580D")

      port map(A => Kt_addr_4_rep1, B => Kt_addr_2_rep2, C => 
        Kt_addr_1_rep2, D => Kt_addr_0_rep2, Y => m311);
    
    \next_rout_31_0_.m19_1_1\ : CFG3
      generic map(INIT => x"27")

      port map(A => Kt_addr(4), B => m17, C => m16, Y => m19_1_1);
    
    \next_rout_31_0_.m124\ : CFG4
      generic map(INIT => x"4F43")

      port map(A => m90, B => Kt_addr(4), C => m124_1_2, D => m16, 
        Y => m124);
    
    \next_rout_31_0_.m73_1_0\ : CFG4
      generic map(INIT => x"41EB")

      port map(A => Kt_addr_3_rep1, B => Kt_addr_0_rep2, C => 
        Kt_addr(1), D => m71, Y => m73_1_0);
    
    \next_rout_31_0_.m120\ : CFG3
      generic map(INIT => x"23")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m120);
    
    \next_rout_31_0_.m281_ns\ : CFG3
      generic map(INIT => x"D8")

      port map(A => Kt_addr(3), B => m281_bm, C => m281_am, Y => 
        m281_ns);
    
    \next_rout_31_0_.m49_bm_1\ : CFG4
      generic map(INIT => x"0A4E")

      port map(A => Kt_addr_fast(4), B => Kt_addr_0_rep1, C => 
        m43, D => hash_control_st_reg_ns_i_0_a2_0(4), Y => 
        m49_bm_1);
    
    \next_rout_31_0_.m122\ : CFG3
      generic map(INIT => x"34")

      port map(A => Kt_addr_2_rep1, B => Kt_addr_1_rep1, C => 
        Kt_addr_0_rep1, Y => m122);
    
    \next_rout_31_0_.m285\ : CFG4
      generic map(INIT => x"02DF")

      port map(A => Kt_addr(3), B => Kt_addr(4), C => m28, D => 
        m285_1_1, Y => m285);
    
    \next_rout_31_0_.m252\ : CFG3
      generic map(INIT => x"2A")

      port map(A => Kt_addr_2_rep2, B => Kt_addr_1_rep2, C => 
        Kt_addr_0_rep2, Y => m252);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity gv_sha256 is

    port( reg_17x32_0_valid_bytes_0                 : in    std_logic_vector(1 downto 0);
          di_o_0                                    : out   std_logic_vector(1 to 1);
          SHA256_BLOCK_0_H0_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o                       : out   std_logic_vector(31 downto 0);
          state_0                                   : in    std_logic;
          state_2                                   : in    std_logic;
          state_3                                   : in    std_logic;
          sha256_controller_0_di_o_3                : in    std_logic;
          sha256_controller_0_di_o_5                : in    std_logic;
          sha256_controller_0_di_o_0                : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0      : in    std_logic;
          SHA256_Module_0_di_req_o                  : out   std_logic;
          SHA256_BLOCK_0_do_valid_o                 : out   std_logic;
          SHA256_Module_0_waiting_data              : in    std_logic;
          SHA256_Module_0_data_available_lastbank_8 : in    std_logic;
          N_484                                     : in    std_logic;
          bytes_sel                                 : in    std_logic;
          SHA256_Module_0_error_o                   : out   std_logic;
          SHA256_BLOCK_0_start_o                    : in    std_logic;
          N_1702                                    : in    std_logic;
          N_1710                                    : in    std_logic;
          ren_pos                                   : in    std_logic;
          N_1690                                    : in    std_logic;
          N_1691                                    : in    std_logic;
          N_1693                                    : in    std_logic;
          N_1692                                    : in    std_logic;
          N_1718                                    : in    std_logic;
          N_1694                                    : in    std_logic;
          N_1698                                    : in    std_logic;
          N_1701                                    : in    std_logic;
          N_1696                                    : in    std_logic;
          N_1697                                    : in    std_logic;
          N_1695                                    : in    std_logic;
          N_1699                                    : in    std_logic;
          N_1707                                    : in    std_logic;
          N_1708                                    : in    std_logic;
          N_1709                                    : in    std_logic;
          N_1706                                    : in    std_logic;
          N_1704                                    : in    std_logic;
          N_1688                                    : in    std_logic;
          N_1687                                    : in    std_logic;
          N_1689                                    : in    std_logic;
          N_1713                                    : in    std_logic;
          N_1716                                    : in    std_logic;
          N_1712                                    : in    std_logic;
          N_1717                                    : in    std_logic;
          N_1715                                    : in    std_logic;
          N_1711                                    : in    std_logic;
          N_1714                                    : in    std_logic
        );

end gv_sha256;

architecture DEF_ARCH of gv_sha256 is 

  component sha256_control
    port( hash_control_st_reg_i                     : out   std_logic_vector(6 to 6);
          msg_bitlen                                : out   std_logic_vector(63 downto 3);
          Kt_addr                                   : out   std_logic_vector(5 downto 0);
          Kt_addr_fast                              : out   std_logic_vector(4 downto 0);
          state                                     : in    std_logic_vector(1 to 1) := (others => 'U');
          hash_control_st_reg_ns_i_0_a2_0           : out   std_logic_vector(4 to 4);
          reg_17x32_0_valid_bytes_0                 : in    std_logic_vector(1 downto 0) := (others => 'U');
          hash_control_st_reg_ns_i_0_a2_2           : in    std_logic_vector(4 to 4) := (others => 'U');
          hash_control_st_reg_2                     : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0      : in    std_logic := 'U';
          one_insert                                : out   std_logic;
          sha_last_blk_reg                          : out   std_logic;
          SHA256_Module_0_di_req_o                  : out   std_logic;
          SHA256_BLOCK_0_do_valid_o                 : out   std_logic;
          Kt_addr_1_rep1                            : out   std_logic;
          Kt_addr_1_rep2                            : out   std_logic;
          Kt_addr_2_rep1                            : out   std_logic;
          Kt_addr_2_rep2                            : out   std_logic;
          Kt_addr_0_rep1                            : out   std_logic;
          Kt_addr_0_rep2                            : out   std_logic;
          Kt_addr_4_rep1                            : out   std_logic;
          Kt_addr_4_rep2                            : out   std_logic;
          Kt_addr_3_rep1                            : out   std_logic;
          Kt_addr_3_rep2                            : out   std_logic;
          N_112                                     : out   std_logic;
          SHA256_Module_0_waiting_data              : in    std_logic := 'U';
          N_223                                     : out   std_logic;
          N_361                                     : out   std_logic;
          N_102                                     : out   std_logic;
          SHA256_Module_0_data_available_lastbank_8 : in    std_logic := 'U';
          N_168_i_0                                 : out   std_logic;
          pad_one_reg_0_0_a2_0                      : out   std_logic;
          oregs_ce_i_a2_0_a2                        : out   std_logic;
          sha_last_blk_next_0_o2_2_out_0            : out   std_logic;
          N_484                                     : in    std_logic := 'U';
          bytes_sel                                 : in    std_logic := 'U';
          sha_last_blk_next_0_a4_0                  : in    std_logic := 'U';
          N_388                                     : in    std_logic := 'U';
          N_111                                     : out   std_logic;
          core_ce_o_iv_i_0                          : out   std_logic;
          N_244_i_0                                 : out   std_logic;
          SHA256_Module_0_error_o                   : out   std_logic;
          ld_i_i_3                                  : out   std_logic;
          SHA256_BLOCK_0_start_o                    : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component sha256_hash_core
    port( R1_data                              : out   std_logic_vector(31 downto 0);
          R2_data                              : out   std_logic_vector(31 downto 0);
          R3_data                              : out   std_logic_vector(31 downto 0);
          R5_data                              : out   std_logic_vector(31 downto 0);
          R6_data                              : out   std_logic_vector(31 downto 0);
          R7_data                              : out   std_logic_vector(31 downto 0);
          R0_data                              : out   std_logic_vector(31 downto 0);
          R4_data                              : out   std_logic_vector(31 downto 0);
          N4_data                              : in    std_logic_vector(31 downto 1) := (others => 'U');
          N0_data                              : in    std_logic_vector(31 downto 1) := (others => 'U');
          W_out_i_1                            : in    std_logic_vector(0 to 0) := (others => 'U');
          Kt_addr                              : in    std_logic_vector(5 to 5) := (others => 'U');
          N3_data                              : in    std_logic_vector(31 downto 1) := (others => 'U');
          N2_data                              : in    std_logic_vector(31 downto 1) := (others => 'U');
          N1_data                              : in    std_logic_vector(31 downto 1) := (others => 'U');
          N7_data                              : in    std_logic_vector(31 downto 1) := (others => 'U');
          N6_data                              : in    std_logic_vector(31 downto 1) := (others => 'U');
          N5_data                              : in    std_logic_vector(31 downto 1) := (others => 'U');
          Wt_data                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          Kt_data_0                            : in    std_logic := 'U';
          Kt_data_9                            : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          core_ce_o_iv_i_0                     : in    std_logic := 'U';
          oregs_ce_i_a2_0_a2                   : in    std_logic := 'U';
          next_reg_H4_cry_0_0_Y                : in    std_logic := 'U';
          next_reg_H0_cry_0_0_Y                : in    std_logic := 'U';
          next_r0_0_cry_0_Y                    : in    std_logic := 'U';
          ld_i_i_3                             : in    std_logic := 'U';
          N_98                                 : in    std_logic := 'U';
          m34                                  : in    std_logic := 'U';
          m49_am                               : in    std_logic := 'U';
          m49_bm                               : in    std_logic := 'U';
          m62_am                               : in    std_logic := 'U';
          m62_bm                               : in    std_logic := 'U';
          m67_ns                               : in    std_logic := 'U';
          m73                                  : in    std_logic := 'U';
          m78                                  : in    std_logic := 'U';
          m83_ns                               : in    std_logic := 'U';
          m95_1_0                              : in    std_logic := 'U';
          m95_1_1                              : in    std_logic := 'U';
          m104_am                              : in    std_logic := 'U';
          m104_bm                              : in    std_logic := 'U';
          m110_ns                              : in    std_logic := 'U';
          m114                                 : in    std_logic := 'U';
          m119_ns                              : in    std_logic := 'U';
          m124                                 : in    std_logic := 'U';
          m137_am                              : in    std_logic := 'U';
          m137_bm                              : in    std_logic := 'U';
          m141                                 : in    std_logic := 'U';
          m144_ns                              : in    std_logic := 'U';
          m157                                 : in    std_logic := 'U';
          m168_1_0                             : in    std_logic := 'U';
          m168_1_1                             : in    std_logic := 'U';
          m172_ns                              : in    std_logic := 'U';
          m177                                 : in    std_logic := 'U';
          m197_1_0                             : in    std_logic := 'U';
          m197_1_1                             : in    std_logic := 'U';
          m207_1_0                             : in    std_logic := 'U';
          m207_1_1                             : in    std_logic := 'U';
          m215_am                              : in    std_logic := 'U';
          m215_bm                              : in    std_logic := 'U';
          m219                                 : in    std_logic := 'U';
          m222_ns                              : in    std_logic := 'U';
          m226_ns                              : in    std_logic := 'U';
          m230                                 : in    std_logic := 'U';
          m235_ns                              : in    std_logic := 'U';
          m239                                 : in    std_logic := 'U';
          m250_am                              : in    std_logic := 'U';
          m250_bm                              : in    std_logic := 'U';
          m254                                 : in    std_logic := 'U';
          m258_ns                              : in    std_logic := 'U';
          m273                                 : in    std_logic := 'U';
          m276_ns                              : in    std_logic := 'U';
          m281_ns                              : in    std_logic := 'U';
          m285                                 : in    std_logic := 'U';
          m289                                 : in    std_logic := 'U';
          m292_ns                              : in    std_logic := 'U';
          m296                                 : in    std_logic := 'U';
          m300_ns                              : in    std_logic := 'U';
          m304                                 : in    std_logic := 'U';
          i3_mux_1                             : in    std_logic := 'U';
          m325                                 : in    std_logic := 'U';
          m316                                 : in    std_logic := 'U';
          next_reg_H3_cry_0_0_Y                : in    std_logic := 'U';
          next_reg_H2_cry_0_0_Y                : in    std_logic := 'U';
          next_reg_H1_cry_0_0_Y                : in    std_logic := 'U';
          next_reg_H7_cry_0_0_Y                : in    std_logic := 'U';
          next_reg_H6_cry_0_0_Y                : in    std_logic := 'U';
          next_reg_H5_cry_0_0_Y                : in    std_logic := 'U';
          m10_ns                               : in    std_logic := 'U';
          m19                                  : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component sha256_regs
    port( SHA256_BLOCK_0_H0_o                  : out   std_logic_vector(31 downto 0);
          N0_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H1_o                  : out   std_logic_vector(31 downto 0);
          N1_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H2_o                  : out   std_logic_vector(31 downto 0);
          N2_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H3_o                  : out   std_logic_vector(31 downto 0);
          N3_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H4_o                  : out   std_logic_vector(31 downto 0);
          N4_data                              : out   std_logic_vector(31 downto 1);
          N5_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H5_o                  : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o                  : out   std_logic_vector(31 downto 0);
          N6_data                              : out   std_logic_vector(31 downto 1);
          SHA256_BLOCK_0_H7_o                  : out   std_logic_vector(31 downto 0);
          N7_data                              : out   std_logic_vector(31 downto 1);
          hash_control_st_reg_i                : in    std_logic_vector(6 to 6) := (others => 'U');
          R0_data                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          R1_data                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          R2_data                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          R3_data                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          R4_data                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          R5_data                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          R6_data                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          R7_data                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          N_168_i_0                            : in    std_logic := 'U';
          next_reg_H0_cry_0_0_Y                : out   std_logic;
          next_reg_H1_cry_0_0_Y                : out   std_logic;
          next_reg_H2_cry_0_0_Y                : out   std_logic;
          next_reg_H3_cry_0_0_Y                : out   std_logic;
          next_reg_H4_cry_0_0_Y                : out   std_logic;
          next_reg_H5_cry_0_0_Y                : out   std_logic;
          next_reg_H6_cry_0_0_Y                : out   std_logic;
          next_reg_H7_cry_0_0_Y                : out   std_logic
        );
  end component;

  component sha256_padding
    port( di_o_0                                    : out   std_logic_vector(1 to 1);
          reg_17x32_0_valid_bytes_0                 : in    std_logic_vector(1 downto 0) := (others => 'U');
          Kt_addr_fast                              : in    std_logic_vector(0 to 0) := (others => 'U');
          hash_control_st_reg                       : in    std_logic_vector(2 to 2) := (others => 'U');
          W_out_2_0                                 : out   std_logic_vector(5 to 5);
          W_out_i_i_2                               : out   std_logic_vector(31 to 31);
          W_out_i_i_1                               : out   std_logic_vector(31 to 31);
          W_out_i_1                                 : out   std_logic_vector(1 downto 0);
          W_out_i_0                                 : out   std_logic_vector(2 to 2);
          msg_bitlen                                : in    std_logic_vector(63 downto 3) := (others => 'U');
          state_2                                   : in    std_logic := 'U';
          state_0                                   : in    std_logic := 'U';
          state_3                                   : in    std_logic := 'U';
          Kt_addr_5                                 : in    std_logic := 'U';
          Kt_addr_0                                 : in    std_logic := 'U';
          W_out_2_0_0_1                             : out   std_logic;
          W_out_2_0_0_0                             : out   std_logic;
          W_out_2_0_0_3                             : out   std_logic;
          W_out_2_0_1_8                             : out   std_logic;
          W_out_2_0_1_0                             : out   std_logic;
          W_out_2_i_0_18                            : out   std_logic;
          W_out_2_i_0_21                            : out   std_logic;
          W_out_2_i_0_17                            : out   std_logic;
          W_out_2_i_0_22                            : out   std_logic;
          W_out_2_i_0_20                            : out   std_logic;
          W_out_2_i_0_16                            : out   std_logic;
          W_out_2_i_0_19                            : out   std_logic;
          W_out_2_0_2_0                             : out   std_logic;
          W_out_2_0_2_8                             : out   std_logic;
          sha256_controller_0_di_o_3                : in    std_logic := 'U';
          sha256_controller_0_di_o_5                : in    std_logic := 'U';
          sha256_controller_0_di_o_0                : in    std_logic := 'U';
          W_out_2_i_1_18                            : out   std_logic;
          W_out_2_i_1_21                            : out   std_logic;
          W_out_2_i_1_17                            : out   std_logic;
          W_out_2_i_1_22                            : out   std_logic;
          W_out_2_i_1_20                            : out   std_logic;
          W_out_2_i_1_16                            : out   std_logic;
          W_out_2_i_1_19                            : out   std_logic;
          W_out_2_i_1_12                            : out   std_logic;
          W_out_2_i_1_8                             : out   std_logic;
          W_out_2_i_1_10                            : out   std_logic;
          W_out_2_i_1_13                            : out   std_logic;
          W_out_2_i_1_14                            : out   std_logic;
          W_out_2_i_1_11                            : out   std_logic;
          W_out_2_i_1_9                             : out   std_logic;
          W_out_2_i_1_1                             : out   std_logic;
          W_out_2_i_1_2                             : out   std_logic;
          W_out_2_i_1_0                             : out   std_logic;
          W_out_2_i_1_4                             : out   std_logic;
          W_out_2_i_1_3                             : out   std_logic;
          W_out_2_i_1_6                             : out   std_logic;
          W_out_2_i_1_5                             : out   std_logic;
          N_223                                     : in    std_logic := 'U';
          N_1702                                    : in    std_logic := 'U';
          N_1710                                    : in    std_logic := 'U';
          SHA256_Module_0_di_req_o                  : in    std_logic := 'U';
          N_388                                     : out   std_logic;
          N_112                                     : in    std_logic := 'U';
          one_insert                                : in    std_logic := 'U';
          Kt_addr_0_rep2                            : in    std_logic := 'U';
          sha_last_blk_reg                          : in    std_logic := 'U';
          Kt_addr_4_rep1                            : in    std_logic := 'U';
          bytes_sel                                 : in    std_logic := 'U';
          ren_pos                                   : in    std_logic := 'U';
          N_102                                     : in    std_logic := 'U';
          sha_last_blk_next_0_o2_2_out_0            : in    std_logic := 'U';
          N_361                                     : in    std_logic := 'U';
          SHA256_Module_0_data_available_lastbank_8 : in    std_logic := 'U';
          N_111                                     : in    std_logic := 'U';
          N_1690                                    : in    std_logic := 'U';
          N_245                                     : out   std_logic;
          N_1691                                    : in    std_logic := 'U';
          N_248                                     : out   std_logic;
          N_1693                                    : in    std_logic := 'U';
          N_251                                     : out   std_logic;
          N_1692                                    : in    std_logic := 'U';
          N_349                                     : out   std_logic;
          N_1718                                    : in    std_logic := 'U';
          N_1694                                    : in    std_logic := 'U';
          N_255                                     : out   std_logic;
          N_1698                                    : in    std_logic := 'U';
          N_1701                                    : in    std_logic := 'U';
          N_98                                      : out   std_logic;
          N_307                                     : out   std_logic;
          N_1696                                    : in    std_logic := 'U';
          N_1697                                    : in    std_logic := 'U';
          N_1695                                    : in    std_logic := 'U';
          N_1699                                    : in    std_logic := 'U';
          N_1707                                    : in    std_logic := 'U';
          N_1708                                    : in    std_logic := 'U';
          N_1709                                    : in    std_logic := 'U';
          N_1706                                    : in    std_logic := 'U';
          N_1704                                    : in    std_logic := 'U';
          N_1688                                    : in    std_logic := 'U';
          N_1687                                    : in    std_logic := 'U';
          N_1689                                    : in    std_logic := 'U';
          N_1713                                    : in    std_logic := 'U';
          N_1716                                    : in    std_logic := 'U';
          N_1712                                    : in    std_logic := 'U';
          N_1717                                    : in    std_logic := 'U';
          N_1715                                    : in    std_logic := 'U';
          N_1711                                    : in    std_logic := 'U';
          N_1714                                    : in    std_logic := 'U';
          N_273                                     : out   std_logic;
          N_266                                     : out   std_logic;
          N_263                                     : out   std_logic;
          N_260                                     : out   std_logic;
          N_287                                     : out   std_logic;
          N_290                                     : out   std_logic;
          N_293                                     : out   std_logic;
          N_296                                     : out   std_logic;
          N_299                                     : out   std_logic;
          N_302                                     : out   std_logic;
          N_305                                     : out   std_logic;
          N_268                                     : out   std_logic;
          N_275                                     : out   std_logic;
          N_278                                     : out   std_logic
        );
  end component;

  component sha256_msg_sch
    port( Wt_data                              : out   std_logic_vector(31 downto 0);
          W_out_2_0                            : in    std_logic_vector(5 to 5) := (others => 'U');
          W_out_i_i_2                          : in    std_logic_vector(31 to 31) := (others => 'U');
          W_out_i_i_1                          : in    std_logic_vector(31 to 31) := (others => 'U');
          W_out_2_i_0                          : in    std_logic_vector(30 downto 24) := (others => 'U');
          W_out_i_0                            : in    std_logic_vector(2 to 2) := (others => 'U');
          W_out_i_1                            : in    std_logic_vector(1 downto 0) := (others => 'U');
          W_out_2_0_0_3                        : in    std_logic := 'U';
          W_out_2_0_0_1                        : in    std_logic := 'U';
          W_out_2_0_0_0                        : in    std_logic := 'U';
          W_out_2_0_2_8                        : in    std_logic := 'U';
          W_out_2_0_2_0                        : in    std_logic := 'U';
          W_out_2_0_1_0                        : in    std_logic := 'U';
          W_out_2_0_1_8                        : in    std_logic := 'U';
          W_out_2_i_1_22                       : in    std_logic := 'U';
          W_out_2_i_1_21                       : in    std_logic := 'U';
          W_out_2_i_1_20                       : in    std_logic := 'U';
          W_out_2_i_1_19                       : in    std_logic := 'U';
          W_out_2_i_1_18                       : in    std_logic := 'U';
          W_out_2_i_1_17                       : in    std_logic := 'U';
          W_out_2_i_1_16                       : in    std_logic := 'U';
          W_out_2_i_1_14                       : in    std_logic := 'U';
          W_out_2_i_1_13                       : in    std_logic := 'U';
          W_out_2_i_1_12                       : in    std_logic := 'U';
          W_out_2_i_1_11                       : in    std_logic := 'U';
          W_out_2_i_1_10                       : in    std_logic := 'U';
          W_out_2_i_1_9                        : in    std_logic := 'U';
          W_out_2_i_1_8                        : in    std_logic := 'U';
          W_out_2_i_1_6                        : in    std_logic := 'U';
          W_out_2_i_1_5                        : in    std_logic := 'U';
          W_out_2_i_1_4                        : in    std_logic := 'U';
          W_out_2_i_1_3                        : in    std_logic := 'U';
          W_out_2_i_1_2                        : in    std_logic := 'U';
          W_out_2_i_1_1                        : in    std_logic := 'U';
          W_out_2_i_1_0                        : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          N_244_i_0                            : in    std_logic := 'U';
          next_r0_0_cry_0_Y                    : out   std_logic;
          N_251                                : in    std_logic := 'U';
          ld_i_i_3                             : in    std_logic := 'U';
          N_349                                : in    std_logic := 'U';
          N_248                                : in    std_logic := 'U';
          N_245                                : in    std_logic := 'U';
          N_255                                : in    std_logic := 'U';
          N_98                                 : in    std_logic := 'U';
          N_307                                : in    std_logic := 'U';
          N_305                                : in    std_logic := 'U';
          N_302                                : in    std_logic := 'U';
          N_299                                : in    std_logic := 'U';
          N_296                                : in    std_logic := 'U';
          N_293                                : in    std_logic := 'U';
          N_290                                : in    std_logic := 'U';
          N_287                                : in    std_logic := 'U';
          N_278                                : in    std_logic := 'U';
          N_275                                : in    std_logic := 'U';
          N_273                                : in    std_logic := 'U';
          N_268                                : in    std_logic := 'U';
          N_266                                : in    std_logic := 'U';
          N_263                                : in    std_logic := 'U';
          N_260                                : in    std_logic := 'U'
        );
  end component;

  component sha256_kt_rom
    port( hash_control_st_reg_ns_i_0_a2_0 : in    std_logic_vector(4 to 4) := (others => 'U');
          Kt_addr_fast                    : in    std_logic_vector(4 downto 0) := (others => 'U');
          hash_control_st_reg_ns_i_0_a2_2 : out   std_logic_vector(4 to 4);
          Kt_addr                         : in    std_logic_vector(5 downto 0) := (others => 'U');
          Kt_data_9                       : out   std_logic;
          Kt_data_0                       : out   std_logic;
          Kt_addr_3_rep1                  : in    std_logic := 'U';
          m62_am                          : out   std_logic;
          Kt_addr_0_rep1                  : in    std_logic := 'U';
          m104_bm                         : out   std_logic;
          Kt_addr_2_rep1                  : in    std_logic := 'U';
          Kt_addr_0_rep2                  : in    std_logic := 'U';
          m49_am                          : out   std_logic;
          Kt_addr_1_rep1                  : in    std_logic := 'U';
          m49_bm                          : out   std_logic;
          m137_am                         : out   std_logic;
          Kt_addr_3_rep2                  : in    std_logic := 'U';
          m137_bm                         : out   std_logic;
          Kt_addr_4_rep2                  : in    std_logic := 'U';
          m215_am                         : out   std_logic;
          Kt_addr_4_rep1                  : in    std_logic := 'U';
          m215_bm                         : out   std_logic;
          Kt_addr_2_rep2                  : in    std_logic := 'U';
          m250_am                         : out   std_logic;
          Kt_addr_1_rep2                  : in    std_logic := 'U';
          m250_bm                         : out   std_logic;
          m207_1_1                        : out   std_logic;
          m207_1_0                        : out   std_logic;
          m157                            : out   std_logic;
          m197_1_1                        : out   std_logic;
          m197_1_0                        : out   std_logic;
          m95_1_1                         : out   std_logic;
          m95_1_0                         : out   std_logic;
          m325                            : out   std_logic;
          m168_1_1                        : out   std_logic;
          m168_1_0                        : out   std_logic;
          m316                            : out   std_logic;
          m34                             : out   std_logic;
          m114                            : out   std_logic;
          m285                            : out   std_logic;
          m289                            : out   std_logic;
          m254                            : out   std_logic;
          m239                            : out   std_logic;
          m124                            : out   std_logic;
          m141                            : out   std_logic;
          m304                            : out   std_logic;
          m19                             : out   std_logic;
          pad_one_reg_0_0_a2_0            : in    std_logic := 'U';
          m296                            : out   std_logic;
          m78                             : out   std_logic;
          m219                            : out   std_logic;
          m230                            : out   std_logic;
          m177                            : out   std_logic;
          m73_0                           : out   std_logic;
          i3_mux_1                        : out   std_logic;
          m10_ns                          : out   std_logic;
          m67_ns                          : out   std_logic;
          m83_ns                          : out   std_logic;
          m110_ns                         : out   std_logic;
          m119_ns                         : out   std_logic;
          m144_ns                         : out   std_logic;
          m172_ns                         : out   std_logic;
          m222_ns                         : out   std_logic;
          m226_ns                         : out   std_logic;
          m235_ns                         : out   std_logic;
          m258_ns                         : out   std_logic;
          m276_ns                         : out   std_logic;
          m281_ns                         : out   std_logic;
          m292_ns                         : out   std_logic;
          m300_ns                         : out   std_logic;
          sha_last_blk_next_0_a4_0        : out   std_logic;
          m273                            : out   std_logic;
          m104_am                         : out   std_logic;
          m62_bm                          : out   std_logic
        );
  end component;

    signal \hash_control_st_reg_i[6]\, \msg_bitlen[3]\, 
        \msg_bitlen[4]\, \msg_bitlen[5]\, \msg_bitlen[6]\, 
        \msg_bitlen[7]\, \msg_bitlen[8]\, \msg_bitlen[9]\, 
        \msg_bitlen[10]\, \msg_bitlen[11]\, \msg_bitlen[12]\, 
        \msg_bitlen[13]\, \msg_bitlen[14]\, \msg_bitlen[15]\, 
        \msg_bitlen[16]\, \msg_bitlen[17]\, \msg_bitlen[18]\, 
        \msg_bitlen[19]\, \msg_bitlen[20]\, \msg_bitlen[21]\, 
        \msg_bitlen[22]\, \msg_bitlen[23]\, \msg_bitlen[24]\, 
        \msg_bitlen[25]\, \msg_bitlen[26]\, \msg_bitlen[27]\, 
        \msg_bitlen[28]\, \msg_bitlen[29]\, \msg_bitlen[30]\, 
        \msg_bitlen[31]\, \msg_bitlen[32]\, \msg_bitlen[33]\, 
        \msg_bitlen[34]\, \msg_bitlen[35]\, \msg_bitlen[36]\, 
        \msg_bitlen[37]\, \msg_bitlen[38]\, \msg_bitlen[39]\, 
        \msg_bitlen[40]\, \msg_bitlen[41]\, \msg_bitlen[42]\, 
        \msg_bitlen[43]\, \msg_bitlen[44]\, \msg_bitlen[45]\, 
        \msg_bitlen[46]\, \msg_bitlen[47]\, \msg_bitlen[48]\, 
        \msg_bitlen[49]\, \msg_bitlen[50]\, \msg_bitlen[51]\, 
        \msg_bitlen[52]\, \msg_bitlen[53]\, \msg_bitlen[54]\, 
        \msg_bitlen[55]\, \msg_bitlen[56]\, \msg_bitlen[57]\, 
        \msg_bitlen[58]\, \msg_bitlen[59]\, \msg_bitlen[60]\, 
        \msg_bitlen[61]\, \msg_bitlen[62]\, \msg_bitlen[63]\, 
        \Kt_addr[0]\, \Kt_addr[1]\, \Kt_addr[2]\, \Kt_addr[3]\, 
        \Kt_addr[4]\, \Kt_addr[5]\, \hash_control_st_reg[2]\, 
        \Kt_addr_fast[0]\, \Kt_addr_fast[1]\, \Kt_addr_fast[2]\, 
        \Kt_addr_fast[3]\, \Kt_addr_fast[4]\, 
        \hash_control_st_reg_ns_i_0_a2_0[4]\, 
        \hash_control_st_reg_ns_i_0_a2_2[4]\, one_insert, 
        sha_last_blk_reg, \SHA256_Module_0_di_req_o\, 
        Kt_addr_1_rep1, Kt_addr_1_rep2, Kt_addr_2_rep1, 
        Kt_addr_2_rep2, Kt_addr_0_rep1, Kt_addr_0_rep2, 
        Kt_addr_4_rep1, Kt_addr_4_rep2, Kt_addr_3_rep1, 
        Kt_addr_3_rep2, N_112, N_223, N_361, N_102, N_168_i_0, 
        pad_one_reg_0_0_a2_0, oregs_ce_i_a2_0_a2, 
        sha_last_blk_next_0_o2_2_out_0, sha_last_blk_next_0_a4_0, 
        N_388, N_111, core_ce_o_iv_i_0, N_244_i_0, ld_i_i_3, 
        \W_out_2_0[5]\, \W_out_2_0_0[4]\, \W_out_2_0_0[3]\, 
        \W_out_2_0_0[6]\, \W_out_i_i_2[31]\, \W_out_i_i_1[31]\, 
        \W_out_2_0_1[15]\, \W_out_2_0_1[7]\, \W_out_i_1[0]\, 
        \W_out_i_1[1]\, \W_out_i_0[2]\, \W_out_2_i_0[26]\, 
        \W_out_2_i_0[29]\, \W_out_2_i_0[25]\, \W_out_2_i_0[30]\, 
        \W_out_2_i_0[28]\, \W_out_2_i_0[24]\, \W_out_2_i_0[27]\, 
        \W_out_2_0_2[15]\, \W_out_2_0_2[23]\, \W_out_2_i_1[26]\, 
        \W_out_2_i_1[29]\, \W_out_2_i_1[25]\, \W_out_2_i_1[30]\, 
        \W_out_2_i_1[28]\, \W_out_2_i_1[24]\, \W_out_2_i_1[27]\, 
        \W_out_2_i_1[20]\, \W_out_2_i_1[16]\, \W_out_2_i_1[18]\, 
        \W_out_2_i_1[21]\, \W_out_2_i_1[22]\, \W_out_2_i_1[19]\, 
        \W_out_2_i_1[17]\, \W_out_2_i_1[9]\, \W_out_2_i_1[10]\, 
        \W_out_2_i_1[8]\, \W_out_2_i_1[12]\, \W_out_2_i_1[11]\, 
        \W_out_2_i_1[14]\, \W_out_2_i_1[13]\, N_245, N_248, N_251, 
        N_349, N_255, N_98, N_307, N_273, N_266, N_263, N_260, 
        N_287, N_290, N_293, N_296, N_299, N_302, N_305, N_268, 
        N_275, N_278, \Wt_data[0]\, \Wt_data[1]\, \Wt_data[2]\, 
        \Wt_data[3]\, \Wt_data[4]\, \Wt_data[5]\, \Wt_data[6]\, 
        \Wt_data[7]\, \Wt_data[8]\, \Wt_data[9]\, \Wt_data[10]\, 
        \Wt_data[11]\, \Wt_data[12]\, \Wt_data[13]\, 
        \Wt_data[14]\, \Wt_data[15]\, \Wt_data[16]\, 
        \Wt_data[17]\, \Wt_data[18]\, \Wt_data[19]\, 
        \Wt_data[20]\, \Wt_data[21]\, \Wt_data[22]\, 
        \Wt_data[23]\, \Wt_data[24]\, \Wt_data[25]\, 
        \Wt_data[26]\, \Wt_data[27]\, \Wt_data[28]\, 
        \Wt_data[29]\, \Wt_data[30]\, \Wt_data[31]\, 
        next_r0_0_cry_0_Y, \R1_data[0]\, \R1_data[1]\, 
        \R1_data[2]\, \R1_data[3]\, \R1_data[4]\, \R1_data[5]\, 
        \R1_data[6]\, \R1_data[7]\, \R1_data[8]\, \R1_data[9]\, 
        \R1_data[10]\, \R1_data[11]\, \R1_data[12]\, 
        \R1_data[13]\, \R1_data[14]\, \R1_data[15]\, 
        \R1_data[16]\, \R1_data[17]\, \R1_data[18]\, 
        \R1_data[19]\, \R1_data[20]\, \R1_data[21]\, 
        \R1_data[22]\, \R1_data[23]\, \R1_data[24]\, 
        \R1_data[25]\, \R1_data[26]\, \R1_data[27]\, 
        \R1_data[28]\, \R1_data[29]\, \R1_data[30]\, 
        \R1_data[31]\, \R2_data[0]\, \R2_data[1]\, \R2_data[2]\, 
        \R2_data[3]\, \R2_data[4]\, \R2_data[5]\, \R2_data[6]\, 
        \R2_data[7]\, \R2_data[8]\, \R2_data[9]\, \R2_data[10]\, 
        \R2_data[11]\, \R2_data[12]\, \R2_data[13]\, 
        \R2_data[14]\, \R2_data[15]\, \R2_data[16]\, 
        \R2_data[17]\, \R2_data[18]\, \R2_data[19]\, 
        \R2_data[20]\, \R2_data[21]\, \R2_data[22]\, 
        \R2_data[23]\, \R2_data[24]\, \R2_data[25]\, 
        \R2_data[26]\, \R2_data[27]\, \R2_data[28]\, 
        \R2_data[29]\, \R2_data[30]\, \R2_data[31]\, \R3_data[0]\, 
        \R3_data[1]\, \R3_data[2]\, \R3_data[3]\, \R3_data[4]\, 
        \R3_data[5]\, \R3_data[6]\, \R3_data[7]\, \R3_data[8]\, 
        \R3_data[9]\, \R3_data[10]\, \R3_data[11]\, \R3_data[12]\, 
        \R3_data[13]\, \R3_data[14]\, \R3_data[15]\, 
        \R3_data[16]\, \R3_data[17]\, \R3_data[18]\, 
        \R3_data[19]\, \R3_data[20]\, \R3_data[21]\, 
        \R3_data[22]\, \R3_data[23]\, \R3_data[24]\, 
        \R3_data[25]\, \R3_data[26]\, \R3_data[27]\, 
        \R3_data[28]\, \R3_data[29]\, \R3_data[30]\, 
        \R3_data[31]\, \R5_data[0]\, \R5_data[1]\, \R5_data[2]\, 
        \R5_data[3]\, \R5_data[4]\, \R5_data[5]\, \R5_data[6]\, 
        \R5_data[7]\, \R5_data[8]\, \R5_data[9]\, \R5_data[10]\, 
        \R5_data[11]\, \R5_data[12]\, \R5_data[13]\, 
        \R5_data[14]\, \R5_data[15]\, \R5_data[16]\, 
        \R5_data[17]\, \R5_data[18]\, \R5_data[19]\, 
        \R5_data[20]\, \R5_data[21]\, \R5_data[22]\, 
        \R5_data[23]\, \R5_data[24]\, \R5_data[25]\, 
        \R5_data[26]\, \R5_data[27]\, \R5_data[28]\, 
        \R5_data[29]\, \R5_data[30]\, \R5_data[31]\, \R6_data[0]\, 
        \R6_data[1]\, \R6_data[2]\, \R6_data[3]\, \R6_data[4]\, 
        \R6_data[5]\, \R6_data[6]\, \R6_data[7]\, \R6_data[8]\, 
        \R6_data[9]\, \R6_data[10]\, \R6_data[11]\, \R6_data[12]\, 
        \R6_data[13]\, \R6_data[14]\, \R6_data[15]\, 
        \R6_data[16]\, \R6_data[17]\, \R6_data[18]\, 
        \R6_data[19]\, \R6_data[20]\, \R6_data[21]\, 
        \R6_data[22]\, \R6_data[23]\, \R6_data[24]\, 
        \R6_data[25]\, \R6_data[26]\, \R6_data[27]\, 
        \R6_data[28]\, \R6_data[29]\, \R6_data[30]\, 
        \R6_data[31]\, \R7_data[0]\, \R7_data[1]\, \R7_data[2]\, 
        \R7_data[3]\, \R7_data[4]\, \R7_data[5]\, \R7_data[6]\, 
        \R7_data[7]\, \R7_data[8]\, \R7_data[9]\, \R7_data[10]\, 
        \R7_data[11]\, \R7_data[12]\, \R7_data[13]\, 
        \R7_data[14]\, \R7_data[15]\, \R7_data[16]\, 
        \R7_data[17]\, \R7_data[18]\, \R7_data[19]\, 
        \R7_data[20]\, \R7_data[21]\, \R7_data[22]\, 
        \R7_data[23]\, \R7_data[24]\, \R7_data[25]\, 
        \R7_data[26]\, \R7_data[27]\, \R7_data[28]\, 
        \R7_data[29]\, \R7_data[30]\, \R7_data[31]\, \R0_data[0]\, 
        \R0_data[1]\, \R0_data[2]\, \R0_data[3]\, \R0_data[4]\, 
        \R0_data[5]\, \R0_data[6]\, \R0_data[7]\, \R0_data[8]\, 
        \R0_data[9]\, \R0_data[10]\, \R0_data[11]\, \R0_data[12]\, 
        \R0_data[13]\, \R0_data[14]\, \R0_data[15]\, 
        \R0_data[16]\, \R0_data[17]\, \R0_data[18]\, 
        \R0_data[19]\, \R0_data[20]\, \R0_data[21]\, 
        \R0_data[22]\, \R0_data[23]\, \R0_data[24]\, 
        \R0_data[25]\, \R0_data[26]\, \R0_data[27]\, 
        \R0_data[28]\, \R0_data[29]\, \R0_data[30]\, 
        \R0_data[31]\, \R4_data[0]\, \R4_data[1]\, \R4_data[2]\, 
        \R4_data[3]\, \R4_data[4]\, \R4_data[5]\, \R4_data[6]\, 
        \R4_data[7]\, \R4_data[8]\, \R4_data[9]\, \R4_data[10]\, 
        \R4_data[11]\, \R4_data[12]\, \R4_data[13]\, 
        \R4_data[14]\, \R4_data[15]\, \R4_data[16]\, 
        \R4_data[17]\, \R4_data[18]\, \R4_data[19]\, 
        \R4_data[20]\, \R4_data[21]\, \R4_data[22]\, 
        \R4_data[23]\, \R4_data[24]\, \R4_data[25]\, 
        \R4_data[26]\, \R4_data[27]\, \R4_data[28]\, 
        \R4_data[29]\, \R4_data[30]\, \R4_data[31]\, \N4_data[1]\, 
        \N4_data[2]\, \N4_data[3]\, \N4_data[4]\, \N4_data[5]\, 
        \N4_data[6]\, \N4_data[7]\, \N4_data[8]\, \N4_data[9]\, 
        \N4_data[10]\, \N4_data[11]\, \N4_data[12]\, 
        \N4_data[13]\, \N4_data[14]\, \N4_data[15]\, 
        \N4_data[16]\, \N4_data[17]\, \N4_data[18]\, 
        \N4_data[19]\, \N4_data[20]\, \N4_data[21]\, 
        \N4_data[22]\, \N4_data[23]\, \N4_data[24]\, 
        \N4_data[25]\, \N4_data[26]\, \N4_data[27]\, 
        \N4_data[28]\, \N4_data[29]\, \N4_data[30]\, 
        \N4_data[31]\, \N0_data[1]\, \N0_data[2]\, \N0_data[3]\, 
        \N0_data[4]\, \N0_data[5]\, \N0_data[6]\, \N0_data[7]\, 
        \N0_data[8]\, \N0_data[9]\, \N0_data[10]\, \N0_data[11]\, 
        \N0_data[12]\, \N0_data[13]\, \N0_data[14]\, 
        \N0_data[15]\, \N0_data[16]\, \N0_data[17]\, 
        \N0_data[18]\, \N0_data[19]\, \N0_data[20]\, 
        \N0_data[21]\, \N0_data[22]\, \N0_data[23]\, 
        \N0_data[24]\, \N0_data[25]\, \N0_data[26]\, 
        \N0_data[27]\, \N0_data[28]\, \N0_data[29]\, 
        \N0_data[30]\, \N0_data[31]\, \Kt_data[15]\, 
        \Kt_data[24]\, \N3_data[1]\, \N3_data[2]\, \N3_data[3]\, 
        \N3_data[4]\, \N3_data[5]\, \N3_data[6]\, \N3_data[7]\, 
        \N3_data[8]\, \N3_data[9]\, \N3_data[10]\, \N3_data[11]\, 
        \N3_data[12]\, \N3_data[13]\, \N3_data[14]\, 
        \N3_data[15]\, \N3_data[16]\, \N3_data[17]\, 
        \N3_data[18]\, \N3_data[19]\, \N3_data[20]\, 
        \N3_data[21]\, \N3_data[22]\, \N3_data[23]\, 
        \N3_data[24]\, \N3_data[25]\, \N3_data[26]\, 
        \N3_data[27]\, \N3_data[28]\, \N3_data[29]\, 
        \N3_data[30]\, \N3_data[31]\, \N2_data[1]\, \N2_data[2]\, 
        \N2_data[3]\, \N2_data[4]\, \N2_data[5]\, \N2_data[6]\, 
        \N2_data[7]\, \N2_data[8]\, \N2_data[9]\, \N2_data[10]\, 
        \N2_data[11]\, \N2_data[12]\, \N2_data[13]\, 
        \N2_data[14]\, \N2_data[15]\, \N2_data[16]\, 
        \N2_data[17]\, \N2_data[18]\, \N2_data[19]\, 
        \N2_data[20]\, \N2_data[21]\, \N2_data[22]\, 
        \N2_data[23]\, \N2_data[24]\, \N2_data[25]\, 
        \N2_data[26]\, \N2_data[27]\, \N2_data[28]\, 
        \N2_data[29]\, \N2_data[30]\, \N2_data[31]\, \N1_data[1]\, 
        \N1_data[2]\, \N1_data[3]\, \N1_data[4]\, \N1_data[5]\, 
        \N1_data[6]\, \N1_data[7]\, \N1_data[8]\, \N1_data[9]\, 
        \N1_data[10]\, \N1_data[11]\, \N1_data[12]\, 
        \N1_data[13]\, \N1_data[14]\, \N1_data[15]\, 
        \N1_data[16]\, \N1_data[17]\, \N1_data[18]\, 
        \N1_data[19]\, \N1_data[20]\, \N1_data[21]\, 
        \N1_data[22]\, \N1_data[23]\, \N1_data[24]\, 
        \N1_data[25]\, \N1_data[26]\, \N1_data[27]\, 
        \N1_data[28]\, \N1_data[29]\, \N1_data[30]\, 
        \N1_data[31]\, \N7_data[1]\, \N7_data[2]\, \N7_data[3]\, 
        \N7_data[4]\, \N7_data[5]\, \N7_data[6]\, \N7_data[7]\, 
        \N7_data[8]\, \N7_data[9]\, \N7_data[10]\, \N7_data[11]\, 
        \N7_data[12]\, \N7_data[13]\, \N7_data[14]\, 
        \N7_data[15]\, \N7_data[16]\, \N7_data[17]\, 
        \N7_data[18]\, \N7_data[19]\, \N7_data[20]\, 
        \N7_data[21]\, \N7_data[22]\, \N7_data[23]\, 
        \N7_data[24]\, \N7_data[25]\, \N7_data[26]\, 
        \N7_data[27]\, \N7_data[28]\, \N7_data[29]\, 
        \N7_data[30]\, \N7_data[31]\, \N6_data[1]\, \N6_data[2]\, 
        \N6_data[3]\, \N6_data[4]\, \N6_data[5]\, \N6_data[6]\, 
        \N6_data[7]\, \N6_data[8]\, \N6_data[9]\, \N6_data[10]\, 
        \N6_data[11]\, \N6_data[12]\, \N6_data[13]\, 
        \N6_data[14]\, \N6_data[15]\, \N6_data[16]\, 
        \N6_data[17]\, \N6_data[18]\, \N6_data[19]\, 
        \N6_data[20]\, \N6_data[21]\, \N6_data[22]\, 
        \N6_data[23]\, \N6_data[24]\, \N6_data[25]\, 
        \N6_data[26]\, \N6_data[27]\, \N6_data[28]\, 
        \N6_data[29]\, \N6_data[30]\, \N6_data[31]\, \N5_data[1]\, 
        \N5_data[2]\, \N5_data[3]\, \N5_data[4]\, \N5_data[5]\, 
        \N5_data[6]\, \N5_data[7]\, \N5_data[8]\, \N5_data[9]\, 
        \N5_data[10]\, \N5_data[11]\, \N5_data[12]\, 
        \N5_data[13]\, \N5_data[14]\, \N5_data[15]\, 
        \N5_data[16]\, \N5_data[17]\, \N5_data[18]\, 
        \N5_data[19]\, \N5_data[20]\, \N5_data[21]\, 
        \N5_data[22]\, \N5_data[23]\, \N5_data[24]\, 
        \N5_data[25]\, \N5_data[26]\, \N5_data[27]\, 
        \N5_data[28]\, \N5_data[29]\, \N5_data[30]\, 
        \N5_data[31]\, next_reg_H4_cry_0_0_Y, 
        next_reg_H0_cry_0_0_Y, m34, m49_am, m49_bm, m62_am, 
        m62_bm, m67_ns, m73, m78, m83_ns, m95_1_0, m95_1_1, 
        m104_am, m104_bm, m110_ns, m114, m119_ns, m124, m137_am, 
        m137_bm, m141, m144_ns, m157, m168_1_0, m168_1_1, m172_ns, 
        m177, m197_1_0, m197_1_1, m207_1_0, m207_1_1, m215_am, 
        m215_bm, m219, m222_ns, m226_ns, m230, m235_ns, m239, 
        m250_am, m250_bm, m254, m258_ns, m273, m276_ns, m281_ns, 
        m285, m289, m292_ns, m296, m300_ns, m304, i3_mux_1, m325, 
        m316, next_reg_H3_cry_0_0_Y, next_reg_H2_cry_0_0_Y, 
        next_reg_H1_cry_0_0_Y, next_reg_H7_cry_0_0_Y, 
        next_reg_H6_cry_0_0_Y, next_reg_H5_cry_0_0_Y, m10_ns, m19, 
        GND_net_1, VCC_net_1 : std_logic;

    for all : sha256_control
	Use entity work.sha256_control(DEF_ARCH);
    for all : sha256_hash_core
	Use entity work.sha256_hash_core(DEF_ARCH);
    for all : sha256_regs
	Use entity work.sha256_regs(DEF_ARCH);
    for all : sha256_padding
	Use entity work.sha256_padding(DEF_ARCH);
    for all : sha256_msg_sch
	Use entity work.sha256_msg_sch(DEF_ARCH);
    for all : sha256_kt_rom
	Use entity work.sha256_kt_rom(DEF_ARCH);
begin 

    SHA256_Module_0_di_req_o <= \SHA256_Module_0_di_req_o\;

    Inst_sha256_control : sha256_control
      port map(hash_control_st_reg_i(6) => 
        \hash_control_st_reg_i[6]\, msg_bitlen(63) => 
        \msg_bitlen[63]\, msg_bitlen(62) => \msg_bitlen[62]\, 
        msg_bitlen(61) => \msg_bitlen[61]\, msg_bitlen(60) => 
        \msg_bitlen[60]\, msg_bitlen(59) => \msg_bitlen[59]\, 
        msg_bitlen(58) => \msg_bitlen[58]\, msg_bitlen(57) => 
        \msg_bitlen[57]\, msg_bitlen(56) => \msg_bitlen[56]\, 
        msg_bitlen(55) => \msg_bitlen[55]\, msg_bitlen(54) => 
        \msg_bitlen[54]\, msg_bitlen(53) => \msg_bitlen[53]\, 
        msg_bitlen(52) => \msg_bitlen[52]\, msg_bitlen(51) => 
        \msg_bitlen[51]\, msg_bitlen(50) => \msg_bitlen[50]\, 
        msg_bitlen(49) => \msg_bitlen[49]\, msg_bitlen(48) => 
        \msg_bitlen[48]\, msg_bitlen(47) => \msg_bitlen[47]\, 
        msg_bitlen(46) => \msg_bitlen[46]\, msg_bitlen(45) => 
        \msg_bitlen[45]\, msg_bitlen(44) => \msg_bitlen[44]\, 
        msg_bitlen(43) => \msg_bitlen[43]\, msg_bitlen(42) => 
        \msg_bitlen[42]\, msg_bitlen(41) => \msg_bitlen[41]\, 
        msg_bitlen(40) => \msg_bitlen[40]\, msg_bitlen(39) => 
        \msg_bitlen[39]\, msg_bitlen(38) => \msg_bitlen[38]\, 
        msg_bitlen(37) => \msg_bitlen[37]\, msg_bitlen(36) => 
        \msg_bitlen[36]\, msg_bitlen(35) => \msg_bitlen[35]\, 
        msg_bitlen(34) => \msg_bitlen[34]\, msg_bitlen(33) => 
        \msg_bitlen[33]\, msg_bitlen(32) => \msg_bitlen[32]\, 
        msg_bitlen(31) => \msg_bitlen[31]\, msg_bitlen(30) => 
        \msg_bitlen[30]\, msg_bitlen(29) => \msg_bitlen[29]\, 
        msg_bitlen(28) => \msg_bitlen[28]\, msg_bitlen(27) => 
        \msg_bitlen[27]\, msg_bitlen(26) => \msg_bitlen[26]\, 
        msg_bitlen(25) => \msg_bitlen[25]\, msg_bitlen(24) => 
        \msg_bitlen[24]\, msg_bitlen(23) => \msg_bitlen[23]\, 
        msg_bitlen(22) => \msg_bitlen[22]\, msg_bitlen(21) => 
        \msg_bitlen[21]\, msg_bitlen(20) => \msg_bitlen[20]\, 
        msg_bitlen(19) => \msg_bitlen[19]\, msg_bitlen(18) => 
        \msg_bitlen[18]\, msg_bitlen(17) => \msg_bitlen[17]\, 
        msg_bitlen(16) => \msg_bitlen[16]\, msg_bitlen(15) => 
        \msg_bitlen[15]\, msg_bitlen(14) => \msg_bitlen[14]\, 
        msg_bitlen(13) => \msg_bitlen[13]\, msg_bitlen(12) => 
        \msg_bitlen[12]\, msg_bitlen(11) => \msg_bitlen[11]\, 
        msg_bitlen(10) => \msg_bitlen[10]\, msg_bitlen(9) => 
        \msg_bitlen[9]\, msg_bitlen(8) => \msg_bitlen[8]\, 
        msg_bitlen(7) => \msg_bitlen[7]\, msg_bitlen(6) => 
        \msg_bitlen[6]\, msg_bitlen(5) => \msg_bitlen[5]\, 
        msg_bitlen(4) => \msg_bitlen[4]\, msg_bitlen(3) => 
        \msg_bitlen[3]\, Kt_addr(5) => \Kt_addr[5]\, Kt_addr(4)
         => \Kt_addr[4]\, Kt_addr(3) => \Kt_addr[3]\, Kt_addr(2)
         => \Kt_addr[2]\, Kt_addr(1) => \Kt_addr[1]\, Kt_addr(0)
         => \Kt_addr[0]\, Kt_addr_fast(4) => \Kt_addr_fast[4]\, 
        Kt_addr_fast(3) => \Kt_addr_fast[3]\, Kt_addr_fast(2) => 
        \Kt_addr_fast[2]\, Kt_addr_fast(1) => \Kt_addr_fast[1]\, 
        Kt_addr_fast(0) => \Kt_addr_fast[0]\, state(1) => state_0, 
        hash_control_st_reg_ns_i_0_a2_0(4) => 
        \hash_control_st_reg_ns_i_0_a2_0[4]\, 
        reg_17x32_0_valid_bytes_0(1) => 
        reg_17x32_0_valid_bytes_0(1), 
        reg_17x32_0_valid_bytes_0(0) => 
        reg_17x32_0_valid_bytes_0(0), 
        hash_control_st_reg_ns_i_0_a2_2(4) => 
        \hash_control_st_reg_ns_i_0_a2_2[4]\, 
        hash_control_st_reg_2 => \hash_control_st_reg[2]\, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, one_insert => 
        one_insert, sha_last_blk_reg => sha_last_blk_reg, 
        SHA256_Module_0_di_req_o => \SHA256_Module_0_di_req_o\, 
        SHA256_BLOCK_0_do_valid_o => SHA256_BLOCK_0_do_valid_o, 
        Kt_addr_1_rep1 => Kt_addr_1_rep1, Kt_addr_1_rep2 => 
        Kt_addr_1_rep2, Kt_addr_2_rep1 => Kt_addr_2_rep1, 
        Kt_addr_2_rep2 => Kt_addr_2_rep2, Kt_addr_0_rep1 => 
        Kt_addr_0_rep1, Kt_addr_0_rep2 => Kt_addr_0_rep2, 
        Kt_addr_4_rep1 => Kt_addr_4_rep1, Kt_addr_4_rep2 => 
        Kt_addr_4_rep2, Kt_addr_3_rep1 => Kt_addr_3_rep1, 
        Kt_addr_3_rep2 => Kt_addr_3_rep2, N_112 => N_112, 
        SHA256_Module_0_waiting_data => 
        SHA256_Module_0_waiting_data, N_223 => N_223, N_361 => 
        N_361, N_102 => N_102, 
        SHA256_Module_0_data_available_lastbank_8 => 
        SHA256_Module_0_data_available_lastbank_8, N_168_i_0 => 
        N_168_i_0, pad_one_reg_0_0_a2_0 => pad_one_reg_0_0_a2_0, 
        oregs_ce_i_a2_0_a2 => oregs_ce_i_a2_0_a2, 
        sha_last_blk_next_0_o2_2_out_0 => 
        sha_last_blk_next_0_o2_2_out_0, N_484 => N_484, bytes_sel
         => bytes_sel, sha_last_blk_next_0_a4_0 => 
        sha_last_blk_next_0_a4_0, N_388 => N_388, N_111 => N_111, 
        core_ce_o_iv_i_0 => core_ce_o_iv_i_0, N_244_i_0 => 
        N_244_i_0, SHA256_Module_0_error_o => 
        SHA256_Module_0_error_o, ld_i_i_3 => ld_i_i_3, 
        SHA256_BLOCK_0_start_o => SHA256_BLOCK_0_start_o);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    Inst_sha256_hash_core : sha256_hash_core
      port map(R1_data(31) => \R1_data[31]\, R1_data(30) => 
        \R1_data[30]\, R1_data(29) => \R1_data[29]\, R1_data(28)
         => \R1_data[28]\, R1_data(27) => \R1_data[27]\, 
        R1_data(26) => \R1_data[26]\, R1_data(25) => 
        \R1_data[25]\, R1_data(24) => \R1_data[24]\, R1_data(23)
         => \R1_data[23]\, R1_data(22) => \R1_data[22]\, 
        R1_data(21) => \R1_data[21]\, R1_data(20) => 
        \R1_data[20]\, R1_data(19) => \R1_data[19]\, R1_data(18)
         => \R1_data[18]\, R1_data(17) => \R1_data[17]\, 
        R1_data(16) => \R1_data[16]\, R1_data(15) => 
        \R1_data[15]\, R1_data(14) => \R1_data[14]\, R1_data(13)
         => \R1_data[13]\, R1_data(12) => \R1_data[12]\, 
        R1_data(11) => \R1_data[11]\, R1_data(10) => 
        \R1_data[10]\, R1_data(9) => \R1_data[9]\, R1_data(8) => 
        \R1_data[8]\, R1_data(7) => \R1_data[7]\, R1_data(6) => 
        \R1_data[6]\, R1_data(5) => \R1_data[5]\, R1_data(4) => 
        \R1_data[4]\, R1_data(3) => \R1_data[3]\, R1_data(2) => 
        \R1_data[2]\, R1_data(1) => \R1_data[1]\, R1_data(0) => 
        \R1_data[0]\, R2_data(31) => \R2_data[31]\, R2_data(30)
         => \R2_data[30]\, R2_data(29) => \R2_data[29]\, 
        R2_data(28) => \R2_data[28]\, R2_data(27) => 
        \R2_data[27]\, R2_data(26) => \R2_data[26]\, R2_data(25)
         => \R2_data[25]\, R2_data(24) => \R2_data[24]\, 
        R2_data(23) => \R2_data[23]\, R2_data(22) => 
        \R2_data[22]\, R2_data(21) => \R2_data[21]\, R2_data(20)
         => \R2_data[20]\, R2_data(19) => \R2_data[19]\, 
        R2_data(18) => \R2_data[18]\, R2_data(17) => 
        \R2_data[17]\, R2_data(16) => \R2_data[16]\, R2_data(15)
         => \R2_data[15]\, R2_data(14) => \R2_data[14]\, 
        R2_data(13) => \R2_data[13]\, R2_data(12) => 
        \R2_data[12]\, R2_data(11) => \R2_data[11]\, R2_data(10)
         => \R2_data[10]\, R2_data(9) => \R2_data[9]\, R2_data(8)
         => \R2_data[8]\, R2_data(7) => \R2_data[7]\, R2_data(6)
         => \R2_data[6]\, R2_data(5) => \R2_data[5]\, R2_data(4)
         => \R2_data[4]\, R2_data(3) => \R2_data[3]\, R2_data(2)
         => \R2_data[2]\, R2_data(1) => \R2_data[1]\, R2_data(0)
         => \R2_data[0]\, R3_data(31) => \R3_data[31]\, 
        R3_data(30) => \R3_data[30]\, R3_data(29) => 
        \R3_data[29]\, R3_data(28) => \R3_data[28]\, R3_data(27)
         => \R3_data[27]\, R3_data(26) => \R3_data[26]\, 
        R3_data(25) => \R3_data[25]\, R3_data(24) => 
        \R3_data[24]\, R3_data(23) => \R3_data[23]\, R3_data(22)
         => \R3_data[22]\, R3_data(21) => \R3_data[21]\, 
        R3_data(20) => \R3_data[20]\, R3_data(19) => 
        \R3_data[19]\, R3_data(18) => \R3_data[18]\, R3_data(17)
         => \R3_data[17]\, R3_data(16) => \R3_data[16]\, 
        R3_data(15) => \R3_data[15]\, R3_data(14) => 
        \R3_data[14]\, R3_data(13) => \R3_data[13]\, R3_data(12)
         => \R3_data[12]\, R3_data(11) => \R3_data[11]\, 
        R3_data(10) => \R3_data[10]\, R3_data(9) => \R3_data[9]\, 
        R3_data(8) => \R3_data[8]\, R3_data(7) => \R3_data[7]\, 
        R3_data(6) => \R3_data[6]\, R3_data(5) => \R3_data[5]\, 
        R3_data(4) => \R3_data[4]\, R3_data(3) => \R3_data[3]\, 
        R3_data(2) => \R3_data[2]\, R3_data(1) => \R3_data[1]\, 
        R3_data(0) => \R3_data[0]\, R5_data(31) => \R5_data[31]\, 
        R5_data(30) => \R5_data[30]\, R5_data(29) => 
        \R5_data[29]\, R5_data(28) => \R5_data[28]\, R5_data(27)
         => \R5_data[27]\, R5_data(26) => \R5_data[26]\, 
        R5_data(25) => \R5_data[25]\, R5_data(24) => 
        \R5_data[24]\, R5_data(23) => \R5_data[23]\, R5_data(22)
         => \R5_data[22]\, R5_data(21) => \R5_data[21]\, 
        R5_data(20) => \R5_data[20]\, R5_data(19) => 
        \R5_data[19]\, R5_data(18) => \R5_data[18]\, R5_data(17)
         => \R5_data[17]\, R5_data(16) => \R5_data[16]\, 
        R5_data(15) => \R5_data[15]\, R5_data(14) => 
        \R5_data[14]\, R5_data(13) => \R5_data[13]\, R5_data(12)
         => \R5_data[12]\, R5_data(11) => \R5_data[11]\, 
        R5_data(10) => \R5_data[10]\, R5_data(9) => \R5_data[9]\, 
        R5_data(8) => \R5_data[8]\, R5_data(7) => \R5_data[7]\, 
        R5_data(6) => \R5_data[6]\, R5_data(5) => \R5_data[5]\, 
        R5_data(4) => \R5_data[4]\, R5_data(3) => \R5_data[3]\, 
        R5_data(2) => \R5_data[2]\, R5_data(1) => \R5_data[1]\, 
        R5_data(0) => \R5_data[0]\, R6_data(31) => \R6_data[31]\, 
        R6_data(30) => \R6_data[30]\, R6_data(29) => 
        \R6_data[29]\, R6_data(28) => \R6_data[28]\, R6_data(27)
         => \R6_data[27]\, R6_data(26) => \R6_data[26]\, 
        R6_data(25) => \R6_data[25]\, R6_data(24) => 
        \R6_data[24]\, R6_data(23) => \R6_data[23]\, R6_data(22)
         => \R6_data[22]\, R6_data(21) => \R6_data[21]\, 
        R6_data(20) => \R6_data[20]\, R6_data(19) => 
        \R6_data[19]\, R6_data(18) => \R6_data[18]\, R6_data(17)
         => \R6_data[17]\, R6_data(16) => \R6_data[16]\, 
        R6_data(15) => \R6_data[15]\, R6_data(14) => 
        \R6_data[14]\, R6_data(13) => \R6_data[13]\, R6_data(12)
         => \R6_data[12]\, R6_data(11) => \R6_data[11]\, 
        R6_data(10) => \R6_data[10]\, R6_data(9) => \R6_data[9]\, 
        R6_data(8) => \R6_data[8]\, R6_data(7) => \R6_data[7]\, 
        R6_data(6) => \R6_data[6]\, R6_data(5) => \R6_data[5]\, 
        R6_data(4) => \R6_data[4]\, R6_data(3) => \R6_data[3]\, 
        R6_data(2) => \R6_data[2]\, R6_data(1) => \R6_data[1]\, 
        R6_data(0) => \R6_data[0]\, R7_data(31) => \R7_data[31]\, 
        R7_data(30) => \R7_data[30]\, R7_data(29) => 
        \R7_data[29]\, R7_data(28) => \R7_data[28]\, R7_data(27)
         => \R7_data[27]\, R7_data(26) => \R7_data[26]\, 
        R7_data(25) => \R7_data[25]\, R7_data(24) => 
        \R7_data[24]\, R7_data(23) => \R7_data[23]\, R7_data(22)
         => \R7_data[22]\, R7_data(21) => \R7_data[21]\, 
        R7_data(20) => \R7_data[20]\, R7_data(19) => 
        \R7_data[19]\, R7_data(18) => \R7_data[18]\, R7_data(17)
         => \R7_data[17]\, R7_data(16) => \R7_data[16]\, 
        R7_data(15) => \R7_data[15]\, R7_data(14) => 
        \R7_data[14]\, R7_data(13) => \R7_data[13]\, R7_data(12)
         => \R7_data[12]\, R7_data(11) => \R7_data[11]\, 
        R7_data(10) => \R7_data[10]\, R7_data(9) => \R7_data[9]\, 
        R7_data(8) => \R7_data[8]\, R7_data(7) => \R7_data[7]\, 
        R7_data(6) => \R7_data[6]\, R7_data(5) => \R7_data[5]\, 
        R7_data(4) => \R7_data[4]\, R7_data(3) => \R7_data[3]\, 
        R7_data(2) => \R7_data[2]\, R7_data(1) => \R7_data[1]\, 
        R7_data(0) => \R7_data[0]\, R0_data(31) => \R0_data[31]\, 
        R0_data(30) => \R0_data[30]\, R0_data(29) => 
        \R0_data[29]\, R0_data(28) => \R0_data[28]\, R0_data(27)
         => \R0_data[27]\, R0_data(26) => \R0_data[26]\, 
        R0_data(25) => \R0_data[25]\, R0_data(24) => 
        \R0_data[24]\, R0_data(23) => \R0_data[23]\, R0_data(22)
         => \R0_data[22]\, R0_data(21) => \R0_data[21]\, 
        R0_data(20) => \R0_data[20]\, R0_data(19) => 
        \R0_data[19]\, R0_data(18) => \R0_data[18]\, R0_data(17)
         => \R0_data[17]\, R0_data(16) => \R0_data[16]\, 
        R0_data(15) => \R0_data[15]\, R0_data(14) => 
        \R0_data[14]\, R0_data(13) => \R0_data[13]\, R0_data(12)
         => \R0_data[12]\, R0_data(11) => \R0_data[11]\, 
        R0_data(10) => \R0_data[10]\, R0_data(9) => \R0_data[9]\, 
        R0_data(8) => \R0_data[8]\, R0_data(7) => \R0_data[7]\, 
        R0_data(6) => \R0_data[6]\, R0_data(5) => \R0_data[5]\, 
        R0_data(4) => \R0_data[4]\, R0_data(3) => \R0_data[3]\, 
        R0_data(2) => \R0_data[2]\, R0_data(1) => \R0_data[1]\, 
        R0_data(0) => \R0_data[0]\, R4_data(31) => \R4_data[31]\, 
        R4_data(30) => \R4_data[30]\, R4_data(29) => 
        \R4_data[29]\, R4_data(28) => \R4_data[28]\, R4_data(27)
         => \R4_data[27]\, R4_data(26) => \R4_data[26]\, 
        R4_data(25) => \R4_data[25]\, R4_data(24) => 
        \R4_data[24]\, R4_data(23) => \R4_data[23]\, R4_data(22)
         => \R4_data[22]\, R4_data(21) => \R4_data[21]\, 
        R4_data(20) => \R4_data[20]\, R4_data(19) => 
        \R4_data[19]\, R4_data(18) => \R4_data[18]\, R4_data(17)
         => \R4_data[17]\, R4_data(16) => \R4_data[16]\, 
        R4_data(15) => \R4_data[15]\, R4_data(14) => 
        \R4_data[14]\, R4_data(13) => \R4_data[13]\, R4_data(12)
         => \R4_data[12]\, R4_data(11) => \R4_data[11]\, 
        R4_data(10) => \R4_data[10]\, R4_data(9) => \R4_data[9]\, 
        R4_data(8) => \R4_data[8]\, R4_data(7) => \R4_data[7]\, 
        R4_data(6) => \R4_data[6]\, R4_data(5) => \R4_data[5]\, 
        R4_data(4) => \R4_data[4]\, R4_data(3) => \R4_data[3]\, 
        R4_data(2) => \R4_data[2]\, R4_data(1) => \R4_data[1]\, 
        R4_data(0) => \R4_data[0]\, N4_data(31) => \N4_data[31]\, 
        N4_data(30) => \N4_data[30]\, N4_data(29) => 
        \N4_data[29]\, N4_data(28) => \N4_data[28]\, N4_data(27)
         => \N4_data[27]\, N4_data(26) => \N4_data[26]\, 
        N4_data(25) => \N4_data[25]\, N4_data(24) => 
        \N4_data[24]\, N4_data(23) => \N4_data[23]\, N4_data(22)
         => \N4_data[22]\, N4_data(21) => \N4_data[21]\, 
        N4_data(20) => \N4_data[20]\, N4_data(19) => 
        \N4_data[19]\, N4_data(18) => \N4_data[18]\, N4_data(17)
         => \N4_data[17]\, N4_data(16) => \N4_data[16]\, 
        N4_data(15) => \N4_data[15]\, N4_data(14) => 
        \N4_data[14]\, N4_data(13) => \N4_data[13]\, N4_data(12)
         => \N4_data[12]\, N4_data(11) => \N4_data[11]\, 
        N4_data(10) => \N4_data[10]\, N4_data(9) => \N4_data[9]\, 
        N4_data(8) => \N4_data[8]\, N4_data(7) => \N4_data[7]\, 
        N4_data(6) => \N4_data[6]\, N4_data(5) => \N4_data[5]\, 
        N4_data(4) => \N4_data[4]\, N4_data(3) => \N4_data[3]\, 
        N4_data(2) => \N4_data[2]\, N4_data(1) => \N4_data[1]\, 
        N0_data(31) => \N0_data[31]\, N0_data(30) => 
        \N0_data[30]\, N0_data(29) => \N0_data[29]\, N0_data(28)
         => \N0_data[28]\, N0_data(27) => \N0_data[27]\, 
        N0_data(26) => \N0_data[26]\, N0_data(25) => 
        \N0_data[25]\, N0_data(24) => \N0_data[24]\, N0_data(23)
         => \N0_data[23]\, N0_data(22) => \N0_data[22]\, 
        N0_data(21) => \N0_data[21]\, N0_data(20) => 
        \N0_data[20]\, N0_data(19) => \N0_data[19]\, N0_data(18)
         => \N0_data[18]\, N0_data(17) => \N0_data[17]\, 
        N0_data(16) => \N0_data[16]\, N0_data(15) => 
        \N0_data[15]\, N0_data(14) => \N0_data[14]\, N0_data(13)
         => \N0_data[13]\, N0_data(12) => \N0_data[12]\, 
        N0_data(11) => \N0_data[11]\, N0_data(10) => 
        \N0_data[10]\, N0_data(9) => \N0_data[9]\, N0_data(8) => 
        \N0_data[8]\, N0_data(7) => \N0_data[7]\, N0_data(6) => 
        \N0_data[6]\, N0_data(5) => \N0_data[5]\, N0_data(4) => 
        \N0_data[4]\, N0_data(3) => \N0_data[3]\, N0_data(2) => 
        \N0_data[2]\, N0_data(1) => \N0_data[1]\, W_out_i_1(0)
         => \W_out_i_1[0]\, Kt_addr(5) => \Kt_addr[5]\, 
        N3_data(31) => \N3_data[31]\, N3_data(30) => 
        \N3_data[30]\, N3_data(29) => \N3_data[29]\, N3_data(28)
         => \N3_data[28]\, N3_data(27) => \N3_data[27]\, 
        N3_data(26) => \N3_data[26]\, N3_data(25) => 
        \N3_data[25]\, N3_data(24) => \N3_data[24]\, N3_data(23)
         => \N3_data[23]\, N3_data(22) => \N3_data[22]\, 
        N3_data(21) => \N3_data[21]\, N3_data(20) => 
        \N3_data[20]\, N3_data(19) => \N3_data[19]\, N3_data(18)
         => \N3_data[18]\, N3_data(17) => \N3_data[17]\, 
        N3_data(16) => \N3_data[16]\, N3_data(15) => 
        \N3_data[15]\, N3_data(14) => \N3_data[14]\, N3_data(13)
         => \N3_data[13]\, N3_data(12) => \N3_data[12]\, 
        N3_data(11) => \N3_data[11]\, N3_data(10) => 
        \N3_data[10]\, N3_data(9) => \N3_data[9]\, N3_data(8) => 
        \N3_data[8]\, N3_data(7) => \N3_data[7]\, N3_data(6) => 
        \N3_data[6]\, N3_data(5) => \N3_data[5]\, N3_data(4) => 
        \N3_data[4]\, N3_data(3) => \N3_data[3]\, N3_data(2) => 
        \N3_data[2]\, N3_data(1) => \N3_data[1]\, N2_data(31) => 
        \N2_data[31]\, N2_data(30) => \N2_data[30]\, N2_data(29)
         => \N2_data[29]\, N2_data(28) => \N2_data[28]\, 
        N2_data(27) => \N2_data[27]\, N2_data(26) => 
        \N2_data[26]\, N2_data(25) => \N2_data[25]\, N2_data(24)
         => \N2_data[24]\, N2_data(23) => \N2_data[23]\, 
        N2_data(22) => \N2_data[22]\, N2_data(21) => 
        \N2_data[21]\, N2_data(20) => \N2_data[20]\, N2_data(19)
         => \N2_data[19]\, N2_data(18) => \N2_data[18]\, 
        N2_data(17) => \N2_data[17]\, N2_data(16) => 
        \N2_data[16]\, N2_data(15) => \N2_data[15]\, N2_data(14)
         => \N2_data[14]\, N2_data(13) => \N2_data[13]\, 
        N2_data(12) => \N2_data[12]\, N2_data(11) => 
        \N2_data[11]\, N2_data(10) => \N2_data[10]\, N2_data(9)
         => \N2_data[9]\, N2_data(8) => \N2_data[8]\, N2_data(7)
         => \N2_data[7]\, N2_data(6) => \N2_data[6]\, N2_data(5)
         => \N2_data[5]\, N2_data(4) => \N2_data[4]\, N2_data(3)
         => \N2_data[3]\, N2_data(2) => \N2_data[2]\, N2_data(1)
         => \N2_data[1]\, N1_data(31) => \N1_data[31]\, 
        N1_data(30) => \N1_data[30]\, N1_data(29) => 
        \N1_data[29]\, N1_data(28) => \N1_data[28]\, N1_data(27)
         => \N1_data[27]\, N1_data(26) => \N1_data[26]\, 
        N1_data(25) => \N1_data[25]\, N1_data(24) => 
        \N1_data[24]\, N1_data(23) => \N1_data[23]\, N1_data(22)
         => \N1_data[22]\, N1_data(21) => \N1_data[21]\, 
        N1_data(20) => \N1_data[20]\, N1_data(19) => 
        \N1_data[19]\, N1_data(18) => \N1_data[18]\, N1_data(17)
         => \N1_data[17]\, N1_data(16) => \N1_data[16]\, 
        N1_data(15) => \N1_data[15]\, N1_data(14) => 
        \N1_data[14]\, N1_data(13) => \N1_data[13]\, N1_data(12)
         => \N1_data[12]\, N1_data(11) => \N1_data[11]\, 
        N1_data(10) => \N1_data[10]\, N1_data(9) => \N1_data[9]\, 
        N1_data(8) => \N1_data[8]\, N1_data(7) => \N1_data[7]\, 
        N1_data(6) => \N1_data[6]\, N1_data(5) => \N1_data[5]\, 
        N1_data(4) => \N1_data[4]\, N1_data(3) => \N1_data[3]\, 
        N1_data(2) => \N1_data[2]\, N1_data(1) => \N1_data[1]\, 
        N7_data(31) => \N7_data[31]\, N7_data(30) => 
        \N7_data[30]\, N7_data(29) => \N7_data[29]\, N7_data(28)
         => \N7_data[28]\, N7_data(27) => \N7_data[27]\, 
        N7_data(26) => \N7_data[26]\, N7_data(25) => 
        \N7_data[25]\, N7_data(24) => \N7_data[24]\, N7_data(23)
         => \N7_data[23]\, N7_data(22) => \N7_data[22]\, 
        N7_data(21) => \N7_data[21]\, N7_data(20) => 
        \N7_data[20]\, N7_data(19) => \N7_data[19]\, N7_data(18)
         => \N7_data[18]\, N7_data(17) => \N7_data[17]\, 
        N7_data(16) => \N7_data[16]\, N7_data(15) => 
        \N7_data[15]\, N7_data(14) => \N7_data[14]\, N7_data(13)
         => \N7_data[13]\, N7_data(12) => \N7_data[12]\, 
        N7_data(11) => \N7_data[11]\, N7_data(10) => 
        \N7_data[10]\, N7_data(9) => \N7_data[9]\, N7_data(8) => 
        \N7_data[8]\, N7_data(7) => \N7_data[7]\, N7_data(6) => 
        \N7_data[6]\, N7_data(5) => \N7_data[5]\, N7_data(4) => 
        \N7_data[4]\, N7_data(3) => \N7_data[3]\, N7_data(2) => 
        \N7_data[2]\, N7_data(1) => \N7_data[1]\, N6_data(31) => 
        \N6_data[31]\, N6_data(30) => \N6_data[30]\, N6_data(29)
         => \N6_data[29]\, N6_data(28) => \N6_data[28]\, 
        N6_data(27) => \N6_data[27]\, N6_data(26) => 
        \N6_data[26]\, N6_data(25) => \N6_data[25]\, N6_data(24)
         => \N6_data[24]\, N6_data(23) => \N6_data[23]\, 
        N6_data(22) => \N6_data[22]\, N6_data(21) => 
        \N6_data[21]\, N6_data(20) => \N6_data[20]\, N6_data(19)
         => \N6_data[19]\, N6_data(18) => \N6_data[18]\, 
        N6_data(17) => \N6_data[17]\, N6_data(16) => 
        \N6_data[16]\, N6_data(15) => \N6_data[15]\, N6_data(14)
         => \N6_data[14]\, N6_data(13) => \N6_data[13]\, 
        N6_data(12) => \N6_data[12]\, N6_data(11) => 
        \N6_data[11]\, N6_data(10) => \N6_data[10]\, N6_data(9)
         => \N6_data[9]\, N6_data(8) => \N6_data[8]\, N6_data(7)
         => \N6_data[7]\, N6_data(6) => \N6_data[6]\, N6_data(5)
         => \N6_data[5]\, N6_data(4) => \N6_data[4]\, N6_data(3)
         => \N6_data[3]\, N6_data(2) => \N6_data[2]\, N6_data(1)
         => \N6_data[1]\, N5_data(31) => \N5_data[31]\, 
        N5_data(30) => \N5_data[30]\, N5_data(29) => 
        \N5_data[29]\, N5_data(28) => \N5_data[28]\, N5_data(27)
         => \N5_data[27]\, N5_data(26) => \N5_data[26]\, 
        N5_data(25) => \N5_data[25]\, N5_data(24) => 
        \N5_data[24]\, N5_data(23) => \N5_data[23]\, N5_data(22)
         => \N5_data[22]\, N5_data(21) => \N5_data[21]\, 
        N5_data(20) => \N5_data[20]\, N5_data(19) => 
        \N5_data[19]\, N5_data(18) => \N5_data[18]\, N5_data(17)
         => \N5_data[17]\, N5_data(16) => \N5_data[16]\, 
        N5_data(15) => \N5_data[15]\, N5_data(14) => 
        \N5_data[14]\, N5_data(13) => \N5_data[13]\, N5_data(12)
         => \N5_data[12]\, N5_data(11) => \N5_data[11]\, 
        N5_data(10) => \N5_data[10]\, N5_data(9) => \N5_data[9]\, 
        N5_data(8) => \N5_data[8]\, N5_data(7) => \N5_data[7]\, 
        N5_data(6) => \N5_data[6]\, N5_data(5) => \N5_data[5]\, 
        N5_data(4) => \N5_data[4]\, N5_data(3) => \N5_data[3]\, 
        N5_data(2) => \N5_data[2]\, N5_data(1) => \N5_data[1]\, 
        Wt_data(31) => \Wt_data[31]\, Wt_data(30) => 
        \Wt_data[30]\, Wt_data(29) => \Wt_data[29]\, Wt_data(28)
         => \Wt_data[28]\, Wt_data(27) => \Wt_data[27]\, 
        Wt_data(26) => \Wt_data[26]\, Wt_data(25) => 
        \Wt_data[25]\, Wt_data(24) => \Wt_data[24]\, Wt_data(23)
         => \Wt_data[23]\, Wt_data(22) => \Wt_data[22]\, 
        Wt_data(21) => \Wt_data[21]\, Wt_data(20) => 
        \Wt_data[20]\, Wt_data(19) => \Wt_data[19]\, Wt_data(18)
         => \Wt_data[18]\, Wt_data(17) => \Wt_data[17]\, 
        Wt_data(16) => \Wt_data[16]\, Wt_data(15) => 
        \Wt_data[15]\, Wt_data(14) => \Wt_data[14]\, Wt_data(13)
         => \Wt_data[13]\, Wt_data(12) => \Wt_data[12]\, 
        Wt_data(11) => \Wt_data[11]\, Wt_data(10) => 
        \Wt_data[10]\, Wt_data(9) => \Wt_data[9]\, Wt_data(8) => 
        \Wt_data[8]\, Wt_data(7) => \Wt_data[7]\, Wt_data(6) => 
        \Wt_data[6]\, Wt_data(5) => \Wt_data[5]\, Wt_data(4) => 
        \Wt_data[4]\, Wt_data(3) => \Wt_data[3]\, Wt_data(2) => 
        \Wt_data[2]\, Wt_data(1) => \Wt_data[1]\, Wt_data(0) => 
        \Wt_data[0]\, Kt_data_0 => \Kt_data[15]\, Kt_data_9 => 
        \Kt_data[24]\, CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, core_ce_o_iv_i_0
         => core_ce_o_iv_i_0, oregs_ce_i_a2_0_a2 => 
        oregs_ce_i_a2_0_a2, next_reg_H4_cry_0_0_Y => 
        next_reg_H4_cry_0_0_Y, next_reg_H0_cry_0_0_Y => 
        next_reg_H0_cry_0_0_Y, next_r0_0_cry_0_Y => 
        next_r0_0_cry_0_Y, ld_i_i_3 => ld_i_i_3, N_98 => N_98, 
        m34 => m34, m49_am => m49_am, m49_bm => m49_bm, m62_am
         => m62_am, m62_bm => m62_bm, m67_ns => m67_ns, m73 => 
        m73, m78 => m78, m83_ns => m83_ns, m95_1_0 => m95_1_0, 
        m95_1_1 => m95_1_1, m104_am => m104_am, m104_bm => 
        m104_bm, m110_ns => m110_ns, m114 => m114, m119_ns => 
        m119_ns, m124 => m124, m137_am => m137_am, m137_bm => 
        m137_bm, m141 => m141, m144_ns => m144_ns, m157 => m157, 
        m168_1_0 => m168_1_0, m168_1_1 => m168_1_1, m172_ns => 
        m172_ns, m177 => m177, m197_1_0 => m197_1_0, m197_1_1 => 
        m197_1_1, m207_1_0 => m207_1_0, m207_1_1 => m207_1_1, 
        m215_am => m215_am, m215_bm => m215_bm, m219 => m219, 
        m222_ns => m222_ns, m226_ns => m226_ns, m230 => m230, 
        m235_ns => m235_ns, m239 => m239, m250_am => m250_am, 
        m250_bm => m250_bm, m254 => m254, m258_ns => m258_ns, 
        m273 => m273, m276_ns => m276_ns, m281_ns => m281_ns, 
        m285 => m285, m289 => m289, m292_ns => m292_ns, m296 => 
        m296, m300_ns => m300_ns, m304 => m304, i3_mux_1 => 
        i3_mux_1, m325 => m325, m316 => m316, 
        next_reg_H3_cry_0_0_Y => next_reg_H3_cry_0_0_Y, 
        next_reg_H2_cry_0_0_Y => next_reg_H2_cry_0_0_Y, 
        next_reg_H1_cry_0_0_Y => next_reg_H1_cry_0_0_Y, 
        next_reg_H7_cry_0_0_Y => next_reg_H7_cry_0_0_Y, 
        next_reg_H6_cry_0_0_Y => next_reg_H6_cry_0_0_Y, 
        next_reg_H5_cry_0_0_Y => next_reg_H5_cry_0_0_Y, m10_ns
         => m10_ns, m19 => m19);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    Inst_sha256_regs : sha256_regs
      port map(SHA256_BLOCK_0_H0_o(31) => SHA256_BLOCK_0_H0_o(31), 
        SHA256_BLOCK_0_H0_o(30) => SHA256_BLOCK_0_H0_o(30), 
        SHA256_BLOCK_0_H0_o(29) => SHA256_BLOCK_0_H0_o(29), 
        SHA256_BLOCK_0_H0_o(28) => SHA256_BLOCK_0_H0_o(28), 
        SHA256_BLOCK_0_H0_o(27) => SHA256_BLOCK_0_H0_o(27), 
        SHA256_BLOCK_0_H0_o(26) => SHA256_BLOCK_0_H0_o(26), 
        SHA256_BLOCK_0_H0_o(25) => SHA256_BLOCK_0_H0_o(25), 
        SHA256_BLOCK_0_H0_o(24) => SHA256_BLOCK_0_H0_o(24), 
        SHA256_BLOCK_0_H0_o(23) => SHA256_BLOCK_0_H0_o(23), 
        SHA256_BLOCK_0_H0_o(22) => SHA256_BLOCK_0_H0_o(22), 
        SHA256_BLOCK_0_H0_o(21) => SHA256_BLOCK_0_H0_o(21), 
        SHA256_BLOCK_0_H0_o(20) => SHA256_BLOCK_0_H0_o(20), 
        SHA256_BLOCK_0_H0_o(19) => SHA256_BLOCK_0_H0_o(19), 
        SHA256_BLOCK_0_H0_o(18) => SHA256_BLOCK_0_H0_o(18), 
        SHA256_BLOCK_0_H0_o(17) => SHA256_BLOCK_0_H0_o(17), 
        SHA256_BLOCK_0_H0_o(16) => SHA256_BLOCK_0_H0_o(16), 
        SHA256_BLOCK_0_H0_o(15) => SHA256_BLOCK_0_H0_o(15), 
        SHA256_BLOCK_0_H0_o(14) => SHA256_BLOCK_0_H0_o(14), 
        SHA256_BLOCK_0_H0_o(13) => SHA256_BLOCK_0_H0_o(13), 
        SHA256_BLOCK_0_H0_o(12) => SHA256_BLOCK_0_H0_o(12), 
        SHA256_BLOCK_0_H0_o(11) => SHA256_BLOCK_0_H0_o(11), 
        SHA256_BLOCK_0_H0_o(10) => SHA256_BLOCK_0_H0_o(10), 
        SHA256_BLOCK_0_H0_o(9) => SHA256_BLOCK_0_H0_o(9), 
        SHA256_BLOCK_0_H0_o(8) => SHA256_BLOCK_0_H0_o(8), 
        SHA256_BLOCK_0_H0_o(7) => SHA256_BLOCK_0_H0_o(7), 
        SHA256_BLOCK_0_H0_o(6) => SHA256_BLOCK_0_H0_o(6), 
        SHA256_BLOCK_0_H0_o(5) => SHA256_BLOCK_0_H0_o(5), 
        SHA256_BLOCK_0_H0_o(4) => SHA256_BLOCK_0_H0_o(4), 
        SHA256_BLOCK_0_H0_o(3) => SHA256_BLOCK_0_H0_o(3), 
        SHA256_BLOCK_0_H0_o(2) => SHA256_BLOCK_0_H0_o(2), 
        SHA256_BLOCK_0_H0_o(1) => SHA256_BLOCK_0_H0_o(1), 
        SHA256_BLOCK_0_H0_o(0) => SHA256_BLOCK_0_H0_o(0), 
        N0_data(31) => \N0_data[31]\, N0_data(30) => 
        \N0_data[30]\, N0_data(29) => \N0_data[29]\, N0_data(28)
         => \N0_data[28]\, N0_data(27) => \N0_data[27]\, 
        N0_data(26) => \N0_data[26]\, N0_data(25) => 
        \N0_data[25]\, N0_data(24) => \N0_data[24]\, N0_data(23)
         => \N0_data[23]\, N0_data(22) => \N0_data[22]\, 
        N0_data(21) => \N0_data[21]\, N0_data(20) => 
        \N0_data[20]\, N0_data(19) => \N0_data[19]\, N0_data(18)
         => \N0_data[18]\, N0_data(17) => \N0_data[17]\, 
        N0_data(16) => \N0_data[16]\, N0_data(15) => 
        \N0_data[15]\, N0_data(14) => \N0_data[14]\, N0_data(13)
         => \N0_data[13]\, N0_data(12) => \N0_data[12]\, 
        N0_data(11) => \N0_data[11]\, N0_data(10) => 
        \N0_data[10]\, N0_data(9) => \N0_data[9]\, N0_data(8) => 
        \N0_data[8]\, N0_data(7) => \N0_data[7]\, N0_data(6) => 
        \N0_data[6]\, N0_data(5) => \N0_data[5]\, N0_data(4) => 
        \N0_data[4]\, N0_data(3) => \N0_data[3]\, N0_data(2) => 
        \N0_data[2]\, N0_data(1) => \N0_data[1]\, 
        SHA256_BLOCK_0_H1_o(31) => SHA256_BLOCK_0_H1_o(31), 
        SHA256_BLOCK_0_H1_o(30) => SHA256_BLOCK_0_H1_o(30), 
        SHA256_BLOCK_0_H1_o(29) => SHA256_BLOCK_0_H1_o(29), 
        SHA256_BLOCK_0_H1_o(28) => SHA256_BLOCK_0_H1_o(28), 
        SHA256_BLOCK_0_H1_o(27) => SHA256_BLOCK_0_H1_o(27), 
        SHA256_BLOCK_0_H1_o(26) => SHA256_BLOCK_0_H1_o(26), 
        SHA256_BLOCK_0_H1_o(25) => SHA256_BLOCK_0_H1_o(25), 
        SHA256_BLOCK_0_H1_o(24) => SHA256_BLOCK_0_H1_o(24), 
        SHA256_BLOCK_0_H1_o(23) => SHA256_BLOCK_0_H1_o(23), 
        SHA256_BLOCK_0_H1_o(22) => SHA256_BLOCK_0_H1_o(22), 
        SHA256_BLOCK_0_H1_o(21) => SHA256_BLOCK_0_H1_o(21), 
        SHA256_BLOCK_0_H1_o(20) => SHA256_BLOCK_0_H1_o(20), 
        SHA256_BLOCK_0_H1_o(19) => SHA256_BLOCK_0_H1_o(19), 
        SHA256_BLOCK_0_H1_o(18) => SHA256_BLOCK_0_H1_o(18), 
        SHA256_BLOCK_0_H1_o(17) => SHA256_BLOCK_0_H1_o(17), 
        SHA256_BLOCK_0_H1_o(16) => SHA256_BLOCK_0_H1_o(16), 
        SHA256_BLOCK_0_H1_o(15) => SHA256_BLOCK_0_H1_o(15), 
        SHA256_BLOCK_0_H1_o(14) => SHA256_BLOCK_0_H1_o(14), 
        SHA256_BLOCK_0_H1_o(13) => SHA256_BLOCK_0_H1_o(13), 
        SHA256_BLOCK_0_H1_o(12) => SHA256_BLOCK_0_H1_o(12), 
        SHA256_BLOCK_0_H1_o(11) => SHA256_BLOCK_0_H1_o(11), 
        SHA256_BLOCK_0_H1_o(10) => SHA256_BLOCK_0_H1_o(10), 
        SHA256_BLOCK_0_H1_o(9) => SHA256_BLOCK_0_H1_o(9), 
        SHA256_BLOCK_0_H1_o(8) => SHA256_BLOCK_0_H1_o(8), 
        SHA256_BLOCK_0_H1_o(7) => SHA256_BLOCK_0_H1_o(7), 
        SHA256_BLOCK_0_H1_o(6) => SHA256_BLOCK_0_H1_o(6), 
        SHA256_BLOCK_0_H1_o(5) => SHA256_BLOCK_0_H1_o(5), 
        SHA256_BLOCK_0_H1_o(4) => SHA256_BLOCK_0_H1_o(4), 
        SHA256_BLOCK_0_H1_o(3) => SHA256_BLOCK_0_H1_o(3), 
        SHA256_BLOCK_0_H1_o(2) => SHA256_BLOCK_0_H1_o(2), 
        SHA256_BLOCK_0_H1_o(1) => SHA256_BLOCK_0_H1_o(1), 
        SHA256_BLOCK_0_H1_o(0) => SHA256_BLOCK_0_H1_o(0), 
        N1_data(31) => \N1_data[31]\, N1_data(30) => 
        \N1_data[30]\, N1_data(29) => \N1_data[29]\, N1_data(28)
         => \N1_data[28]\, N1_data(27) => \N1_data[27]\, 
        N1_data(26) => \N1_data[26]\, N1_data(25) => 
        \N1_data[25]\, N1_data(24) => \N1_data[24]\, N1_data(23)
         => \N1_data[23]\, N1_data(22) => \N1_data[22]\, 
        N1_data(21) => \N1_data[21]\, N1_data(20) => 
        \N1_data[20]\, N1_data(19) => \N1_data[19]\, N1_data(18)
         => \N1_data[18]\, N1_data(17) => \N1_data[17]\, 
        N1_data(16) => \N1_data[16]\, N1_data(15) => 
        \N1_data[15]\, N1_data(14) => \N1_data[14]\, N1_data(13)
         => \N1_data[13]\, N1_data(12) => \N1_data[12]\, 
        N1_data(11) => \N1_data[11]\, N1_data(10) => 
        \N1_data[10]\, N1_data(9) => \N1_data[9]\, N1_data(8) => 
        \N1_data[8]\, N1_data(7) => \N1_data[7]\, N1_data(6) => 
        \N1_data[6]\, N1_data(5) => \N1_data[5]\, N1_data(4) => 
        \N1_data[4]\, N1_data(3) => \N1_data[3]\, N1_data(2) => 
        \N1_data[2]\, N1_data(1) => \N1_data[1]\, 
        SHA256_BLOCK_0_H2_o(31) => SHA256_BLOCK_0_H2_o(31), 
        SHA256_BLOCK_0_H2_o(30) => SHA256_BLOCK_0_H2_o(30), 
        SHA256_BLOCK_0_H2_o(29) => SHA256_BLOCK_0_H2_o(29), 
        SHA256_BLOCK_0_H2_o(28) => SHA256_BLOCK_0_H2_o(28), 
        SHA256_BLOCK_0_H2_o(27) => SHA256_BLOCK_0_H2_o(27), 
        SHA256_BLOCK_0_H2_o(26) => SHA256_BLOCK_0_H2_o(26), 
        SHA256_BLOCK_0_H2_o(25) => SHA256_BLOCK_0_H2_o(25), 
        SHA256_BLOCK_0_H2_o(24) => SHA256_BLOCK_0_H2_o(24), 
        SHA256_BLOCK_0_H2_o(23) => SHA256_BLOCK_0_H2_o(23), 
        SHA256_BLOCK_0_H2_o(22) => SHA256_BLOCK_0_H2_o(22), 
        SHA256_BLOCK_0_H2_o(21) => SHA256_BLOCK_0_H2_o(21), 
        SHA256_BLOCK_0_H2_o(20) => SHA256_BLOCK_0_H2_o(20), 
        SHA256_BLOCK_0_H2_o(19) => SHA256_BLOCK_0_H2_o(19), 
        SHA256_BLOCK_0_H2_o(18) => SHA256_BLOCK_0_H2_o(18), 
        SHA256_BLOCK_0_H2_o(17) => SHA256_BLOCK_0_H2_o(17), 
        SHA256_BLOCK_0_H2_o(16) => SHA256_BLOCK_0_H2_o(16), 
        SHA256_BLOCK_0_H2_o(15) => SHA256_BLOCK_0_H2_o(15), 
        SHA256_BLOCK_0_H2_o(14) => SHA256_BLOCK_0_H2_o(14), 
        SHA256_BLOCK_0_H2_o(13) => SHA256_BLOCK_0_H2_o(13), 
        SHA256_BLOCK_0_H2_o(12) => SHA256_BLOCK_0_H2_o(12), 
        SHA256_BLOCK_0_H2_o(11) => SHA256_BLOCK_0_H2_o(11), 
        SHA256_BLOCK_0_H2_o(10) => SHA256_BLOCK_0_H2_o(10), 
        SHA256_BLOCK_0_H2_o(9) => SHA256_BLOCK_0_H2_o(9), 
        SHA256_BLOCK_0_H2_o(8) => SHA256_BLOCK_0_H2_o(8), 
        SHA256_BLOCK_0_H2_o(7) => SHA256_BLOCK_0_H2_o(7), 
        SHA256_BLOCK_0_H2_o(6) => SHA256_BLOCK_0_H2_o(6), 
        SHA256_BLOCK_0_H2_o(5) => SHA256_BLOCK_0_H2_o(5), 
        SHA256_BLOCK_0_H2_o(4) => SHA256_BLOCK_0_H2_o(4), 
        SHA256_BLOCK_0_H2_o(3) => SHA256_BLOCK_0_H2_o(3), 
        SHA256_BLOCK_0_H2_o(2) => SHA256_BLOCK_0_H2_o(2), 
        SHA256_BLOCK_0_H2_o(1) => SHA256_BLOCK_0_H2_o(1), 
        SHA256_BLOCK_0_H2_o(0) => SHA256_BLOCK_0_H2_o(0), 
        N2_data(31) => \N2_data[31]\, N2_data(30) => 
        \N2_data[30]\, N2_data(29) => \N2_data[29]\, N2_data(28)
         => \N2_data[28]\, N2_data(27) => \N2_data[27]\, 
        N2_data(26) => \N2_data[26]\, N2_data(25) => 
        \N2_data[25]\, N2_data(24) => \N2_data[24]\, N2_data(23)
         => \N2_data[23]\, N2_data(22) => \N2_data[22]\, 
        N2_data(21) => \N2_data[21]\, N2_data(20) => 
        \N2_data[20]\, N2_data(19) => \N2_data[19]\, N2_data(18)
         => \N2_data[18]\, N2_data(17) => \N2_data[17]\, 
        N2_data(16) => \N2_data[16]\, N2_data(15) => 
        \N2_data[15]\, N2_data(14) => \N2_data[14]\, N2_data(13)
         => \N2_data[13]\, N2_data(12) => \N2_data[12]\, 
        N2_data(11) => \N2_data[11]\, N2_data(10) => 
        \N2_data[10]\, N2_data(9) => \N2_data[9]\, N2_data(8) => 
        \N2_data[8]\, N2_data(7) => \N2_data[7]\, N2_data(6) => 
        \N2_data[6]\, N2_data(5) => \N2_data[5]\, N2_data(4) => 
        \N2_data[4]\, N2_data(3) => \N2_data[3]\, N2_data(2) => 
        \N2_data[2]\, N2_data(1) => \N2_data[1]\, 
        SHA256_BLOCK_0_H3_o(31) => SHA256_BLOCK_0_H3_o(31), 
        SHA256_BLOCK_0_H3_o(30) => SHA256_BLOCK_0_H3_o(30), 
        SHA256_BLOCK_0_H3_o(29) => SHA256_BLOCK_0_H3_o(29), 
        SHA256_BLOCK_0_H3_o(28) => SHA256_BLOCK_0_H3_o(28), 
        SHA256_BLOCK_0_H3_o(27) => SHA256_BLOCK_0_H3_o(27), 
        SHA256_BLOCK_0_H3_o(26) => SHA256_BLOCK_0_H3_o(26), 
        SHA256_BLOCK_0_H3_o(25) => SHA256_BLOCK_0_H3_o(25), 
        SHA256_BLOCK_0_H3_o(24) => SHA256_BLOCK_0_H3_o(24), 
        SHA256_BLOCK_0_H3_o(23) => SHA256_BLOCK_0_H3_o(23), 
        SHA256_BLOCK_0_H3_o(22) => SHA256_BLOCK_0_H3_o(22), 
        SHA256_BLOCK_0_H3_o(21) => SHA256_BLOCK_0_H3_o(21), 
        SHA256_BLOCK_0_H3_o(20) => SHA256_BLOCK_0_H3_o(20), 
        SHA256_BLOCK_0_H3_o(19) => SHA256_BLOCK_0_H3_o(19), 
        SHA256_BLOCK_0_H3_o(18) => SHA256_BLOCK_0_H3_o(18), 
        SHA256_BLOCK_0_H3_o(17) => SHA256_BLOCK_0_H3_o(17), 
        SHA256_BLOCK_0_H3_o(16) => SHA256_BLOCK_0_H3_o(16), 
        SHA256_BLOCK_0_H3_o(15) => SHA256_BLOCK_0_H3_o(15), 
        SHA256_BLOCK_0_H3_o(14) => SHA256_BLOCK_0_H3_o(14), 
        SHA256_BLOCK_0_H3_o(13) => SHA256_BLOCK_0_H3_o(13), 
        SHA256_BLOCK_0_H3_o(12) => SHA256_BLOCK_0_H3_o(12), 
        SHA256_BLOCK_0_H3_o(11) => SHA256_BLOCK_0_H3_o(11), 
        SHA256_BLOCK_0_H3_o(10) => SHA256_BLOCK_0_H3_o(10), 
        SHA256_BLOCK_0_H3_o(9) => SHA256_BLOCK_0_H3_o(9), 
        SHA256_BLOCK_0_H3_o(8) => SHA256_BLOCK_0_H3_o(8), 
        SHA256_BLOCK_0_H3_o(7) => SHA256_BLOCK_0_H3_o(7), 
        SHA256_BLOCK_0_H3_o(6) => SHA256_BLOCK_0_H3_o(6), 
        SHA256_BLOCK_0_H3_o(5) => SHA256_BLOCK_0_H3_o(5), 
        SHA256_BLOCK_0_H3_o(4) => SHA256_BLOCK_0_H3_o(4), 
        SHA256_BLOCK_0_H3_o(3) => SHA256_BLOCK_0_H3_o(3), 
        SHA256_BLOCK_0_H3_o(2) => SHA256_BLOCK_0_H3_o(2), 
        SHA256_BLOCK_0_H3_o(1) => SHA256_BLOCK_0_H3_o(1), 
        SHA256_BLOCK_0_H3_o(0) => SHA256_BLOCK_0_H3_o(0), 
        N3_data(31) => \N3_data[31]\, N3_data(30) => 
        \N3_data[30]\, N3_data(29) => \N3_data[29]\, N3_data(28)
         => \N3_data[28]\, N3_data(27) => \N3_data[27]\, 
        N3_data(26) => \N3_data[26]\, N3_data(25) => 
        \N3_data[25]\, N3_data(24) => \N3_data[24]\, N3_data(23)
         => \N3_data[23]\, N3_data(22) => \N3_data[22]\, 
        N3_data(21) => \N3_data[21]\, N3_data(20) => 
        \N3_data[20]\, N3_data(19) => \N3_data[19]\, N3_data(18)
         => \N3_data[18]\, N3_data(17) => \N3_data[17]\, 
        N3_data(16) => \N3_data[16]\, N3_data(15) => 
        \N3_data[15]\, N3_data(14) => \N3_data[14]\, N3_data(13)
         => \N3_data[13]\, N3_data(12) => \N3_data[12]\, 
        N3_data(11) => \N3_data[11]\, N3_data(10) => 
        \N3_data[10]\, N3_data(9) => \N3_data[9]\, N3_data(8) => 
        \N3_data[8]\, N3_data(7) => \N3_data[7]\, N3_data(6) => 
        \N3_data[6]\, N3_data(5) => \N3_data[5]\, N3_data(4) => 
        \N3_data[4]\, N3_data(3) => \N3_data[3]\, N3_data(2) => 
        \N3_data[2]\, N3_data(1) => \N3_data[1]\, 
        SHA256_BLOCK_0_H4_o(31) => SHA256_BLOCK_0_H4_o(31), 
        SHA256_BLOCK_0_H4_o(30) => SHA256_BLOCK_0_H4_o(30), 
        SHA256_BLOCK_0_H4_o(29) => SHA256_BLOCK_0_H4_o(29), 
        SHA256_BLOCK_0_H4_o(28) => SHA256_BLOCK_0_H4_o(28), 
        SHA256_BLOCK_0_H4_o(27) => SHA256_BLOCK_0_H4_o(27), 
        SHA256_BLOCK_0_H4_o(26) => SHA256_BLOCK_0_H4_o(26), 
        SHA256_BLOCK_0_H4_o(25) => SHA256_BLOCK_0_H4_o(25), 
        SHA256_BLOCK_0_H4_o(24) => SHA256_BLOCK_0_H4_o(24), 
        SHA256_BLOCK_0_H4_o(23) => SHA256_BLOCK_0_H4_o(23), 
        SHA256_BLOCK_0_H4_o(22) => SHA256_BLOCK_0_H4_o(22), 
        SHA256_BLOCK_0_H4_o(21) => SHA256_BLOCK_0_H4_o(21), 
        SHA256_BLOCK_0_H4_o(20) => SHA256_BLOCK_0_H4_o(20), 
        SHA256_BLOCK_0_H4_o(19) => SHA256_BLOCK_0_H4_o(19), 
        SHA256_BLOCK_0_H4_o(18) => SHA256_BLOCK_0_H4_o(18), 
        SHA256_BLOCK_0_H4_o(17) => SHA256_BLOCK_0_H4_o(17), 
        SHA256_BLOCK_0_H4_o(16) => SHA256_BLOCK_0_H4_o(16), 
        SHA256_BLOCK_0_H4_o(15) => SHA256_BLOCK_0_H4_o(15), 
        SHA256_BLOCK_0_H4_o(14) => SHA256_BLOCK_0_H4_o(14), 
        SHA256_BLOCK_0_H4_o(13) => SHA256_BLOCK_0_H4_o(13), 
        SHA256_BLOCK_0_H4_o(12) => SHA256_BLOCK_0_H4_o(12), 
        SHA256_BLOCK_0_H4_o(11) => SHA256_BLOCK_0_H4_o(11), 
        SHA256_BLOCK_0_H4_o(10) => SHA256_BLOCK_0_H4_o(10), 
        SHA256_BLOCK_0_H4_o(9) => SHA256_BLOCK_0_H4_o(9), 
        SHA256_BLOCK_0_H4_o(8) => SHA256_BLOCK_0_H4_o(8), 
        SHA256_BLOCK_0_H4_o(7) => SHA256_BLOCK_0_H4_o(7), 
        SHA256_BLOCK_0_H4_o(6) => SHA256_BLOCK_0_H4_o(6), 
        SHA256_BLOCK_0_H4_o(5) => SHA256_BLOCK_0_H4_o(5), 
        SHA256_BLOCK_0_H4_o(4) => SHA256_BLOCK_0_H4_o(4), 
        SHA256_BLOCK_0_H4_o(3) => SHA256_BLOCK_0_H4_o(3), 
        SHA256_BLOCK_0_H4_o(2) => SHA256_BLOCK_0_H4_o(2), 
        SHA256_BLOCK_0_H4_o(1) => SHA256_BLOCK_0_H4_o(1), 
        SHA256_BLOCK_0_H4_o(0) => SHA256_BLOCK_0_H4_o(0), 
        N4_data(31) => \N4_data[31]\, N4_data(30) => 
        \N4_data[30]\, N4_data(29) => \N4_data[29]\, N4_data(28)
         => \N4_data[28]\, N4_data(27) => \N4_data[27]\, 
        N4_data(26) => \N4_data[26]\, N4_data(25) => 
        \N4_data[25]\, N4_data(24) => \N4_data[24]\, N4_data(23)
         => \N4_data[23]\, N4_data(22) => \N4_data[22]\, 
        N4_data(21) => \N4_data[21]\, N4_data(20) => 
        \N4_data[20]\, N4_data(19) => \N4_data[19]\, N4_data(18)
         => \N4_data[18]\, N4_data(17) => \N4_data[17]\, 
        N4_data(16) => \N4_data[16]\, N4_data(15) => 
        \N4_data[15]\, N4_data(14) => \N4_data[14]\, N4_data(13)
         => \N4_data[13]\, N4_data(12) => \N4_data[12]\, 
        N4_data(11) => \N4_data[11]\, N4_data(10) => 
        \N4_data[10]\, N4_data(9) => \N4_data[9]\, N4_data(8) => 
        \N4_data[8]\, N4_data(7) => \N4_data[7]\, N4_data(6) => 
        \N4_data[6]\, N4_data(5) => \N4_data[5]\, N4_data(4) => 
        \N4_data[4]\, N4_data(3) => \N4_data[3]\, N4_data(2) => 
        \N4_data[2]\, N4_data(1) => \N4_data[1]\, N5_data(31) => 
        \N5_data[31]\, N5_data(30) => \N5_data[30]\, N5_data(29)
         => \N5_data[29]\, N5_data(28) => \N5_data[28]\, 
        N5_data(27) => \N5_data[27]\, N5_data(26) => 
        \N5_data[26]\, N5_data(25) => \N5_data[25]\, N5_data(24)
         => \N5_data[24]\, N5_data(23) => \N5_data[23]\, 
        N5_data(22) => \N5_data[22]\, N5_data(21) => 
        \N5_data[21]\, N5_data(20) => \N5_data[20]\, N5_data(19)
         => \N5_data[19]\, N5_data(18) => \N5_data[18]\, 
        N5_data(17) => \N5_data[17]\, N5_data(16) => 
        \N5_data[16]\, N5_data(15) => \N5_data[15]\, N5_data(14)
         => \N5_data[14]\, N5_data(13) => \N5_data[13]\, 
        N5_data(12) => \N5_data[12]\, N5_data(11) => 
        \N5_data[11]\, N5_data(10) => \N5_data[10]\, N5_data(9)
         => \N5_data[9]\, N5_data(8) => \N5_data[8]\, N5_data(7)
         => \N5_data[7]\, N5_data(6) => \N5_data[6]\, N5_data(5)
         => \N5_data[5]\, N5_data(4) => \N5_data[4]\, N5_data(3)
         => \N5_data[3]\, N5_data(2) => \N5_data[2]\, N5_data(1)
         => \N5_data[1]\, SHA256_BLOCK_0_H5_o(31) => 
        SHA256_BLOCK_0_H5_o(31), SHA256_BLOCK_0_H5_o(30) => 
        SHA256_BLOCK_0_H5_o(30), SHA256_BLOCK_0_H5_o(29) => 
        SHA256_BLOCK_0_H5_o(29), SHA256_BLOCK_0_H5_o(28) => 
        SHA256_BLOCK_0_H5_o(28), SHA256_BLOCK_0_H5_o(27) => 
        SHA256_BLOCK_0_H5_o(27), SHA256_BLOCK_0_H5_o(26) => 
        SHA256_BLOCK_0_H5_o(26), SHA256_BLOCK_0_H5_o(25) => 
        SHA256_BLOCK_0_H5_o(25), SHA256_BLOCK_0_H5_o(24) => 
        SHA256_BLOCK_0_H5_o(24), SHA256_BLOCK_0_H5_o(23) => 
        SHA256_BLOCK_0_H5_o(23), SHA256_BLOCK_0_H5_o(22) => 
        SHA256_BLOCK_0_H5_o(22), SHA256_BLOCK_0_H5_o(21) => 
        SHA256_BLOCK_0_H5_o(21), SHA256_BLOCK_0_H5_o(20) => 
        SHA256_BLOCK_0_H5_o(20), SHA256_BLOCK_0_H5_o(19) => 
        SHA256_BLOCK_0_H5_o(19), SHA256_BLOCK_0_H5_o(18) => 
        SHA256_BLOCK_0_H5_o(18), SHA256_BLOCK_0_H5_o(17) => 
        SHA256_BLOCK_0_H5_o(17), SHA256_BLOCK_0_H5_o(16) => 
        SHA256_BLOCK_0_H5_o(16), SHA256_BLOCK_0_H5_o(15) => 
        SHA256_BLOCK_0_H5_o(15), SHA256_BLOCK_0_H5_o(14) => 
        SHA256_BLOCK_0_H5_o(14), SHA256_BLOCK_0_H5_o(13) => 
        SHA256_BLOCK_0_H5_o(13), SHA256_BLOCK_0_H5_o(12) => 
        SHA256_BLOCK_0_H5_o(12), SHA256_BLOCK_0_H5_o(11) => 
        SHA256_BLOCK_0_H5_o(11), SHA256_BLOCK_0_H5_o(10) => 
        SHA256_BLOCK_0_H5_o(10), SHA256_BLOCK_0_H5_o(9) => 
        SHA256_BLOCK_0_H5_o(9), SHA256_BLOCK_0_H5_o(8) => 
        SHA256_BLOCK_0_H5_o(8), SHA256_BLOCK_0_H5_o(7) => 
        SHA256_BLOCK_0_H5_o(7), SHA256_BLOCK_0_H5_o(6) => 
        SHA256_BLOCK_0_H5_o(6), SHA256_BLOCK_0_H5_o(5) => 
        SHA256_BLOCK_0_H5_o(5), SHA256_BLOCK_0_H5_o(4) => 
        SHA256_BLOCK_0_H5_o(4), SHA256_BLOCK_0_H5_o(3) => 
        SHA256_BLOCK_0_H5_o(3), SHA256_BLOCK_0_H5_o(2) => 
        SHA256_BLOCK_0_H5_o(2), SHA256_BLOCK_0_H5_o(1) => 
        SHA256_BLOCK_0_H5_o(1), SHA256_BLOCK_0_H5_o(0) => 
        SHA256_BLOCK_0_H5_o(0), SHA256_BLOCK_0_H6_o(31) => 
        SHA256_BLOCK_0_H6_o(31), SHA256_BLOCK_0_H6_o(30) => 
        SHA256_BLOCK_0_H6_o(30), SHA256_BLOCK_0_H6_o(29) => 
        SHA256_BLOCK_0_H6_o(29), SHA256_BLOCK_0_H6_o(28) => 
        SHA256_BLOCK_0_H6_o(28), SHA256_BLOCK_0_H6_o(27) => 
        SHA256_BLOCK_0_H6_o(27), SHA256_BLOCK_0_H6_o(26) => 
        SHA256_BLOCK_0_H6_o(26), SHA256_BLOCK_0_H6_o(25) => 
        SHA256_BLOCK_0_H6_o(25), SHA256_BLOCK_0_H6_o(24) => 
        SHA256_BLOCK_0_H6_o(24), SHA256_BLOCK_0_H6_o(23) => 
        SHA256_BLOCK_0_H6_o(23), SHA256_BLOCK_0_H6_o(22) => 
        SHA256_BLOCK_0_H6_o(22), SHA256_BLOCK_0_H6_o(21) => 
        SHA256_BLOCK_0_H6_o(21), SHA256_BLOCK_0_H6_o(20) => 
        SHA256_BLOCK_0_H6_o(20), SHA256_BLOCK_0_H6_o(19) => 
        SHA256_BLOCK_0_H6_o(19), SHA256_BLOCK_0_H6_o(18) => 
        SHA256_BLOCK_0_H6_o(18), SHA256_BLOCK_0_H6_o(17) => 
        SHA256_BLOCK_0_H6_o(17), SHA256_BLOCK_0_H6_o(16) => 
        SHA256_BLOCK_0_H6_o(16), SHA256_BLOCK_0_H6_o(15) => 
        SHA256_BLOCK_0_H6_o(15), SHA256_BLOCK_0_H6_o(14) => 
        SHA256_BLOCK_0_H6_o(14), SHA256_BLOCK_0_H6_o(13) => 
        SHA256_BLOCK_0_H6_o(13), SHA256_BLOCK_0_H6_o(12) => 
        SHA256_BLOCK_0_H6_o(12), SHA256_BLOCK_0_H6_o(11) => 
        SHA256_BLOCK_0_H6_o(11), SHA256_BLOCK_0_H6_o(10) => 
        SHA256_BLOCK_0_H6_o(10), SHA256_BLOCK_0_H6_o(9) => 
        SHA256_BLOCK_0_H6_o(9), SHA256_BLOCK_0_H6_o(8) => 
        SHA256_BLOCK_0_H6_o(8), SHA256_BLOCK_0_H6_o(7) => 
        SHA256_BLOCK_0_H6_o(7), SHA256_BLOCK_0_H6_o(6) => 
        SHA256_BLOCK_0_H6_o(6), SHA256_BLOCK_0_H6_o(5) => 
        SHA256_BLOCK_0_H6_o(5), SHA256_BLOCK_0_H6_o(4) => 
        SHA256_BLOCK_0_H6_o(4), SHA256_BLOCK_0_H6_o(3) => 
        SHA256_BLOCK_0_H6_o(3), SHA256_BLOCK_0_H6_o(2) => 
        SHA256_BLOCK_0_H6_o(2), SHA256_BLOCK_0_H6_o(1) => 
        SHA256_BLOCK_0_H6_o(1), SHA256_BLOCK_0_H6_o(0) => 
        SHA256_BLOCK_0_H6_o(0), N6_data(31) => \N6_data[31]\, 
        N6_data(30) => \N6_data[30]\, N6_data(29) => 
        \N6_data[29]\, N6_data(28) => \N6_data[28]\, N6_data(27)
         => \N6_data[27]\, N6_data(26) => \N6_data[26]\, 
        N6_data(25) => \N6_data[25]\, N6_data(24) => 
        \N6_data[24]\, N6_data(23) => \N6_data[23]\, N6_data(22)
         => \N6_data[22]\, N6_data(21) => \N6_data[21]\, 
        N6_data(20) => \N6_data[20]\, N6_data(19) => 
        \N6_data[19]\, N6_data(18) => \N6_data[18]\, N6_data(17)
         => \N6_data[17]\, N6_data(16) => \N6_data[16]\, 
        N6_data(15) => \N6_data[15]\, N6_data(14) => 
        \N6_data[14]\, N6_data(13) => \N6_data[13]\, N6_data(12)
         => \N6_data[12]\, N6_data(11) => \N6_data[11]\, 
        N6_data(10) => \N6_data[10]\, N6_data(9) => \N6_data[9]\, 
        N6_data(8) => \N6_data[8]\, N6_data(7) => \N6_data[7]\, 
        N6_data(6) => \N6_data[6]\, N6_data(5) => \N6_data[5]\, 
        N6_data(4) => \N6_data[4]\, N6_data(3) => \N6_data[3]\, 
        N6_data(2) => \N6_data[2]\, N6_data(1) => \N6_data[1]\, 
        SHA256_BLOCK_0_H7_o(31) => SHA256_BLOCK_0_H7_o(31), 
        SHA256_BLOCK_0_H7_o(30) => SHA256_BLOCK_0_H7_o(30), 
        SHA256_BLOCK_0_H7_o(29) => SHA256_BLOCK_0_H7_o(29), 
        SHA256_BLOCK_0_H7_o(28) => SHA256_BLOCK_0_H7_o(28), 
        SHA256_BLOCK_0_H7_o(27) => SHA256_BLOCK_0_H7_o(27), 
        SHA256_BLOCK_0_H7_o(26) => SHA256_BLOCK_0_H7_o(26), 
        SHA256_BLOCK_0_H7_o(25) => SHA256_BLOCK_0_H7_o(25), 
        SHA256_BLOCK_0_H7_o(24) => SHA256_BLOCK_0_H7_o(24), 
        SHA256_BLOCK_0_H7_o(23) => SHA256_BLOCK_0_H7_o(23), 
        SHA256_BLOCK_0_H7_o(22) => SHA256_BLOCK_0_H7_o(22), 
        SHA256_BLOCK_0_H7_o(21) => SHA256_BLOCK_0_H7_o(21), 
        SHA256_BLOCK_0_H7_o(20) => SHA256_BLOCK_0_H7_o(20), 
        SHA256_BLOCK_0_H7_o(19) => SHA256_BLOCK_0_H7_o(19), 
        SHA256_BLOCK_0_H7_o(18) => SHA256_BLOCK_0_H7_o(18), 
        SHA256_BLOCK_0_H7_o(17) => SHA256_BLOCK_0_H7_o(17), 
        SHA256_BLOCK_0_H7_o(16) => SHA256_BLOCK_0_H7_o(16), 
        SHA256_BLOCK_0_H7_o(15) => SHA256_BLOCK_0_H7_o(15), 
        SHA256_BLOCK_0_H7_o(14) => SHA256_BLOCK_0_H7_o(14), 
        SHA256_BLOCK_0_H7_o(13) => SHA256_BLOCK_0_H7_o(13), 
        SHA256_BLOCK_0_H7_o(12) => SHA256_BLOCK_0_H7_o(12), 
        SHA256_BLOCK_0_H7_o(11) => SHA256_BLOCK_0_H7_o(11), 
        SHA256_BLOCK_0_H7_o(10) => SHA256_BLOCK_0_H7_o(10), 
        SHA256_BLOCK_0_H7_o(9) => SHA256_BLOCK_0_H7_o(9), 
        SHA256_BLOCK_0_H7_o(8) => SHA256_BLOCK_0_H7_o(8), 
        SHA256_BLOCK_0_H7_o(7) => SHA256_BLOCK_0_H7_o(7), 
        SHA256_BLOCK_0_H7_o(6) => SHA256_BLOCK_0_H7_o(6), 
        SHA256_BLOCK_0_H7_o(5) => SHA256_BLOCK_0_H7_o(5), 
        SHA256_BLOCK_0_H7_o(4) => SHA256_BLOCK_0_H7_o(4), 
        SHA256_BLOCK_0_H7_o(3) => SHA256_BLOCK_0_H7_o(3), 
        SHA256_BLOCK_0_H7_o(2) => SHA256_BLOCK_0_H7_o(2), 
        SHA256_BLOCK_0_H7_o(1) => SHA256_BLOCK_0_H7_o(1), 
        SHA256_BLOCK_0_H7_o(0) => SHA256_BLOCK_0_H7_o(0), 
        N7_data(31) => \N7_data[31]\, N7_data(30) => 
        \N7_data[30]\, N7_data(29) => \N7_data[29]\, N7_data(28)
         => \N7_data[28]\, N7_data(27) => \N7_data[27]\, 
        N7_data(26) => \N7_data[26]\, N7_data(25) => 
        \N7_data[25]\, N7_data(24) => \N7_data[24]\, N7_data(23)
         => \N7_data[23]\, N7_data(22) => \N7_data[22]\, 
        N7_data(21) => \N7_data[21]\, N7_data(20) => 
        \N7_data[20]\, N7_data(19) => \N7_data[19]\, N7_data(18)
         => \N7_data[18]\, N7_data(17) => \N7_data[17]\, 
        N7_data(16) => \N7_data[16]\, N7_data(15) => 
        \N7_data[15]\, N7_data(14) => \N7_data[14]\, N7_data(13)
         => \N7_data[13]\, N7_data(12) => \N7_data[12]\, 
        N7_data(11) => \N7_data[11]\, N7_data(10) => 
        \N7_data[10]\, N7_data(9) => \N7_data[9]\, N7_data(8) => 
        \N7_data[8]\, N7_data(7) => \N7_data[7]\, N7_data(6) => 
        \N7_data[6]\, N7_data(5) => \N7_data[5]\, N7_data(4) => 
        \N7_data[4]\, N7_data(3) => \N7_data[3]\, N7_data(2) => 
        \N7_data[2]\, N7_data(1) => \N7_data[1]\, 
        hash_control_st_reg_i(6) => \hash_control_st_reg_i[6]\, 
        R0_data(31) => \R0_data[31]\, R0_data(30) => 
        \R0_data[30]\, R0_data(29) => \R0_data[29]\, R0_data(28)
         => \R0_data[28]\, R0_data(27) => \R0_data[27]\, 
        R0_data(26) => \R0_data[26]\, R0_data(25) => 
        \R0_data[25]\, R0_data(24) => \R0_data[24]\, R0_data(23)
         => \R0_data[23]\, R0_data(22) => \R0_data[22]\, 
        R0_data(21) => \R0_data[21]\, R0_data(20) => 
        \R0_data[20]\, R0_data(19) => \R0_data[19]\, R0_data(18)
         => \R0_data[18]\, R0_data(17) => \R0_data[17]\, 
        R0_data(16) => \R0_data[16]\, R0_data(15) => 
        \R0_data[15]\, R0_data(14) => \R0_data[14]\, R0_data(13)
         => \R0_data[13]\, R0_data(12) => \R0_data[12]\, 
        R0_data(11) => \R0_data[11]\, R0_data(10) => 
        \R0_data[10]\, R0_data(9) => \R0_data[9]\, R0_data(8) => 
        \R0_data[8]\, R0_data(7) => \R0_data[7]\, R0_data(6) => 
        \R0_data[6]\, R0_data(5) => \R0_data[5]\, R0_data(4) => 
        \R0_data[4]\, R0_data(3) => \R0_data[3]\, R0_data(2) => 
        \R0_data[2]\, R0_data(1) => \R0_data[1]\, R0_data(0) => 
        \R0_data[0]\, R1_data(31) => \R1_data[31]\, R1_data(30)
         => \R1_data[30]\, R1_data(29) => \R1_data[29]\, 
        R1_data(28) => \R1_data[28]\, R1_data(27) => 
        \R1_data[27]\, R1_data(26) => \R1_data[26]\, R1_data(25)
         => \R1_data[25]\, R1_data(24) => \R1_data[24]\, 
        R1_data(23) => \R1_data[23]\, R1_data(22) => 
        \R1_data[22]\, R1_data(21) => \R1_data[21]\, R1_data(20)
         => \R1_data[20]\, R1_data(19) => \R1_data[19]\, 
        R1_data(18) => \R1_data[18]\, R1_data(17) => 
        \R1_data[17]\, R1_data(16) => \R1_data[16]\, R1_data(15)
         => \R1_data[15]\, R1_data(14) => \R1_data[14]\, 
        R1_data(13) => \R1_data[13]\, R1_data(12) => 
        \R1_data[12]\, R1_data(11) => \R1_data[11]\, R1_data(10)
         => \R1_data[10]\, R1_data(9) => \R1_data[9]\, R1_data(8)
         => \R1_data[8]\, R1_data(7) => \R1_data[7]\, R1_data(6)
         => \R1_data[6]\, R1_data(5) => \R1_data[5]\, R1_data(4)
         => \R1_data[4]\, R1_data(3) => \R1_data[3]\, R1_data(2)
         => \R1_data[2]\, R1_data(1) => \R1_data[1]\, R1_data(0)
         => \R1_data[0]\, R2_data(31) => \R2_data[31]\, 
        R2_data(30) => \R2_data[30]\, R2_data(29) => 
        \R2_data[29]\, R2_data(28) => \R2_data[28]\, R2_data(27)
         => \R2_data[27]\, R2_data(26) => \R2_data[26]\, 
        R2_data(25) => \R2_data[25]\, R2_data(24) => 
        \R2_data[24]\, R2_data(23) => \R2_data[23]\, R2_data(22)
         => \R2_data[22]\, R2_data(21) => \R2_data[21]\, 
        R2_data(20) => \R2_data[20]\, R2_data(19) => 
        \R2_data[19]\, R2_data(18) => \R2_data[18]\, R2_data(17)
         => \R2_data[17]\, R2_data(16) => \R2_data[16]\, 
        R2_data(15) => \R2_data[15]\, R2_data(14) => 
        \R2_data[14]\, R2_data(13) => \R2_data[13]\, R2_data(12)
         => \R2_data[12]\, R2_data(11) => \R2_data[11]\, 
        R2_data(10) => \R2_data[10]\, R2_data(9) => \R2_data[9]\, 
        R2_data(8) => \R2_data[8]\, R2_data(7) => \R2_data[7]\, 
        R2_data(6) => \R2_data[6]\, R2_data(5) => \R2_data[5]\, 
        R2_data(4) => \R2_data[4]\, R2_data(3) => \R2_data[3]\, 
        R2_data(2) => \R2_data[2]\, R2_data(1) => \R2_data[1]\, 
        R2_data(0) => \R2_data[0]\, R3_data(31) => \R3_data[31]\, 
        R3_data(30) => \R3_data[30]\, R3_data(29) => 
        \R3_data[29]\, R3_data(28) => \R3_data[28]\, R3_data(27)
         => \R3_data[27]\, R3_data(26) => \R3_data[26]\, 
        R3_data(25) => \R3_data[25]\, R3_data(24) => 
        \R3_data[24]\, R3_data(23) => \R3_data[23]\, R3_data(22)
         => \R3_data[22]\, R3_data(21) => \R3_data[21]\, 
        R3_data(20) => \R3_data[20]\, R3_data(19) => 
        \R3_data[19]\, R3_data(18) => \R3_data[18]\, R3_data(17)
         => \R3_data[17]\, R3_data(16) => \R3_data[16]\, 
        R3_data(15) => \R3_data[15]\, R3_data(14) => 
        \R3_data[14]\, R3_data(13) => \R3_data[13]\, R3_data(12)
         => \R3_data[12]\, R3_data(11) => \R3_data[11]\, 
        R3_data(10) => \R3_data[10]\, R3_data(9) => \R3_data[9]\, 
        R3_data(8) => \R3_data[8]\, R3_data(7) => \R3_data[7]\, 
        R3_data(6) => \R3_data[6]\, R3_data(5) => \R3_data[5]\, 
        R3_data(4) => \R3_data[4]\, R3_data(3) => \R3_data[3]\, 
        R3_data(2) => \R3_data[2]\, R3_data(1) => \R3_data[1]\, 
        R3_data(0) => \R3_data[0]\, R4_data(31) => \R4_data[31]\, 
        R4_data(30) => \R4_data[30]\, R4_data(29) => 
        \R4_data[29]\, R4_data(28) => \R4_data[28]\, R4_data(27)
         => \R4_data[27]\, R4_data(26) => \R4_data[26]\, 
        R4_data(25) => \R4_data[25]\, R4_data(24) => 
        \R4_data[24]\, R4_data(23) => \R4_data[23]\, R4_data(22)
         => \R4_data[22]\, R4_data(21) => \R4_data[21]\, 
        R4_data(20) => \R4_data[20]\, R4_data(19) => 
        \R4_data[19]\, R4_data(18) => \R4_data[18]\, R4_data(17)
         => \R4_data[17]\, R4_data(16) => \R4_data[16]\, 
        R4_data(15) => \R4_data[15]\, R4_data(14) => 
        \R4_data[14]\, R4_data(13) => \R4_data[13]\, R4_data(12)
         => \R4_data[12]\, R4_data(11) => \R4_data[11]\, 
        R4_data(10) => \R4_data[10]\, R4_data(9) => \R4_data[9]\, 
        R4_data(8) => \R4_data[8]\, R4_data(7) => \R4_data[7]\, 
        R4_data(6) => \R4_data[6]\, R4_data(5) => \R4_data[5]\, 
        R4_data(4) => \R4_data[4]\, R4_data(3) => \R4_data[3]\, 
        R4_data(2) => \R4_data[2]\, R4_data(1) => \R4_data[1]\, 
        R4_data(0) => \R4_data[0]\, R5_data(31) => \R5_data[31]\, 
        R5_data(30) => \R5_data[30]\, R5_data(29) => 
        \R5_data[29]\, R5_data(28) => \R5_data[28]\, R5_data(27)
         => \R5_data[27]\, R5_data(26) => \R5_data[26]\, 
        R5_data(25) => \R5_data[25]\, R5_data(24) => 
        \R5_data[24]\, R5_data(23) => \R5_data[23]\, R5_data(22)
         => \R5_data[22]\, R5_data(21) => \R5_data[21]\, 
        R5_data(20) => \R5_data[20]\, R5_data(19) => 
        \R5_data[19]\, R5_data(18) => \R5_data[18]\, R5_data(17)
         => \R5_data[17]\, R5_data(16) => \R5_data[16]\, 
        R5_data(15) => \R5_data[15]\, R5_data(14) => 
        \R5_data[14]\, R5_data(13) => \R5_data[13]\, R5_data(12)
         => \R5_data[12]\, R5_data(11) => \R5_data[11]\, 
        R5_data(10) => \R5_data[10]\, R5_data(9) => \R5_data[9]\, 
        R5_data(8) => \R5_data[8]\, R5_data(7) => \R5_data[7]\, 
        R5_data(6) => \R5_data[6]\, R5_data(5) => \R5_data[5]\, 
        R5_data(4) => \R5_data[4]\, R5_data(3) => \R5_data[3]\, 
        R5_data(2) => \R5_data[2]\, R5_data(1) => \R5_data[1]\, 
        R5_data(0) => \R5_data[0]\, R6_data(31) => \R6_data[31]\, 
        R6_data(30) => \R6_data[30]\, R6_data(29) => 
        \R6_data[29]\, R6_data(28) => \R6_data[28]\, R6_data(27)
         => \R6_data[27]\, R6_data(26) => \R6_data[26]\, 
        R6_data(25) => \R6_data[25]\, R6_data(24) => 
        \R6_data[24]\, R6_data(23) => \R6_data[23]\, R6_data(22)
         => \R6_data[22]\, R6_data(21) => \R6_data[21]\, 
        R6_data(20) => \R6_data[20]\, R6_data(19) => 
        \R6_data[19]\, R6_data(18) => \R6_data[18]\, R6_data(17)
         => \R6_data[17]\, R6_data(16) => \R6_data[16]\, 
        R6_data(15) => \R6_data[15]\, R6_data(14) => 
        \R6_data[14]\, R6_data(13) => \R6_data[13]\, R6_data(12)
         => \R6_data[12]\, R6_data(11) => \R6_data[11]\, 
        R6_data(10) => \R6_data[10]\, R6_data(9) => \R6_data[9]\, 
        R6_data(8) => \R6_data[8]\, R6_data(7) => \R6_data[7]\, 
        R6_data(6) => \R6_data[6]\, R6_data(5) => \R6_data[5]\, 
        R6_data(4) => \R6_data[4]\, R6_data(3) => \R6_data[3]\, 
        R6_data(2) => \R6_data[2]\, R6_data(1) => \R6_data[1]\, 
        R6_data(0) => \R6_data[0]\, R7_data(31) => \R7_data[31]\, 
        R7_data(30) => \R7_data[30]\, R7_data(29) => 
        \R7_data[29]\, R7_data(28) => \R7_data[28]\, R7_data(27)
         => \R7_data[27]\, R7_data(26) => \R7_data[26]\, 
        R7_data(25) => \R7_data[25]\, R7_data(24) => 
        \R7_data[24]\, R7_data(23) => \R7_data[23]\, R7_data(22)
         => \R7_data[22]\, R7_data(21) => \R7_data[21]\, 
        R7_data(20) => \R7_data[20]\, R7_data(19) => 
        \R7_data[19]\, R7_data(18) => \R7_data[18]\, R7_data(17)
         => \R7_data[17]\, R7_data(16) => \R7_data[16]\, 
        R7_data(15) => \R7_data[15]\, R7_data(14) => 
        \R7_data[14]\, R7_data(13) => \R7_data[13]\, R7_data(12)
         => \R7_data[12]\, R7_data(11) => \R7_data[11]\, 
        R7_data(10) => \R7_data[10]\, R7_data(9) => \R7_data[9]\, 
        R7_data(8) => \R7_data[8]\, R7_data(7) => \R7_data[7]\, 
        R7_data(6) => \R7_data[6]\, R7_data(5) => \R7_data[5]\, 
        R7_data(4) => \R7_data[4]\, R7_data(3) => \R7_data[3]\, 
        R7_data(2) => \R7_data[2]\, R7_data(1) => \R7_data[1]\, 
        R7_data(0) => \R7_data[0]\, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, N_168_i_0 => 
        N_168_i_0, next_reg_H0_cry_0_0_Y => next_reg_H0_cry_0_0_Y, 
        next_reg_H1_cry_0_0_Y => next_reg_H1_cry_0_0_Y, 
        next_reg_H2_cry_0_0_Y => next_reg_H2_cry_0_0_Y, 
        next_reg_H3_cry_0_0_Y => next_reg_H3_cry_0_0_Y, 
        next_reg_H4_cry_0_0_Y => next_reg_H4_cry_0_0_Y, 
        next_reg_H5_cry_0_0_Y => next_reg_H5_cry_0_0_Y, 
        next_reg_H6_cry_0_0_Y => next_reg_H6_cry_0_0_Y, 
        next_reg_H7_cry_0_0_Y => next_reg_H7_cry_0_0_Y);
    
    Inst_sha256_padding : sha256_padding
      port map(di_o_0(1) => di_o_0(1), 
        reg_17x32_0_valid_bytes_0(1) => 
        reg_17x32_0_valid_bytes_0(1), 
        reg_17x32_0_valid_bytes_0(0) => 
        reg_17x32_0_valid_bytes_0(0), Kt_addr_fast(0) => 
        \Kt_addr_fast[0]\, hash_control_st_reg(2) => 
        \hash_control_st_reg[2]\, W_out_2_0(5) => \W_out_2_0[5]\, 
        W_out_i_i_2(31) => \W_out_i_i_2[31]\, W_out_i_i_1(31) => 
        \W_out_i_i_1[31]\, W_out_i_1(1) => \W_out_i_1[1]\, 
        W_out_i_1(0) => \W_out_i_1[0]\, W_out_i_0(2) => 
        \W_out_i_0[2]\, msg_bitlen(63) => \msg_bitlen[63]\, 
        msg_bitlen(62) => \msg_bitlen[62]\, msg_bitlen(61) => 
        \msg_bitlen[61]\, msg_bitlen(60) => \msg_bitlen[60]\, 
        msg_bitlen(59) => \msg_bitlen[59]\, msg_bitlen(58) => 
        \msg_bitlen[58]\, msg_bitlen(57) => \msg_bitlen[57]\, 
        msg_bitlen(56) => \msg_bitlen[56]\, msg_bitlen(55) => 
        \msg_bitlen[55]\, msg_bitlen(54) => \msg_bitlen[54]\, 
        msg_bitlen(53) => \msg_bitlen[53]\, msg_bitlen(52) => 
        \msg_bitlen[52]\, msg_bitlen(51) => \msg_bitlen[51]\, 
        msg_bitlen(50) => \msg_bitlen[50]\, msg_bitlen(49) => 
        \msg_bitlen[49]\, msg_bitlen(48) => \msg_bitlen[48]\, 
        msg_bitlen(47) => \msg_bitlen[47]\, msg_bitlen(46) => 
        \msg_bitlen[46]\, msg_bitlen(45) => \msg_bitlen[45]\, 
        msg_bitlen(44) => \msg_bitlen[44]\, msg_bitlen(43) => 
        \msg_bitlen[43]\, msg_bitlen(42) => \msg_bitlen[42]\, 
        msg_bitlen(41) => \msg_bitlen[41]\, msg_bitlen(40) => 
        \msg_bitlen[40]\, msg_bitlen(39) => \msg_bitlen[39]\, 
        msg_bitlen(38) => \msg_bitlen[38]\, msg_bitlen(37) => 
        \msg_bitlen[37]\, msg_bitlen(36) => \msg_bitlen[36]\, 
        msg_bitlen(35) => \msg_bitlen[35]\, msg_bitlen(34) => 
        \msg_bitlen[34]\, msg_bitlen(33) => \msg_bitlen[33]\, 
        msg_bitlen(32) => \msg_bitlen[32]\, msg_bitlen(31) => 
        \msg_bitlen[31]\, msg_bitlen(30) => \msg_bitlen[30]\, 
        msg_bitlen(29) => \msg_bitlen[29]\, msg_bitlen(28) => 
        \msg_bitlen[28]\, msg_bitlen(27) => \msg_bitlen[27]\, 
        msg_bitlen(26) => \msg_bitlen[26]\, msg_bitlen(25) => 
        \msg_bitlen[25]\, msg_bitlen(24) => \msg_bitlen[24]\, 
        msg_bitlen(23) => \msg_bitlen[23]\, msg_bitlen(22) => 
        \msg_bitlen[22]\, msg_bitlen(21) => \msg_bitlen[21]\, 
        msg_bitlen(20) => \msg_bitlen[20]\, msg_bitlen(19) => 
        \msg_bitlen[19]\, msg_bitlen(18) => \msg_bitlen[18]\, 
        msg_bitlen(17) => \msg_bitlen[17]\, msg_bitlen(16) => 
        \msg_bitlen[16]\, msg_bitlen(15) => \msg_bitlen[15]\, 
        msg_bitlen(14) => \msg_bitlen[14]\, msg_bitlen(13) => 
        \msg_bitlen[13]\, msg_bitlen(12) => \msg_bitlen[12]\, 
        msg_bitlen(11) => \msg_bitlen[11]\, msg_bitlen(10) => 
        \msg_bitlen[10]\, msg_bitlen(9) => \msg_bitlen[9]\, 
        msg_bitlen(8) => \msg_bitlen[8]\, msg_bitlen(7) => 
        \msg_bitlen[7]\, msg_bitlen(6) => \msg_bitlen[6]\, 
        msg_bitlen(5) => \msg_bitlen[5]\, msg_bitlen(4) => 
        \msg_bitlen[4]\, msg_bitlen(3) => \msg_bitlen[3]\, 
        state_2 => state_2, state_0 => state_0, state_3 => 
        state_3, Kt_addr_5 => \Kt_addr[5]\, Kt_addr_0 => 
        \Kt_addr[0]\, W_out_2_0_0_1 => \W_out_2_0_0[4]\, 
        W_out_2_0_0_0 => \W_out_2_0_0[3]\, W_out_2_0_0_3 => 
        \W_out_2_0_0[6]\, W_out_2_0_1_8 => \W_out_2_0_1[15]\, 
        W_out_2_0_1_0 => \W_out_2_0_1[7]\, W_out_2_i_0_18 => 
        \W_out_2_i_0[26]\, W_out_2_i_0_21 => \W_out_2_i_0[29]\, 
        W_out_2_i_0_17 => \W_out_2_i_0[25]\, W_out_2_i_0_22 => 
        \W_out_2_i_0[30]\, W_out_2_i_0_20 => \W_out_2_i_0[28]\, 
        W_out_2_i_0_16 => \W_out_2_i_0[24]\, W_out_2_i_0_19 => 
        \W_out_2_i_0[27]\, W_out_2_0_2_0 => \W_out_2_0_2[15]\, 
        W_out_2_0_2_8 => \W_out_2_0_2[23]\, 
        sha256_controller_0_di_o_3 => sha256_controller_0_di_o_3, 
        sha256_controller_0_di_o_5 => sha256_controller_0_di_o_5, 
        sha256_controller_0_di_o_0 => sha256_controller_0_di_o_0, 
        W_out_2_i_1_18 => \W_out_2_i_1[26]\, W_out_2_i_1_21 => 
        \W_out_2_i_1[29]\, W_out_2_i_1_17 => \W_out_2_i_1[25]\, 
        W_out_2_i_1_22 => \W_out_2_i_1[30]\, W_out_2_i_1_20 => 
        \W_out_2_i_1[28]\, W_out_2_i_1_16 => \W_out_2_i_1[24]\, 
        W_out_2_i_1_19 => \W_out_2_i_1[27]\, W_out_2_i_1_12 => 
        \W_out_2_i_1[20]\, W_out_2_i_1_8 => \W_out_2_i_1[16]\, 
        W_out_2_i_1_10 => \W_out_2_i_1[18]\, W_out_2_i_1_13 => 
        \W_out_2_i_1[21]\, W_out_2_i_1_14 => \W_out_2_i_1[22]\, 
        W_out_2_i_1_11 => \W_out_2_i_1[19]\, W_out_2_i_1_9 => 
        \W_out_2_i_1[17]\, W_out_2_i_1_1 => \W_out_2_i_1[9]\, 
        W_out_2_i_1_2 => \W_out_2_i_1[10]\, W_out_2_i_1_0 => 
        \W_out_2_i_1[8]\, W_out_2_i_1_4 => \W_out_2_i_1[12]\, 
        W_out_2_i_1_3 => \W_out_2_i_1[11]\, W_out_2_i_1_6 => 
        \W_out_2_i_1[14]\, W_out_2_i_1_5 => \W_out_2_i_1[13]\, 
        N_223 => N_223, N_1702 => N_1702, N_1710 => N_1710, 
        SHA256_Module_0_di_req_o => \SHA256_Module_0_di_req_o\, 
        N_388 => N_388, N_112 => N_112, one_insert => one_insert, 
        Kt_addr_0_rep2 => Kt_addr_0_rep2, sha_last_blk_reg => 
        sha_last_blk_reg, Kt_addr_4_rep1 => Kt_addr_4_rep1, 
        bytes_sel => bytes_sel, ren_pos => ren_pos, N_102 => 
        N_102, sha_last_blk_next_0_o2_2_out_0 => 
        sha_last_blk_next_0_o2_2_out_0, N_361 => N_361, 
        SHA256_Module_0_data_available_lastbank_8 => 
        SHA256_Module_0_data_available_lastbank_8, N_111 => N_111, 
        N_1690 => N_1690, N_245 => N_245, N_1691 => N_1691, N_248
         => N_248, N_1693 => N_1693, N_251 => N_251, N_1692 => 
        N_1692, N_349 => N_349, N_1718 => N_1718, N_1694 => 
        N_1694, N_255 => N_255, N_1698 => N_1698, N_1701 => 
        N_1701, N_98 => N_98, N_307 => N_307, N_1696 => N_1696, 
        N_1697 => N_1697, N_1695 => N_1695, N_1699 => N_1699, 
        N_1707 => N_1707, N_1708 => N_1708, N_1709 => N_1709, 
        N_1706 => N_1706, N_1704 => N_1704, N_1688 => N_1688, 
        N_1687 => N_1687, N_1689 => N_1689, N_1713 => N_1713, 
        N_1716 => N_1716, N_1712 => N_1712, N_1717 => N_1717, 
        N_1715 => N_1715, N_1711 => N_1711, N_1714 => N_1714, 
        N_273 => N_273, N_266 => N_266, N_263 => N_263, N_260 => 
        N_260, N_287 => N_287, N_290 => N_290, N_293 => N_293, 
        N_296 => N_296, N_299 => N_299, N_302 => N_302, N_305 => 
        N_305, N_268 => N_268, N_275 => N_275, N_278 => N_278);
    
    Inst_sha256_msg_sch : sha256_msg_sch
      port map(Wt_data(31) => \Wt_data[31]\, Wt_data(30) => 
        \Wt_data[30]\, Wt_data(29) => \Wt_data[29]\, Wt_data(28)
         => \Wt_data[28]\, Wt_data(27) => \Wt_data[27]\, 
        Wt_data(26) => \Wt_data[26]\, Wt_data(25) => 
        \Wt_data[25]\, Wt_data(24) => \Wt_data[24]\, Wt_data(23)
         => \Wt_data[23]\, Wt_data(22) => \Wt_data[22]\, 
        Wt_data(21) => \Wt_data[21]\, Wt_data(20) => 
        \Wt_data[20]\, Wt_data(19) => \Wt_data[19]\, Wt_data(18)
         => \Wt_data[18]\, Wt_data(17) => \Wt_data[17]\, 
        Wt_data(16) => \Wt_data[16]\, Wt_data(15) => 
        \Wt_data[15]\, Wt_data(14) => \Wt_data[14]\, Wt_data(13)
         => \Wt_data[13]\, Wt_data(12) => \Wt_data[12]\, 
        Wt_data(11) => \Wt_data[11]\, Wt_data(10) => 
        \Wt_data[10]\, Wt_data(9) => \Wt_data[9]\, Wt_data(8) => 
        \Wt_data[8]\, Wt_data(7) => \Wt_data[7]\, Wt_data(6) => 
        \Wt_data[6]\, Wt_data(5) => \Wt_data[5]\, Wt_data(4) => 
        \Wt_data[4]\, Wt_data(3) => \Wt_data[3]\, Wt_data(2) => 
        \Wt_data[2]\, Wt_data(1) => \Wt_data[1]\, Wt_data(0) => 
        \Wt_data[0]\, W_out_2_0(5) => \W_out_2_0[5]\, 
        W_out_i_i_2(31) => \W_out_i_i_2[31]\, W_out_i_i_1(31) => 
        \W_out_i_i_1[31]\, W_out_2_i_0(30) => \W_out_2_i_0[30]\, 
        W_out_2_i_0(29) => \W_out_2_i_0[29]\, W_out_2_i_0(28) => 
        \W_out_2_i_0[28]\, W_out_2_i_0(27) => \W_out_2_i_0[27]\, 
        W_out_2_i_0(26) => \W_out_2_i_0[26]\, W_out_2_i_0(25) => 
        \W_out_2_i_0[25]\, W_out_2_i_0(24) => \W_out_2_i_0[24]\, 
        W_out_i_0(2) => \W_out_i_0[2]\, W_out_i_1(1) => 
        \W_out_i_1[1]\, W_out_i_1(0) => \W_out_i_1[0]\, 
        W_out_2_0_0_3 => \W_out_2_0_0[6]\, W_out_2_0_0_1 => 
        \W_out_2_0_0[4]\, W_out_2_0_0_0 => \W_out_2_0_0[3]\, 
        W_out_2_0_2_8 => \W_out_2_0_2[23]\, W_out_2_0_2_0 => 
        \W_out_2_0_2[15]\, W_out_2_0_1_0 => \W_out_2_0_1[7]\, 
        W_out_2_0_1_8 => \W_out_2_0_1[15]\, W_out_2_i_1_22 => 
        \W_out_2_i_1[30]\, W_out_2_i_1_21 => \W_out_2_i_1[29]\, 
        W_out_2_i_1_20 => \W_out_2_i_1[28]\, W_out_2_i_1_19 => 
        \W_out_2_i_1[27]\, W_out_2_i_1_18 => \W_out_2_i_1[26]\, 
        W_out_2_i_1_17 => \W_out_2_i_1[25]\, W_out_2_i_1_16 => 
        \W_out_2_i_1[24]\, W_out_2_i_1_14 => \W_out_2_i_1[22]\, 
        W_out_2_i_1_13 => \W_out_2_i_1[21]\, W_out_2_i_1_12 => 
        \W_out_2_i_1[20]\, W_out_2_i_1_11 => \W_out_2_i_1[19]\, 
        W_out_2_i_1_10 => \W_out_2_i_1[18]\, W_out_2_i_1_9 => 
        \W_out_2_i_1[17]\, W_out_2_i_1_8 => \W_out_2_i_1[16]\, 
        W_out_2_i_1_6 => \W_out_2_i_1[14]\, W_out_2_i_1_5 => 
        \W_out_2_i_1[13]\, W_out_2_i_1_4 => \W_out_2_i_1[12]\, 
        W_out_2_i_1_3 => \W_out_2_i_1[11]\, W_out_2_i_1_2 => 
        \W_out_2_i_1[10]\, W_out_2_i_1_1 => \W_out_2_i_1[9]\, 
        W_out_2_i_1_0 => \W_out_2_i_1[8]\, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, N_244_i_0 => 
        N_244_i_0, next_r0_0_cry_0_Y => next_r0_0_cry_0_Y, N_251
         => N_251, ld_i_i_3 => ld_i_i_3, N_349 => N_349, N_248
         => N_248, N_245 => N_245, N_255 => N_255, N_98 => N_98, 
        N_307 => N_307, N_305 => N_305, N_302 => N_302, N_299 => 
        N_299, N_296 => N_296, N_293 => N_293, N_290 => N_290, 
        N_287 => N_287, N_278 => N_278, N_275 => N_275, N_273 => 
        N_273, N_268 => N_268, N_266 => N_266, N_263 => N_263, 
        N_260 => N_260);
    
    Inst_sha256_kt_rom : sha256_kt_rom
      port map(hash_control_st_reg_ns_i_0_a2_0(4) => 
        \hash_control_st_reg_ns_i_0_a2_0[4]\, Kt_addr_fast(4) => 
        \Kt_addr_fast[4]\, Kt_addr_fast(3) => \Kt_addr_fast[3]\, 
        Kt_addr_fast(2) => \Kt_addr_fast[2]\, Kt_addr_fast(1) => 
        \Kt_addr_fast[1]\, Kt_addr_fast(0) => \Kt_addr_fast[0]\, 
        hash_control_st_reg_ns_i_0_a2_2(4) => 
        \hash_control_st_reg_ns_i_0_a2_2[4]\, Kt_addr(5) => 
        \Kt_addr[5]\, Kt_addr(4) => \Kt_addr[4]\, Kt_addr(3) => 
        \Kt_addr[3]\, Kt_addr(2) => \Kt_addr[2]\, Kt_addr(1) => 
        \Kt_addr[1]\, Kt_addr(0) => \Kt_addr[0]\, Kt_data_9 => 
        \Kt_data[24]\, Kt_data_0 => \Kt_data[15]\, Kt_addr_3_rep1
         => Kt_addr_3_rep1, m62_am => m62_am, Kt_addr_0_rep1 => 
        Kt_addr_0_rep1, m104_bm => m104_bm, Kt_addr_2_rep1 => 
        Kt_addr_2_rep1, Kt_addr_0_rep2 => Kt_addr_0_rep2, m49_am
         => m49_am, Kt_addr_1_rep1 => Kt_addr_1_rep1, m49_bm => 
        m49_bm, m137_am => m137_am, Kt_addr_3_rep2 => 
        Kt_addr_3_rep2, m137_bm => m137_bm, Kt_addr_4_rep2 => 
        Kt_addr_4_rep2, m215_am => m215_am, Kt_addr_4_rep1 => 
        Kt_addr_4_rep1, m215_bm => m215_bm, Kt_addr_2_rep2 => 
        Kt_addr_2_rep2, m250_am => m250_am, Kt_addr_1_rep2 => 
        Kt_addr_1_rep2, m250_bm => m250_bm, m207_1_1 => m207_1_1, 
        m207_1_0 => m207_1_0, m157 => m157, m197_1_1 => m197_1_1, 
        m197_1_0 => m197_1_0, m95_1_1 => m95_1_1, m95_1_0 => 
        m95_1_0, m325 => m325, m168_1_1 => m168_1_1, m168_1_0 => 
        m168_1_0, m316 => m316, m34 => m34, m114 => m114, m285
         => m285, m289 => m289, m254 => m254, m239 => m239, m124
         => m124, m141 => m141, m304 => m304, m19 => m19, 
        pad_one_reg_0_0_a2_0 => pad_one_reg_0_0_a2_0, m296 => 
        m296, m78 => m78, m219 => m219, m230 => m230, m177 => 
        m177, m73_0 => m73, i3_mux_1 => i3_mux_1, m10_ns => 
        m10_ns, m67_ns => m67_ns, m83_ns => m83_ns, m110_ns => 
        m110_ns, m119_ns => m119_ns, m144_ns => m144_ns, m172_ns
         => m172_ns, m222_ns => m222_ns, m226_ns => m226_ns, 
        m235_ns => m235_ns, m258_ns => m258_ns, m276_ns => 
        m276_ns, m281_ns => m281_ns, m292_ns => m292_ns, m300_ns
         => m300_ns, sha_last_blk_next_0_a4_0 => 
        sha_last_blk_next_0_a4_0, m273 => m273, m104_am => 
        m104_am, m62_bm => m62_bm);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity limiter_1cycle is

    port( prev_sig                             : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          first_block                          : in    std_logic
        );

end limiter_1cycle;

architecture DEF_ARCH of limiter_1cycle is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \prev_sig\ : SLE
      port map(D => first_block, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => prev_sig);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity limiter_1cycle_0 is

    port( prev_sig                             : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          data_out_ready                       : in    std_logic
        );

end limiter_1cycle_0;

architecture DEF_ARCH of limiter_1cycle_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \prev_sig\ : SLE
      port map(D => data_out_ready, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => prev_sig);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_17x32 is

    port( reg_17x32_0_last_word                     : out   std_logic_vector(3 downto 0);
          reg_17x32_0_valid_bytes_0                 : out   std_logic_vector(1 downto 0);
          sha256_controller_0_read_addr_0           : in    std_logic_vector(3 downto 0);
          waddr_in_net_0                            : in    std_logic_vector(4 downto 0);
          data_out_ready                            : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0      : in    std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F       : in    std_logic;
          SHA256_Module_0_data_available            : out   std_logic;
          ren_pos                                   : out   std_logic;
          N_111_i_0                                 : in    std_logic;
          N_109_i_0                                 : in    std_logic;
          N_168_i_0                                 : in    std_logic;
          N_107_i_0                                 : in    std_logic;
          N_99_i_0                                  : in    std_logic;
          N_97_i_0                                  : in    std_logic;
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic;
          N_67_i_0                                  : in    std_logic;
          first_block                               : out   std_logic;
          N_65_i_0                                  : in    std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F_i_0   : in    std_logic;
          N_105_i_0                                 : in    std_logic;
          N_103_i_0                                 : in    std_logic;
          N_158_i_0                                 : in    std_logic;
          N_156_i_0                                 : in    std_logic;
          N_101_i_0                                 : in    std_logic;
          N_152_i_0                                 : in    std_logic;
          N_95_i_0                                  : in    std_logic;
          N_93_i_0                                  : in    std_logic;
          N_91_i_0                                  : in    std_logic;
          N_140_i_0                                 : in    std_logic;
          N_89_i_0                                  : in    std_logic;
          N_87_i_0                                  : in    std_logic;
          N_133_i_0                                 : in    std_logic;
          N_85_i_0                                  : in    std_logic;
          N_83_i_0                                  : in    std_logic;
          N_77_i_0                                  : in    std_logic;
          N_75_i_0                                  : in    std_logic;
          N_73_i_0                                  : in    std_logic;
          N_71_i_0                                  : in    std_logic;
          N_69_i_0                                  : in    std_logic;
          N_116_i_0                                 : in    std_logic;
          N_114_i_0                                 : in    std_logic;
          N_112_i_0                                 : in    std_logic;
          N_110_i_0                                 : in    std_logic;
          N_1687                                    : out   std_logic;
          N_1717                                    : out   std_logic;
          N_1690                                    : out   std_logic;
          N_1689                                    : out   std_logic;
          N_1688                                    : out   std_logic;
          N_1715                                    : out   std_logic;
          N_1713                                    : out   std_logic;
          N_1710                                    : out   std_logic;
          N_1701                                    : out   std_logic;
          N_1714                                    : out   std_logic;
          N_1712                                    : out   std_logic;
          N_1716                                    : out   std_logic;
          N_1700                                    : out   std_logic;
          N_1698                                    : out   std_logic;
          N_1697                                    : out   std_logic;
          N_1692                                    : out   std_logic;
          N_1691                                    : out   std_logic;
          N_1704                                    : out   std_logic;
          N_1694                                    : out   std_logic;
          N_1709                                    : out   std_logic;
          N_1708                                    : out   std_logic;
          N_1707                                    : out   std_logic;
          N_1718                                    : out   std_logic;
          N_1703                                    : out   std_logic;
          N_1696                                    : out   std_logic;
          N_1699                                    : out   std_logic;
          N_1705                                    : out   std_logic;
          N_1695                                    : out   std_logic;
          N_1693                                    : out   std_logic;
          N_1706                                    : out   std_logic;
          N_1702                                    : out   std_logic;
          N_1711                                    : out   std_logic;
          CertificationSystem_sb_0_GPIO_1_M2F       : in    std_logic;
          AHB_slave_dummy_0_write_en                : in    std_logic
        );

end reg_17x32;

architecture DEF_ARCH of reg_17x32 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal data_out_ready_net_1, VCC_net_1, \data_out_ready_1\, 
        GND_net_1, \SHA256_Module_0_data_available\, N_12_0_i_0, 
        data_out_ready_0_sqmuxa, \line8_or[0]_net_1\, line8_0_62, 
        \line7[63]_net_1\, \line7_or[32]_net_1\, 
        \line7[62]_net_1\, \line7[61]_net_1\, \line7[60]_net_1\, 
        \line7[59]_net_1\, \line7[58]_net_1\, \line7[57]_net_1\, 
        \line7[56]_net_1\, \line7[55]_net_1\, \line7[54]_net_1\, 
        \line7[53]_net_1\, \line7[52]_net_1\, \line7[51]_net_1\, 
        \line7[50]_net_1\, \line7[49]_net_1\, \line7[48]_net_1\, 
        \line7[47]_net_1\, \line7[46]_net_1\, \line7[45]_net_1\, 
        \line7[44]_net_1\, \line7[43]_net_1\, \line7[42]_net_1\, 
        \line7[41]_net_1\, \line7[40]_net_1\, \line7[39]_net_1\, 
        \line7[38]_net_1\, \line7[37]_net_1\, \line7[36]_net_1\, 
        \line7[35]_net_1\, \line7[34]_net_1\, \line7[33]_net_1\, 
        \line7[32]_net_1\, line7_0, \line7[31]_net_1\, 
        \line7_or[0]_net_1\, \line7[30]_net_1\, \line7[29]_net_1\, 
        \line7[28]_net_1\, \line7[27]_net_1\, \line7[26]_net_1\, 
        \line7[25]_net_1\, \line7[24]_net_1\, \line7[23]_net_1\, 
        \line7[22]_net_1\, \line7[21]_net_1\, \line7[20]_net_1\, 
        \line7[19]_net_1\, \line7[18]_net_1\, \line7[17]_net_1\, 
        \line7[16]_net_1\, \line7[15]_net_1\, \line7[14]_net_1\, 
        \line7[13]_net_1\, \line7[12]_net_1\, \line7[11]_net_1\, 
        \line7[10]_net_1\, \line7[9]_net_1\, \line7[8]_net_1\, 
        \line7[7]_net_1\, \line7[6]_net_1\, \line7[5]_net_1\, 
        \line7[4]_net_1\, \line7[3]_net_1\, \line7[2]_net_1\, 
        \line7[1]_net_1\, \line7[0]_net_1\, line7_0_62, 
        \line6[63]_net_1\, \line6_or[32]_net_1\, 
        \line6[62]_net_1\, \line6[61]_net_1\, \line6[60]_net_1\, 
        \line6[59]_net_1\, \line6[58]_net_1\, \line6[57]_net_1\, 
        \line6[56]_net_1\, \line6[55]_net_1\, \line6[54]_net_1\, 
        \line6[53]_net_1\, \line6[52]_net_1\, \line6[51]_net_1\, 
        \line6[50]_net_1\, \line6[49]_net_1\, \line6[48]_net_1\, 
        \line6[47]_net_1\, \line6[46]_net_1\, \line6[45]_net_1\, 
        \line6[44]_net_1\, \line6[43]_net_1\, \line6[42]_net_1\, 
        \line6[41]_net_1\, \line6[40]_net_1\, \line6[39]_net_1\, 
        \line6[38]_net_1\, \line6[37]_net_1\, \line6[36]_net_1\, 
        \line6[35]_net_1\, \line6[34]_net_1\, \line6[33]_net_1\, 
        \line6[32]_net_1\, line6_0, \line6[31]_net_1\, 
        \line6_or[0]_net_1\, \line6[30]_net_1\, \line6[29]_net_1\, 
        \line6[28]_net_1\, \line6[27]_net_1\, \line6[26]_net_1\, 
        \line6[25]_net_1\, \line6[24]_net_1\, \line6[23]_net_1\, 
        \line6[22]_net_1\, \line6[21]_net_1\, \line6[20]_net_1\, 
        \line6[19]_net_1\, \line6[18]_net_1\, \line6[17]_net_1\, 
        \line6[16]_net_1\, \line6[15]_net_1\, \line6[14]_net_1\, 
        \line6[13]_net_1\, \line6[12]_net_1\, \line6[11]_net_1\, 
        \line6[10]_net_1\, \line6[9]_net_1\, \line6[8]_net_1\, 
        \line6[7]_net_1\, \line6[6]_net_1\, \line6[5]_net_1\, 
        \line6[4]_net_1\, \line6[3]_net_1\, \line6[2]_net_1\, 
        \line6[1]_net_1\, \line6[0]_net_1\, line6_0_62, 
        \line5[63]_net_1\, \line5_or[32]_net_1\, 
        \line5[62]_net_1\, \line5[61]_net_1\, \line5[60]_net_1\, 
        \line5[59]_net_1\, \line5[58]_net_1\, \line5[57]_net_1\, 
        \line5[56]_net_1\, \line5[55]_net_1\, \line5[54]_net_1\, 
        \line5[53]_net_1\, \line5[52]_net_1\, \line5[51]_net_1\, 
        \line5[50]_net_1\, \line5[49]_net_1\, \line5[48]_net_1\, 
        \line5[47]_net_1\, \line5[46]_net_1\, \line5[45]_net_1\, 
        \line5[44]_net_1\, \line5[43]_net_1\, \line5[42]_net_1\, 
        \line5[41]_net_1\, \line5[40]_net_1\, \line5[39]_net_1\, 
        \line5[38]_net_1\, \line5[37]_net_1\, \line5[36]_net_1\, 
        \line5[35]_net_1\, \line5[34]_net_1\, \line5[33]_net_1\, 
        \line5[32]_net_1\, line5_0, \line5[31]_net_1\, 
        \line5_or[0]_net_1\, \line5[30]_net_1\, \line5[29]_net_1\, 
        \line5[28]_net_1\, \line5[27]_net_1\, \line5[26]_net_1\, 
        \line5[25]_net_1\, \line5[24]_net_1\, \line5[23]_net_1\, 
        \line5[22]_net_1\, \line5[21]_net_1\, \line5[20]_net_1\, 
        \line5[19]_net_1\, \line5[18]_net_1\, \line5[17]_net_1\, 
        \line5[16]_net_1\, \line5[15]_net_1\, \line5[14]_net_1\, 
        \line5[13]_net_1\, \line5[12]_net_1\, \line5[11]_net_1\, 
        \line5[10]_net_1\, \line5[9]_net_1\, \line5[8]_net_1\, 
        \line5[7]_net_1\, \line5[6]_net_1\, \line5[5]_net_1\, 
        \line5[4]_net_1\, \line5[3]_net_1\, \line5[2]_net_1\, 
        \line5[1]_net_1\, \line5[0]_net_1\, line5_0_62, 
        \line4[63]_net_1\, \line4_or[32]_net_1\, 
        \line4[62]_net_1\, \line4[61]_net_1\, \line4[60]_net_1\, 
        \line4[59]_net_1\, \line4[58]_net_1\, \line4[57]_net_1\, 
        \line4[56]_net_1\, \line4[55]_net_1\, \line4[54]_net_1\, 
        \line4[53]_net_1\, \line4[52]_net_1\, \line4[51]_net_1\, 
        \line4[50]_net_1\, \line4[49]_net_1\, \line4[48]_net_1\, 
        \line4[47]_net_1\, \line4[46]_net_1\, \line4[45]_net_1\, 
        \line4[44]_net_1\, \line4[43]_net_1\, \line4[42]_net_1\, 
        \line4[41]_net_1\, \line4[40]_net_1\, \line4[39]_net_1\, 
        \line4[38]_net_1\, \line4[37]_net_1\, \line4[36]_net_1\, 
        \line4[35]_net_1\, \line4[34]_net_1\, \line4[33]_net_1\, 
        \line4[32]_net_1\, line4_0, \line4[31]_net_1\, 
        \line4_or[0]_net_1\, \line4[30]_net_1\, \line4[29]_net_1\, 
        \line4[28]_net_1\, \line4[27]_net_1\, \line4[26]_net_1\, 
        \line4[25]_net_1\, \line4[24]_net_1\, \line4[23]_net_1\, 
        \line4[22]_net_1\, \line4[21]_net_1\, \line4[20]_net_1\, 
        \line4[19]_net_1\, \line4[18]_net_1\, \line4[17]_net_1\, 
        \line4[16]_net_1\, \line4[15]_net_1\, \line4[14]_net_1\, 
        \line4[13]_net_1\, \line4[12]_net_1\, \line4[11]_net_1\, 
        \line4[10]_net_1\, \line4[9]_net_1\, \line4[8]_net_1\, 
        \line4[7]_net_1\, \line4[6]_net_1\, \line4[5]_net_1\, 
        \line4[4]_net_1\, \line4[3]_net_1\, \line4[2]_net_1\, 
        \line4[1]_net_1\, \line4[0]_net_1\, line4_0_62, 
        \line3[63]_net_1\, \line3_or[32]_net_1\, 
        \line3[62]_net_1\, \line3[61]_net_1\, \line3[60]_net_1\, 
        \line3[59]_net_1\, \line3[58]_net_1\, \line3[57]_net_1\, 
        \line3[56]_net_1\, \line3[55]_net_1\, \line3[54]_net_1\, 
        \line3[53]_net_1\, \line3[52]_net_1\, \line3[51]_net_1\, 
        \line3[50]_net_1\, \line3[49]_net_1\, \line3[48]_net_1\, 
        \line3[47]_net_1\, \line3[46]_net_1\, \line3[45]_net_1\, 
        \line3[44]_net_1\, \line3[43]_net_1\, \line3[42]_net_1\, 
        \line3[41]_net_1\, \line3[40]_net_1\, \line3[39]_net_1\, 
        \line3[38]_net_1\, \line3[37]_net_1\, \line3[36]_net_1\, 
        \line3[35]_net_1\, \line3[34]_net_1\, \line3[33]_net_1\, 
        \line3[32]_net_1\, line3_0, \line3[31]_net_1\, 
        \line3_or[0]_net_1\, \line3[30]_net_1\, \line3[29]_net_1\, 
        \line3[28]_net_1\, \line3[27]_net_1\, \line3[26]_net_1\, 
        \line3[25]_net_1\, \line3[24]_net_1\, \line3[23]_net_1\, 
        \line3[22]_net_1\, \line3[21]_net_1\, \line3[20]_net_1\, 
        \line3[19]_net_1\, \line3[18]_net_1\, \line3[17]_net_1\, 
        \line3[16]_net_1\, \line3[15]_net_1\, \line3[14]_net_1\, 
        \line3[13]_net_1\, \line3[12]_net_1\, \line3[11]_net_1\, 
        \line3[10]_net_1\, \line3[9]_net_1\, \line3[8]_net_1\, 
        \line3[7]_net_1\, \line3[6]_net_1\, \line3[5]_net_1\, 
        \line3[4]_net_1\, \line3[3]_net_1\, \line3[2]_net_1\, 
        \line3[1]_net_1\, \line3[0]_net_1\, line3_0_62, 
        \line2[63]_net_1\, \line2_or[32]_net_1\, 
        \line2[62]_net_1\, \line2[61]_net_1\, \line2[60]_net_1\, 
        \line2[59]_net_1\, \line2[58]_net_1\, \line2[57]_net_1\, 
        \line2[56]_net_1\, \line2[55]_net_1\, \line2[54]_net_1\, 
        \line2[53]_net_1\, \line2[52]_net_1\, \line2[51]_net_1\, 
        \line2[50]_net_1\, \line2[49]_net_1\, \line2[48]_net_1\, 
        \line2[47]_net_1\, \line2[46]_net_1\, \line2[45]_net_1\, 
        \line2[44]_net_1\, \line2[43]_net_1\, \line2[42]_net_1\, 
        \line2[41]_net_1\, \line2[40]_net_1\, \line2[39]_net_1\, 
        \line2[38]_net_1\, \line2[37]_net_1\, \line2[36]_net_1\, 
        \line2[35]_net_1\, \line2[34]_net_1\, \line2[33]_net_1\, 
        \line2[32]_net_1\, line2_0, \line2[31]_net_1\, 
        \line2_or[0]_net_1\, \line2[30]_net_1\, \line2[29]_net_1\, 
        \line2[28]_net_1\, \line2[27]_net_1\, \line2[26]_net_1\, 
        \line2[25]_net_1\, \line2[24]_net_1\, \line2[23]_net_1\, 
        \line2[22]_net_1\, \line2[21]_net_1\, \line2[20]_net_1\, 
        \line2[19]_net_1\, \line2[18]_net_1\, \line2[17]_net_1\, 
        \line2[16]_net_1\, \line2[15]_net_1\, \line2[14]_net_1\, 
        \line2[13]_net_1\, \line2[12]_net_1\, \line2[11]_net_1\, 
        \line2[10]_net_1\, \line2[9]_net_1\, \line2[8]_net_1\, 
        \line2[7]_net_1\, \line2[6]_net_1\, \line2[5]_net_1\, 
        \line2[4]_net_1\, \line2[3]_net_1\, \line2[2]_net_1\, 
        \line2[1]_net_1\, \line2[0]_net_1\, line2_0_62, 
        \line1[63]_net_1\, \line1_or[32]_net_1\, 
        \line1[62]_net_1\, \line1[61]_net_1\, \line1[60]_net_1\, 
        \line1[59]_net_1\, \line1[58]_net_1\, \line1[57]_net_1\, 
        \line1[56]_net_1\, \line1[55]_net_1\, \line1[54]_net_1\, 
        \line1[53]_net_1\, \line1[52]_net_1\, \line1[51]_net_1\, 
        \line1[50]_net_1\, \line1[49]_net_1\, \line1[48]_net_1\, 
        \line1[47]_net_1\, \line1[46]_net_1\, \line1[45]_net_1\, 
        \line1[44]_net_1\, \line1[43]_net_1\, \line1[42]_net_1\, 
        \line1[41]_net_1\, \line1[40]_net_1\, \line1[39]_net_1\, 
        \line1[38]_net_1\, \line1[37]_net_1\, \line1[36]_net_1\, 
        \line1[35]_net_1\, \line1[34]_net_1\, \line1[33]_net_1\, 
        \line1[32]_net_1\, line1_0, \line1[31]_net_1\, 
        \line1_or[0]_net_1\, \line1[30]_net_1\, \line1[29]_net_1\, 
        \line1[28]_net_1\, \line1[27]_net_1\, \line1[26]_net_1\, 
        \line1[25]_net_1\, \line1[24]_net_1\, \line1[23]_net_1\, 
        \line1[22]_net_1\, \line1[21]_net_1\, \line1[20]_net_1\, 
        \line1[19]_net_1\, \line1[18]_net_1\, \line1[17]_net_1\, 
        \line1[16]_net_1\, \line1[15]_net_1\, \line1[14]_net_1\, 
        \line1[13]_net_1\, \line1[12]_net_1\, \line1[11]_net_1\, 
        \line1[10]_net_1\, \line1[9]_net_1\, \line1[8]_net_1\, 
        \line1[7]_net_1\, \line1[6]_net_1\, \line1[5]_net_1\, 
        \line1[4]_net_1\, \line1[3]_net_1\, \line1[2]_net_1\, 
        \line1[1]_net_1\, \line1[0]_net_1\, line1_0_62, 
        \line0[63]_net_1\, \line0_or[32]_net_1\, 
        \line0[62]_net_1\, \line0[61]_net_1\, \line0[60]_net_1\, 
        \line0[59]_net_1\, \line0[58]_net_1\, \line0[57]_net_1\, 
        \line0[56]_net_1\, \line0[55]_net_1\, \line0[54]_net_1\, 
        \line0[53]_net_1\, \line0[52]_net_1\, \line0[51]_net_1\, 
        \line0[50]_net_1\, \line0[49]_net_1\, \line0[48]_net_1\, 
        \line0[47]_net_1\, \line0[46]_net_1\, \line0[45]_net_1\, 
        \line0[44]_net_1\, \line0[43]_net_1\, \line0[42]_net_1\, 
        \line0[41]_net_1\, \line0[40]_net_1\, \line0[39]_net_1\, 
        \line0[38]_net_1\, \line0[37]_net_1\, \line0[36]_net_1\, 
        \line0[35]_net_1\, \line0[34]_net_1\, \line0[33]_net_1\, 
        \line0[32]_net_1\, line0_0, \line0[31]_net_1\, 
        \line0_or[0]_net_1\, \line0[30]_net_1\, \line0[29]_net_1\, 
        \line0[28]_net_1\, \line0[27]_net_1\, \line0[26]_net_1\, 
        \line0[25]_net_1\, \line0[24]_net_1\, \line0[23]_net_1\, 
        \line0[22]_net_1\, \line0[21]_net_1\, \line0[20]_net_1\, 
        \line0[19]_net_1\, \line0[18]_net_1\, \line0[17]_net_1\, 
        \line0[16]_net_1\, \line0[15]_net_1\, \line0[14]_net_1\, 
        \line0[13]_net_1\, \line0[12]_net_1\, \line0[11]_net_1\, 
        \line0[10]_net_1\, \line0[9]_net_1\, \line0[8]_net_1\, 
        \line0[7]_net_1\, \line0[6]_net_1\, \line0[5]_net_1\, 
        \line0[4]_net_1\, \line0[3]_net_1\, \line0[2]_net_1\, 
        \line0[1]_net_1\, \line0[0]_net_1\, line0_0_62, 
        \raddr_pos[3]_net_1\, N_3_0, \raddr_pos[2]_net_1\, 
        \raddr_pos[1]_net_1\, \raddr_pos[0]_net_1\, 
        \raddr_pos_fast[0]_net_1\, \raddr_pos_0_rep1\, 
        \raddr_pos_0_rep2\, \raddr_pos_fast[1]_net_1\, 
        \raddr_pos_1_rep1\, \raddr_pos_1_rep2\, 
        \raddr_pos_fast_fast[0]_net_1\, \raddr_pos_fast_0_rep1\, 
        \raddr_pos_fast_0_rep2\, N_1623, \data_out_31_1_1[0]\, 
        N_1399, N_919, N_1143, N_1653, \data_out_31_1_1[30]\, 
        N_1429, N_949, N_1173, N_1626, \data_out_31_1_1[3]\, 
        N_1402, N_922, N_1146, N_1625, \data_out_31_1_1[2]\, 
        N_1401, N_921, N_1145, N_1624, \data_out_31_1_1[1]\, 
        N_1400, N_920, N_1144, N_1651, \data_out_31_1_1[28]\, 
        N_1427, N_947, N_1171, N_1649, \data_out_31_1_1[26]\, 
        N_1425, N_945, N_1169, N_1646, \data_out_31_1_1[23]\, 
        N_1422, N_942, N_1166, N_1637, \data_out_31_1_1[14]\, 
        N_1413, N_933, N_1157, N_1650, \data_out_31_1_1[27]\, 
        N_1426, N_946, N_1170, N_1648, \data_out_31_1_1[25]\, 
        N_1424, N_944, N_1168, N_1652, \data_out_31_1_1[29]\, 
        N_1428, N_948, N_1172, N_1636, \data_out_31_1_1[13]\, 
        N_1412, N_932, N_1156, N_1634, \data_out_31_1_1[11]\, 
        N_1410, N_930, N_1154, N_1633, \data_out_31_1_1[10]\, 
        N_1409, N_929, N_1153, N_1628, \data_out_31_1_1[5]\, 
        N_1404, N_924, N_1148, N_1627, \data_out_31_1_1[4]\, 
        N_1403, N_923, N_1147, N_1640, \data_out_31_1_1[17]\, 
        N_1416, N_936, N_1160, N_1630, \data_out_31_1_1[7]\, 
        N_1406, N_926, N_1150, N_1645, \data_out_31_1_1[22]\, 
        N_1421, N_941, N_1165, N_1644, \data_out_31_1_1[21]\, 
        N_1420, N_940, N_1164, N_1643, \data_out_31_1_1[20]\, 
        N_1419, N_939, N_1163, N_1654, \data_out_31_1_1[31]\, 
        N_1430, N_950, N_1174, N_1639, \data_out_31_1_1[16]\, 
        N_1415, N_935, N_1159, N_1632, \data_out_31_1_1[9]\, 
        N_1408, N_928, N_1152, N_1635, \data_out_31_1_1[12]\, 
        N_1411, N_931, N_1155, N_1641, \data_out_31_1_1[18]\, 
        N_1417, N_937, N_1161, N_1631, \data_out_31_1_1[8]\, 
        N_1407, N_927, N_1151, N_1629, \data_out_31_1_1[6]\, 
        N_1405, N_925, N_1149, N_1642, \data_out_31_1_1[19]\, 
        N_1418, N_938, N_1162, N_1638, \data_out_31_1_1[15]\, 
        N_1414, N_934, N_1158, N_1647, \data_out_31_1_1[24]\, 
        N_1423, N_943, N_1167, \data_out_7_1_1[7]\, 
        \data_out_29_1_1[4]\, \data_out_29_1_1[3]\, 
        \data_out_29_1_1[11]\, \data_out_22_1_1[7]\, 
        \data_out_29_1_1[10]\, \data_out_29_1_1[8]\, 
        \data_out_29_1_1[5]\, \data_out_29_1_1[0]\, 
        \data_out_29_1_1[23]\, \data_out_29_1_1[9]\, 
        \data_out_29_1_1[6]\, \data_out_29_1_1[7]\, 
        \data_out_29_1_1[17]\, \data_out_29_1_1[12]\, 
        \data_out_29_1_1[14]\, \data_out_29_1_1[13]\, 
        \data_out_29_1_1[1]\, \data_out_7_1_1[29]\, 
        \data_out_22_1_1[9]\, \data_out_22_1_1[4]\, 
        \data_out_29_1_1[26]\, \data_out_14_1_1[7]\, 
        \data_out_29_1_1[22]\, \data_out_29_1_1[21]\, 
        \data_out_29_1_1[16]\, \data_out_22_1_1[12]\, 
        \data_out_22_1_1[11]\, \data_out_22_1_1[5]\, 
        \data_out_22_1_1[1]\, \data_out_29_1_1[25]\, 
        \data_out_29_1_1[18]\, \data_out_14_1_1[23]\, 
        \data_out_29_1_1[15]\, \data_out_22_1_1[23]\, 
        \data_out_29_1_1[2]\, \data_out_7_1_1[31]\, 
        \data_out_7_1_1[30]\, \data_out_22_1_1[10]\, 
        \data_out_14_1_1[14]\, \data_out_14_1_1[10]\, 
        \data_out_22_1_1[2]\, \data_out_29_1_1[24]\, 
        \data_out_7_1_1[23]\, \data_out_14_1_1[17]\, 
        \data_out_14_1_1[15]\, \data_out_14_1_1[13]\, 
        \data_out_7_1_1[26]\, \data_out_14_1_1[9]\, 
        \data_out_14_1_1[5]\, \data_out_14_1_1[3]\, 
        \data_out_29_1_1[20]\, \data_out_29_1_1[19]\, 
        \data_out_22_1_1[25]\, \data_out_14_1_1[20]\, 
        \data_out_22_1_1[13]\, \data_out_7_1_1[28]\, 
        \data_out_7_1_1[27]\, \data_out_7_1_1[24]\, 
        \data_out_14_1_1[8]\, \data_out_7_1_1[21]\, 
        \data_out_7_1_1[20]\, \data_out_14_1_1[4]\, 
        \data_out_29_1_1[28]\, \data_out_29_1_1[27]\, 
        \data_out_14_1_1[0]\, \data_out_7_1_1[14]\, 
        \data_out_7_1_1[13]\, \data_out_7_1_1[12]\, 
        \data_out_7_1_1[9]\, \data_out_22_1_1[31]\, 
        \data_out_22_1_1[26]\, \data_out_14_1_1[30]\, 
        \data_out_22_1_1[24]\, \data_out_14_1_1[21]\, 
        \data_out_22_1_1[15]\, \data_out_22_1_1[14]\, 
        \data_out_14_1_1[18]\, \data_out_7_1_1[19]\, 
        \data_out_29_1_1[30]\, \data_out_7_1_1[17]\, 
        \data_out_7_1_1[16]\, \data_out_7_1_1[15]\, 
        \data_out_14_1_1[1]\, \data_out_7_1_1[11]\, 
        \data_out_7_1_1[10]\, \data_out_22_1_1[30]\, 
        \data_out_22_1_1[29]\, \data_out_14_1_1[29]\, 
        \data_out_22_1_1[19]\, \data_out_7_1_1[22]\, 
        \data_out_22_1_1[17]\, \data_out_14_1_1[19]\, 
        \data_out_22_1_1[16]\, \data_out_14_1_1[16]\, 
        \data_out_22_1_1[8]\, \data_out_14_1_1[25]\, 
        \data_out_29_1_1[29]\, \data_out_14_1_1[2]\, 
        \data_out_7_1_1[25]\, \data_out_22_1_1[18]\, 
        \data_out_22_1_1[21]\, \data_out_22_1_1[20]\, 
        \data_out_14_1_1[26]\, \data_out_7_1_1[18]\, 
        \data_out_22_1_1[6]\, \data_out_14_1_1[24]\, 
        \data_out_7_1_1[4]\, \data_out_7_1_1[6]\, 
        \data_out_22_1_1[28]\, \data_out_14_1_1[11]\, 
        \data_out_22_1_1[0]\, \data_out_7_1_1[8]\, 
        \data_out_29_1_1[31]\, \data_out_22_1_1[27]\, 
        \data_out_7_1_1[3]\, \data_out_22_1_1[3]\, 
        \data_out_14_1_1[12]\, \data_out_7_1_1[5]\, 
        \data_out_7_1_1[1]\, \data_out_22_1_1[22]\, 
        \data_out_14_1_1[6]\, \data_out_14_1_1[22]\, 
        \data_out_14_1_1[27]\, \data_out_14_1_1[31]\, 
        \data_out_7_1_1[0]\, \data_out_7_1_1[2]\, 
        \data_out_14_1_1[28]\, N_49, N_49_mux, N_13_0, N_39, N_30, 
        N_23_0, N_15_0 : std_logic;

begin 

    data_out_ready <= data_out_ready_net_1;
    SHA256_Module_0_data_available <= 
        \SHA256_Module_0_data_available\;

    \raddr_pos_RNI0KE04[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_947, D => N_1171, Y => 
        \data_out_31_1_1[28]\);
    
    m43 : CFG4
      generic map(INIT => x"1054")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_39, D => CertificationSystem_sb_0_GPIO_9_M2F, Y => 
        line6_0_62);
    
    \line3[15]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[15]_net_1\);
    
    \line5[19]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[19]_net_1\);
    
    \line3[41]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[41]_net_1\);
    
    \line1[30]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[30]_net_1\);
    
    \line1[16]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[16]_net_1\);
    
    \line6[17]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[17]_net_1\);
    
    \line1[22]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[22]_net_1\);
    
    \line0_RNIJAC11[20]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[20]_net_1\, B => \line0[20]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[20]\);
    
    \line2_RNI793I[19]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[19]_net_1\, B => \line2[19]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[19]\);
    
    \line7[61]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[61]_net_1\);
    
    \line5[33]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[33]_net_1\);
    
    \line3[0]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[0]_net_1\);
    
    \line6[45]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[45]_net_1\);
    
    \line1[14]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[14]_net_1\);
    
    \raddr_pos_fast[1]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_fast[1]_net_1\);
    
    \line6_RNIUUED1[55]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[23]\, C => \line7[55]_net_1\, D => 
        \line6[55]_net_1\, Y => N_1646);
    
    \raddr_pos_RNI2R7D7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1646, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[23]\, D => N_1422, Y => N_1710);
    
    \line7[27]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[27]_net_1\);
    
    \line4_RNI9JQE2[59]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[27]\, C => \line5[59]_net_1\, D => 
        \line4[59]_net_1\, Y => N_1426);
    
    \line1[11]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[11]_net_1\);
    
    \line7[47]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[47]_net_1\);
    
    \line6_RNISQCD1[50]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[18]\, C => \line7[50]_net_1\, D => 
        \line6[50]_net_1\, Y => N_1641);
    
    \line2_RNIJ6151[9]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[9]_net_1\, B => \line2[9]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[9]\);
    
    \raddr_pos_RNIHVHC4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_920, D => N_1144, Y => 
        \data_out_31_1_1[1]\);
    
    \line2_RNI7J3U[55]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[23]\, C => \line3[55]_net_1\, D => 
        \line2[55]_net_1\, Y => N_1166);
    
    \line2[50]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[50]_net_1\);
    
    \raddr_pos_RNIBD6B3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_933, D => N_1157, Y => 
        \data_out_31_1_1[14]\);
    
    \line0_RNI6QE81[21]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[21]_net_1\, B => \line0[21]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[21]\);
    
    \raddr_pos_RNIE53C7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1626, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[3]\, D => N_1402, Y => N_1690);
    
    \line0[32]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[32]_net_1\);
    
    m40 : CFG4
      generic map(INIT => x"4051")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_39, D => CertificationSystem_sb_0_GPIO_9_M2F, Y => 
        line7_0_62);
    
    m14 : CFG4
      generic map(INIT => x"40FB")

      port map(A => waddr_in_net_0(2), B => waddr_in_net_0(3), C
         => N_13_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => N_15_0);
    
    \line8[21]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line8_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        reg_17x32_0_valid_bytes_0(1));
    
    \line6[20]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[20]_net_1\);
    
    \line1[56]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[56]_net_1\);
    
    \line3[36]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[36]_net_1\);
    
    \line3[4]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[4]_net_1\);
    
    \line0[20]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[20]_net_1\);
    
    \line6[55]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[55]_net_1\);
    
    \line2_RNIRADA1[58]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[26]\, C => \line3[58]_net_1\, D => 
        \line2[58]_net_1\, Y => N_1169);
    
    \line6_RNIG22K[9]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[9]_net_1\, B => \line6[9]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[9]\);
    
    \line0[56]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[56]_net_1\);
    
    \line0_RNIV9O01[10]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[10]_net_1\, B => \line0[10]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[10]\);
    
    \line0_RNIFG4A1[7]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[7]_net_1\, B => \line0[7]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[7]\);
    
    \line2[49]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[49]_net_1\);
    
    \line2[20]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[20]_net_1\);
    
    \line7[12]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[12]_net_1\);
    
    \line6_RNIHAN61[43]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[11]\, C => \line7[43]_net_1\, D => 
        \line6[43]_net_1\, Y => N_1634);
    
    \line5[22]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[22]_net_1\);
    
    \line4_RNIKC4F1[36]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[4]\, C => \line5[36]_net_1\, D => 
        \line4[36]_net_1\, Y => N_1403);
    
    \line3[61]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[61]_net_1\);
    
    \line3[29]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[29]_net_1\);
    
    \line1[54]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[54]_net_1\);
    
    \line5[38]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[38]_net_1\);
    
    \line3[34]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[34]_net_1\);
    
    \line3[7]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[7]_net_1\);
    
    \line4[61]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[61]_net_1\);
    
    \line0[54]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[54]_net_1\);
    
    \line0[8]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[8]_net_1\);
    
    \line0[49]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[49]_net_1\);
    
    \line7[52]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[52]_net_1\);
    
    \raddr_pos_RNIJ0AG4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_924, D => N_1148, Y => 
        \data_out_31_1_1[5]\);
    
    \line1[51]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[51]_net_1\);
    
    \line4[50]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[50]_net_1\);
    
    \line3[31]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[31]_net_1\);
    
    \line0[51]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[51]_net_1\);
    
    \line5[42]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[42]_net_1\);
    
    \line2[16]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[16]_net_1\);
    
    \raddr_pos_RNIEOBU6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1634, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[11]\, D => N_1410, Y => N_1698);
    
    \raddr_pos_RNI6AJB8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1647, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[24]\, D => N_1423, Y => N_1711);
    
    \ren_pos\ : SLE
      port map(D => data_out_ready_0_sqmuxa, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => ren_pos);
    
    \line0_RNIB2652[35]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[3]\, 
        C => \line1[35]_net_1\, D => \line0[35]_net_1\, Y => 
        N_922);
    
    \line6[60]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[60]_net_1\);
    
    m16 : CFG4
      generic map(INIT => x"4051")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_15_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => line5_0_62);
    
    \line1[23]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[23]_net_1\);
    
    \line6_RNI52AP[12]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[12]_net_1\, B => \line6[12]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[12]\);
    
    \line4[8]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[8]_net_1\);
    
    \line3[55]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[55]_net_1\);
    
    \line7[30]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[30]_net_1\);
    
    \line0_RNIR60V1[41]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_7_1_1[9]\, C => \line1[41]_net_1\, D => 
        \line0[41]_net_1\, Y => N_928);
    
    \line6[2]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[2]_net_1\);
    
    \line4[0]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[0]_net_1\);
    
    \line4[42]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[42]_net_1\);
    
    \line2[14]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[14]_net_1\);
    
    \line0_RNIE6752[61]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[29]\, C => \line1[61]_net_1\, D => 
        \line0[61]_net_1\, Y => N_948);
    
    \line7[4]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[4]_net_1\);
    
    \line0_RNI6ASR1[44]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[12]\, 
        C => \line1[44]_net_1\, D => \line0[44]_net_1\, Y => 
        N_931);
    
    \raddr_pos_RNI6LBR7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1644, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[21]\, D => N_1420, Y => N_1708);
    
    \line0_RNI26SR1[43]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[11]\, 
        C => \line1[43]_net_1\, D => \line0[43]_net_1\, Y => 
        N_930);
    
    \line1[49]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[49]_net_1\);
    
    \line2[11]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[11]_net_1\);
    
    raddr_pos_fast_0_rep1 : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_fast_0_rep1\);
    
    \line3[2]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[2]_net_1\);
    
    \line0_RNIN20V1[40]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_7_1_1[8]\, C => \line1[40]_net_1\, D => 
        \line0[40]_net_1\, Y => N_927);
    
    \line4[32]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[32]_net_1\);
    
    \line4[16]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[16]_net_1\);
    
    \line2[32]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[32]_net_1\);
    
    \line6_RNIHEAP[18]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[18]_net_1\, B => \line6[18]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[18]\);
    
    \line4[7]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[7]_net_1\);
    
    \line6_RNIOO8S[29]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[29]_net_1\, B => \line6[29]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[29]\);
    
    \line5[17]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[17]_net_1\);
    
    \line3[9]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[9]_net_1\);
    
    \line0[33]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[33]_net_1\);
    
    \line4_RNI9A652[43]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[11]\, C => \line5[43]_net_1\, D => 
        \line4[43]_net_1\, Y => N_1410);
    
    \line4[1]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[1]_net_1\);
    
    \line1[35]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[35]_net_1\);
    
    \line3[49]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[49]_net_1\);
    
    \line2_RNIDI4K[28]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line2[28]_net_1\, B => \line3[28]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_14_1_1[28]\);
    
    \line0[12]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[12]_net_1\);
    
    \line2_RNI4UKC1[0]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[0]_net_1\, B => \line2[0]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[0]\);
    
    \line0_RNIVIIS1[55]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[23]\, 
        C => \line1[55]_net_1\, D => \line0[55]_net_1\, Y => 
        N_942);
    
    \raddr_pos_RNI8BKB8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1649, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[26]\, D => N_1425, Y => N_1713);
    
    \line4[14]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[14]_net_1\);
    
    \line2_RNICC7P[22]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[22]_net_1\, B => \line2[22]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[22]\);
    
    \line7[13]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[13]_net_1\);
    
    \line4_RNIOQ652[47]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[15]\, C => \line5[47]_net_1\, D => 
        \line4[47]_net_1\, Y => N_1414);
    
    \line1[28]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[28]_net_1\);
    
    \line5[23]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[23]_net_1\);
    
    m2 : CFG2
      generic map(INIT => x"B")

      port map(A => CertificationSystem_sb_0_GPIO_1_M2F, B => 
        CertificationSystem_sb_0_GPIO_9_M2F, Y => N_3_0);
    
    \line2[4]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[4]_net_1\);
    
    \line6_RNI54CP[21]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[21]_net_1\, B => \line6[21]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[21]\);
    
    \line6[1]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[1]_net_1\);
    
    \line0_RNI2PA11[19]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[19]_net_1\, B => \line0[19]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[19]\);
    
    \line4[11]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[11]_net_1\);
    
    \line6[30]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[30]_net_1\);
    
    \raddr_pos_RNIGLAB3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_938, D => N_1162, Y => 
        \data_out_31_1_1[19]\);
    
    \line6_RNIPUEG1[62]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[30]\, C => \line7[62]_net_1\, D => 
        \line6[62]_net_1\, Y => N_1653);
    
    \line7[53]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[53]_net_1\);
    
    \line6_RNI7BDG1[61]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[29]\, C => \line7[61]_net_1\, D => 
        \line6[61]_net_1\, Y => N_1652);
    
    \line0_RNIRI652[39]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[7]\, 
        C => \line1[39]_net_1\, D => \line0[39]_net_1\, Y => 
        N_926);
    
    \line2_RNI8QP61[62]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[30]\, C => \line3[62]_net_1\, D => 
        \line2[62]_net_1\, Y => N_1173);
    
    \line7[7]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[7]_net_1\);
    
    \line1[19]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[19]_net_1\);
    
    \line1[0]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[0]_net_1\);
    
    \line0_RNIUKA11[17]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[17]_net_1\, B => \line0[17]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[17]\);
    
    \line5[43]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[43]_net_1\);
    
    \line4[20]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[20]_net_1\);
    
    \line2[55]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[55]_net_1\);
    
    \line0_RNIVEES1[46]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[14]\, 
        C => \line1[46]_net_1\, D => \line0[46]_net_1\, Y => 
        N_933);
    
    \line6_RNI8L941[39]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[7]\, C => \line7[39]_net_1\, D => 
        \line6[39]_net_1\, Y => N_1630);
    
    \line5[50]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[50]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \raddr_pos_RNI7GRP3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_950, D => N_1174, Y => 
        \data_out_31_1_1[31]\);
    
    \line6[25]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[25]_net_1\);
    
    \line3[1]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[1]_net_1\);
    
    \line0[38]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[38]_net_1\);
    
    \line2[47]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[47]_net_1\);
    
    \line8[29]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line8_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        reg_17x32_0_last_word(1));
    
    \line7_or[32]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line7_0, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line7_or[32]_net_1\);
    
    \line4_RNI9QH81[16]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[16]_net_1\, B => \line4[16]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[16]\);
    
    \line0[25]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[25]_net_1\);
    
    \line2_RNIL0A51[63]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[31]\, C => \line3[63]_net_1\, D => 
        \line2[63]_net_1\, Y => N_1174);
    
    \line0_RNINE652[38]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[6]\, 
        C => \line1[38]_net_1\, D => \line0[38]_net_1\, Y => 
        N_925);
    
    \line3[27]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[27]_net_1\);
    
    \line4_RNIHI652[45]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[13]\, C => \line5[45]_net_1\, D => 
        \line4[45]_net_1\, Y => N_1412);
    
    \line0_RNI784A1[3]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[3]_net_1\, B => \line0[3]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[3]\);
    
    \line2[25]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[25]_net_1\);
    
    \line4[43]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[43]_net_1\);
    
    \line7[18]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[18]_net_1\);
    
    \line3[12]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[12]_net_1\);
    
    \line5[28]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[28]_net_1\);
    
    \line0[47]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[47]_net_1\);
    
    \line2_RNI8ERN[26]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[26]_net_1\, B => \line2[26]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep2\, Y => 
        \data_out_14_1_1[26]\);
    
    \line5[36]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[36]_net_1\);
    
    \line4[33]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[33]_net_1\);
    
    \line2[33]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[33]_net_1\);
    
    \raddr_pos_RNIVVIP3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_940, D => N_1164, Y => 
        \data_out_31_1_1[21]\);
    
    \line7[58]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[58]_net_1\);
    
    \line6_RNIMMED1[53]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[21]\, C => \line7[53]_net_1\, D => 
        \line6[53]_net_1\, Y => N_1644);
    
    \line4[55]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[55]_net_1\);
    
    \line1[59]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[59]_net_1\);
    
    \line3[39]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[39]_net_1\);
    
    \raddr_pos_RNI04IV6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1639, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[16]\, D => N_1415, Y => N_1703);
    
    \line0[59]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[59]_net_1\);
    
    \line4_RNIRCTI[9]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line5[9]_net_1\, B => \line4[9]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_22_1_1[9]\);
    
    \line5[48]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[48]_net_1\);
    
    \line0[13]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[13]_net_1\);
    
    \line6[42]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[42]_net_1\);
    
    \line6_RNIKK8S[27]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[27]_net_1\, B => \line6[27]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[27]\);
    
    \line5[34]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[34]_net_1\);
    
    \line4_RNISDH81[10]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[10]_net_1\, B => \line4[10]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[10]\);
    
    \line1[9]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[9]_net_1\);
    
    \line1_or[32]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line1_0, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line1_or[32]_net_1\);
    
    \raddr_pos_RNIHS2A3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_934, D => N_1158, Y => 
        \data_out_31_1_1[15]\);
    
    \line4_RNIBSH81[17]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[17]_net_1\, B => \line4[17]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[17]\);
    
    \line3[5]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[5]_net_1\);
    
    \raddr_pos_RNIMLSR7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1654, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[31]\, D => N_1430, Y => N_1718);
    
    \line3[8]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[8]_net_1\);
    
    \line6_RNIO4941[35]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[3]\, C => \line7[35]_net_1\, D => 
        \line6[35]_net_1\, Y => N_1626);
    
    \line2_RNI7FVT[46]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[14]\, C => \line3[46]_net_1\, D => 
        \line2[46]_net_1\, Y => N_1157);
    
    \line7[35]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[35]_net_1\);
    
    \line5[31]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[31]_net_1\);
    
    \line4_RNI1KJ81[21]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[21]_net_1\, B => \line4[21]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[21]\);
    
    \line1[47]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[47]_net_1\);
    
    \line6[10]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[10]_net_1\);
    
    \line1[7]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[7]_net_1\);
    
    \line1[60]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[60]_net_1\);
    
    \raddr_pos_RNIC4B87[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1624, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[1]\, D => N_1400, Y => N_1688);
    
    \line4[48]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[48]_net_1\);
    
    \line0[62]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[62]_net_1\);
    
    \line0_RNIDE4A1[6]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[6]_net_1\, B => \line0[6]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[6]\);
    
    \line2[6]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[6]_net_1\);
    
    \line6[52]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[52]_net_1\);
    
    \line2[19]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[19]_net_1\);
    
    \line6_RNI74AP[13]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[13]_net_1\, B => \line6[13]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[13]\);
    
    \line2_RNI5F1U[50]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[18]\, C => \line3[50]_net_1\, D => 
        \line2[50]_net_1\, Y => N_1161);
    
    \line2_RNIQS2I[13]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[13]_net_1\, B => \line2[13]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[13]\);
    
    \line4[38]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[38]_net_1\);
    
    \line3[47]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[47]_net_1\);
    
    \line2[38]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[38]_net_1\);
    
    \line7[20]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[20]_net_1\);
    
    \line6_RNIBQAG[5]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[5]_net_1\, B => \line7[5]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[5]\);
    
    \line6_RNIFUAG[7]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[7]_net_1\, B => \line7[7]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[7]\);
    
    \line7[40]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[40]_net_1\);
    
    \line0_RNI82371[28]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[28]_net_1\, B => \line0[28]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep2\, Y => 
        \data_out_7_1_1[28]\);
    
    \line0[18]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[18]_net_1\);
    
    \line2_RNI335K1[41]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_14_1_1[9]\, C => \line3[41]_net_1\, D => 
        \line2[41]_net_1\, Y => N_1152);
    
    \line2[3]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[3]_net_1\);
    
    \line0_RNI2S271[25]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[25]_net_1\, B => \line0[25]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep2\, Y => 
        \data_out_7_1_1[25]\);
    
    \line3[13]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[13]_net_1\);
    
    \line7[0]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[0]_net_1\);
    
    \line1[26]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[26]_net_1\);
    
    \line4_RNIK8GB1[29]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[29]_net_1\, B => \line4[29]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[29]\);
    
    \line4[19]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[19]_net_1\);
    
    \line2_RNINQ4I[20]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[20]_net_1\, B => \line2[20]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[20]\);
    
    \line7[1]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[1]_net_1\);
    
    \line6[35]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[35]_net_1\);
    
    \line1[17]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[17]_net_1\);
    
    \line5[9]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[9]_net_1\);
    
    \raddr_pos_RNID3RS3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_949, D => N_1173, Y => 
        \data_out_31_1_1[30]\);
    
    \raddr_pos_RNI3G9G4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_922, D => N_1146, Y => 
        \data_out_31_1_1[3]\);
    
    \line4[25]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[25]_net_1\);
    
    \line3[52]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[52]_net_1\);
    
    \line5[62]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[62]_net_1\);
    
    \line1[24]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[24]_net_1\);
    
    \line5[55]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[55]_net_1\);
    
    \line6[43]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[43]_net_1\);
    
    \raddr_pos_RNIU8CU6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1635, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[12]\, D => N_1411, Y => N_1699);
    
    m27 : CFG4
      generic map(INIT => x"1054")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_23_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => line2_0_62);
    
    \line6[5]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[5]_net_1\);
    
    \line0_RNI60371[27]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[27]_net_1\, B => \line0[27]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep2\, Y => 
        \data_out_7_1_1[27]\);
    
    \raddr_pos_RNIE75C7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1630, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[7]\, D => N_1406, Y => N_1694);
    
    \line1[21]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[21]_net_1\);
    
    \line0[36]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[36]_net_1\);
    
    \line4_RNIHUTE2[62]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[30]\, C => \line5[62]_net_1\, D => 
        \line4[62]_net_1\, Y => N_1429);
    
    \line0_RNIU5A32[32]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[0]\, 
        C => \line1[32]_net_1\, D => \line0[32]_net_1\, Y => 
        N_919);
    
    \line4_RNIMUTB2[55]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[23]\, C => \line5[55]_net_1\, D => 
        \line4[55]_net_1\, Y => N_1422);
    
    \line0_RNIDSK32[54]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[22]\, 
        C => \line1[54]_net_1\, D => \line0[54]_net_1\, Y => 
        N_941);
    
    \line7[5]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[5]_net_1\);
    
    \line1[2]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[2]_net_1\);
    
    \line6_RNI1GAG[0]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[0]_net_1\, B => \line7[0]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[0]\);
    
    \raddr_pos_RNIBO9G4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_923, D => N_1147, Y => 
        \data_out_31_1_1[4]\);
    
    \line0_RNI9A4A1[4]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[4]_net_1\, B => \line0[4]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[4]\);
    
    \line0[63]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[63]_net_1\);
    
    \raddr_pos_RNI9NHC4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_919, D => N_1143, Y => 
        \data_out_31_1_1[0]\);
    
    \line6_RNIDAAP[16]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[16]_net_1\, B => \line6[16]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[16]\);
    
    \line3[18]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[18]_net_1\);
    
    \line7[16]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[16]_net_1\);
    
    \line5[26]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[26]_net_1\);
    
    \line1[32]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[32]_net_1\);
    
    \line1[57]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[57]_net_1\);
    
    \line6[53]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[53]_net_1\);
    
    \line0[34]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[34]_net_1\);
    
    \line3[37]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[37]_net_1\);
    
    \line6_RNI0D941[37]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[5]\, C => \line7[37]_net_1\, D => 
        \line6[37]_net_1\, Y => N_1628);
    
    \line0[57]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[57]_net_1\);
    
    \line4_RNI5OJ81[23]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[23]_net_1\, B => \line4[23]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[23]\);
    
    \line8_or[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line8_0_62, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line8_or[0]_net_1\);
    
    \line6_RNI9BBG1[57]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[25]\, C => \line7[57]_net_1\, D => 
        \line6[57]_net_1\, Y => N_1648);
    
    \line0[31]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[31]_net_1\);
    
    \line7[56]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[56]_net_1\);
    
    \line6_or[32]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line6_0, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line6_or[32]_net_1\);
    
    \line2_RNIBG4K[27]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line2[27]_net_1\, B => \line3[27]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_14_1_1[27]\);
    
    \line0_RNI4M881[2]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[2]_net_1\, B => \line0[2]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[2]\);
    
    \line7[14]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[14]_net_1\);
    
    \line5[24]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[24]_net_1\);
    
    \line8[1]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line8_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        SHA256_Module_0_data_available_lastbank_8);
    
    \line6[48]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[48]_net_1\);
    
    \line5[10]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[10]_net_1\);
    
    \line5[46]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[46]_net_1\);
    
    \line2_RNIH4151[8]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[8]_net_1\, B => \line2[8]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[8]\);
    
    \line2[7]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[7]_net_1\);
    
    \raddr_pos_RNIE64C7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1628, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[5]\, D => N_1404, Y => N_1692);
    
    \line2_RNI0FM61[59]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[27]\, C => \line3[59]_net_1\, D => 
        \line2[59]_net_1\, Y => N_1170);
    
    \line7[11]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[11]_net_1\);
    
    m32 : CFG4
      generic map(INIT => x"80A2")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_30, D => CertificationSystem_sb_0_GPIO_9_M2F, Y => 
        line1_0);
    
    \line0_RNI92U82[60]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[28]\, C => \line1[60]_net_1\, D => 
        \line0[60]_net_1\, Y => N_947);
    
    \line5[21]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[21]_net_1\);
    
    \line4[6]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[6]_net_1\);
    
    \line7[54]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[54]_net_1\);
    
    \line0_RNIJAS82[58]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[26]\, C => \line1[58]_net_1\, D => 
        \line0[58]_net_1\, Y => N_945);
    
    \line5[39]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[39]_net_1\);
    
    \line4_RNI46652[42]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[10]\, C => \line5[42]_net_1\, D => 
        \line4[42]_net_1\, Y => N_1409);
    
    \line2[52]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[52]_net_1\);
    
    \line2_RNICE9P[31]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[31]_net_1\, B => \line2[31]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[31]\);
    
    \line6[15]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[15]_net_1\);
    
    \line2[17]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[17]_net_1\);
    
    \line5[44]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[44]_net_1\);
    
    \line4_RNIF0I81[19]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[19]_net_1\, B => \line4[19]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[19]\);
    
    \line7[51]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[51]_net_1\);
    
    \line6[22]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[22]_net_1\);
    
    \line0_RNI4U271[26]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[26]_net_1\, B => \line0[26]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep2\, Y => 
        \data_out_7_1_1[26]\);
    
    \line4[46]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[46]_net_1\);
    
    \line4_RNIVHJ81[20]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[20]_net_1\, B => \line4[20]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[20]\);
    
    \line0[22]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[22]_net_1\);
    
    \line2_RNIFQAQ1[34]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[2]\, 
        C => \line3[34]_net_1\, D => \line2[34]_net_1\, Y => 
        N_1145);
    
    \line6[58]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[58]_net_1\);
    
    \line3[53]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[53]_net_1\);
    
    \line5[63]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[63]_net_1\);
    
    \line5[41]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[41]_net_1\);
    
    \raddr_pos_RNIS7BU6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1633, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[10]\, D => N_1409, Y => N_1697);
    
    \line6_RNI57BG1[56]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[24]\, C => \line7[56]_net_1\, D => 
        \line6[56]_net_1\, Y => N_1647);
    
    \line2[22]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[22]_net_1\);
    
    \line7[25]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[25]_net_1\);
    
    \line4_RNITUHF1[40]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_22_1_1[8]\, 
        C => \line5[40]_net_1\, D => \line4[40]_net_1\, Y => 
        N_1407);
    
    \line4[36]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[36]_net_1\);
    
    \line2[36]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[36]_net_1\);
    
    \line4_RNI5FQE2[58]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[26]\, C => \line5[58]_net_1\, D => 
        \line4[58]_net_1\, Y => N_1425);
    
    \line4_RNISK4F1[38]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[6]\, C => \line5[38]_net_1\, D => 
        \line4[38]_net_1\, Y => N_1405);
    
    \line2[2]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[2]_net_1\);
    
    \line4[9]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[9]_net_1\);
    
    \line7[45]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[45]_net_1\);
    
    \line4[44]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[44]_net_1\);
    
    \line0[16]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[16]_net_1\);
    
    \line4[17]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[17]_net_1\);
    
    \line4[41]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[41]_net_1\);
    
    \line2[40]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[40]_net_1\);
    
    \line6_RNIMM8S[28]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[28]_net_1\, B => \line6[28]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[28]\);
    
    \line4[52]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[52]_net_1\);
    
    \raddr_pos_RNIBLEB3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_942, D => N_1166, Y => 
        \data_out_31_1_1[23]\);
    
    \line4[34]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[34]_net_1\);
    
    \line0[0]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[0]_net_1\);
    
    \line2[34]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[34]_net_1\);
    
    \line4_RNIOG4F1[37]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[5]\, C => \line5[37]_net_1\, D => 
        \line4[37]_net_1\, Y => N_1404);
    
    \line6[6]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[6]_net_1\);
    
    \line1[33]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[33]_net_1\);
    
    \line3[20]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[20]_net_1\);
    
    \line2_RNIQMDT[47]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[15]\, C => \line3[47]_net_1\, D => 
        \line2[47]_net_1\, Y => N_1158);
    
    \line0_RNI2K881[1]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[1]_net_1\, B => \line0[1]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[1]\);
    
    \line4[31]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[31]_net_1\);
    
    \line2[31]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[31]_net_1\);
    
    \line6[62]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[62]_net_1\);
    
    \line0[14]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[14]_net_1\);
    
    \line6_RNIQQED1[54]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[22]\, C => \line7[54]_net_1\, D => 
        \line6[54]_net_1\, Y => N_1645);
    
    \line2_RNIFNVT[48]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[16]\, C => \line3[48]_net_1\, D => 
        \line2[48]_net_1\, Y => N_1159);
    
    \line0[40]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[40]_net_1\);
    
    \line0_RNI0Q852[62]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[30]\, C => \line1[62]_net_1\, D => 
        \line0[62]_net_1\, Y => N_949);
    
    \line6_RNIGG8S[25]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[25]_net_1\, B => \line6[25]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[25]\);
    
    \line7[32]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[32]_net_1\);
    
    \line3[58]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[58]_net_1\);
    
    \line0_RNIDOK01[8]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[8]_net_1\, B => \line0[8]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[8]\);
    
    \line5_or[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line5_0_62, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line5_or[0]_net_1\);
    
    \line0[11]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[11]_net_1\);
    
    m22 : CFG4
      generic map(INIT => x"20FD")

      port map(A => waddr_in_net_0(2), B => waddr_in_net_0(3), C
         => N_13_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => N_23_0);
    
    m29 : CFG4
      generic map(INIT => x"10FE")

      port map(A => waddr_in_net_0(2), B => waddr_in_net_0(3), C
         => N_13_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => N_30);
    
    \line5[1]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[1]_net_1\);
    
    \line1[29]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[29]_net_1\);
    
    \line2[60]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[60]_net_1\);
    
    \line6[0]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[0]_net_1\);
    
    m34 : CFG4
      generic map(INIT => x"1054")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_30, D => CertificationSystem_sb_0_GPIO_9_M2F, Y => 
        line0_0_62);
    
    \line2[53]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[53]_net_1\);
    
    \line1[8]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[8]_net_1\);
    
    \line5[8]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[8]_net_1\);
    
    \line6_RNIFCAP[17]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[17]_net_1\, B => \line6[17]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[17]\);
    
    \line6[23]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[23]_net_1\);
    
    \line0[23]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[23]_net_1\);
    
    \line3[16]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[16]_net_1\);
    
    \line4_RNI0P4F1[39]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[7]\, C => \line5[39]_net_1\, D => 
        \line4[39]_net_1\, Y => N_1406);
    
    \line1[38]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[38]_net_1\);
    
    \raddr_pos_RNIDQDU6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1638, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[15]\, D => N_1414, Y => N_1702);
    
    \line1[40]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[40]_net_1\);
    
    \line4_RNIT6QE2[56]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[24]\, C => \line5[56]_net_1\, D => 
        \line4[56]_net_1\, Y => N_1423);
    
    \line4_RNIT3UB[0]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[0]_net_1\, B => \line5[0]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[0]\);
    
    \line4_RNIV5UB[1]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[1]_net_1\, B => \line5[1]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[1]\);
    
    \line2[23]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[23]_net_1\);
    
    raddr_pos_fast_0_rep2 : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_fast_0_rep2\);
    
    \line0_RNI9KO01[15]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[15]_net_1\, B => \line0[15]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[15]\);
    
    \line2_RNIHQGE1[6]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[6]_net_1\, B => \line2[6]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[6]\);
    
    \line0[39]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[39]_net_1\);
    
    \line6_RNIK0941[34]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[2]\, C => \line7[34]_net_1\, D => 
        \line6[34]_net_1\, Y => N_1625);
    
    \line3[14]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[14]_net_1\);
    
    \line5[15]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[15]_net_1\);
    
    \line6[32]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[32]_net_1\);
    
    \line4_RNI5MH81[14]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[14]_net_1\, B => \line4[14]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[14]\);
    
    \line3[40]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[40]_net_1\);
    
    \line5[37]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[37]_net_1\);
    
    \line6[46]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[46]_net_1\);
    
    \line2_RNIJSGE1[7]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[7]_net_1\, B => \line2[7]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[7]\);
    
    \line0_RNI8SE81[22]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[22]_net_1\, B => \line0[22]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[22]\);
    
    \line4[53]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[53]_net_1\);
    
    \line7[19]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[19]_net_1\);
    
    \line5[29]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[29]_net_1\);
    
    \line3[11]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[11]_net_1\);
    
    \line4[22]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[22]_net_1\);
    
    m36 : CFG2
      generic map(INIT => x"2")

      port map(A => N_49_mux, B => waddr_in_net_0(0), Y => 
        line8_0_62);
    
    \line7[60]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[60]_net_1\);
    
    \line5[52]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[52]_net_1\);
    
    \line2[58]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[58]_net_1\);
    
    \line0_RNIOGC11[23]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[23]_net_1\, B => \line0[23]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[23]\);
    
    \raddr_pos_RNIBS144[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_944, D => N_1168, Y => 
        \data_out_31_1_1[25]\);
    
    \line7[6]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[6]_net_1\);
    
    \line5[5]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[5]_net_1\);
    
    \line0_RNID0P32[63]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[31]\, 
        C => \line1[63]_net_1\, D => \line0[63]_net_1\, Y => 
        N_950);
    
    \line7[59]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[59]_net_1\);
    
    \line6[63]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[63]_net_1\);
    
    \line6[28]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[28]_net_1\);
    
    \line6[44]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[44]_net_1\);
    
    \line2[8]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[8]_net_1\);
    
    \line0[28]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[28]_net_1\);
    
    \raddr_pos_RNIT47A7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1625, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[2]\, D => N_1401, Y => N_1689);
    
    \raddr_pos_RNI3HAG4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_926, D => N_1150, Y => 
        \data_out_31_1_1[7]\);
    
    \line6_RNIII8S[26]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[26]_net_1\, B => \line6[26]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[26]\);
    
    \line4_RNIDUH81[18]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[18]_net_1\, B => \line4[18]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[18]\);
    
    \line0_RNIA2S82[56]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[24]\, C => \line1[56]_net_1\, D => 
        \line0[56]_net_1\, Y => N_943);
    
    \line7[33]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[33]_net_1\);
    
    \line5[49]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[49]_net_1\);
    
    \line6[56]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[56]_net_1\);
    
    \line1[10]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[10]_net_1\);
    
    m9_e : CFG4
      generic map(INIT => x"0002")

      port map(A => waddr_in_net_0(4), B => waddr_in_net_0(3), C
         => waddr_in_net_0(2), D => waddr_in_net_0(1), Y => N_49);
    
    \line6[41]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[41]_net_1\);
    
    \line0_RNIFQK01[9]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[9]_net_1\, B => \line0[9]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[9]\);
    
    \line4_RNIBIUB[7]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[7]_net_1\, B => \line5[7]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[7]\);
    
    \line2[28]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[28]_net_1\);
    
    m24 : CFG4
      generic map(INIT => x"4051")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_23_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => line3_0_62);
    
    \line4_RNI3MJ81[22]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[22]_net_1\, B => \line4[22]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[22]\);
    
    \line0[6]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[6]_net_1\);
    
    \line2_RNI6CRN[25]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[25]_net_1\, B => \line2[25]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep2\, Y => 
        \data_out_14_1_1[25]\);
    
    \line6_RNIIIED1[52]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[20]\, C => \line7[52]_net_1\, D => 
        \line6[52]_net_1\, Y => N_1643);
    
    \line8[20]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line8_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        reg_17x32_0_valid_bytes_0(0));
    
    \line6_RNI32CP[20]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[20]_net_1\, B => \line6[20]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[20]\);
    
    \line5[4]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[4]_net_1\);
    
    \line2[1]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[1]_net_1\);
    
    \line6[54]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[54]_net_1\);
    
    \line2_RNI473I[18]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[18]_net_1\, B => \line2[18]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[18]\);
    
    \line2[45]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[45]_net_1\);
    
    \line0_RNI1JGS1[51]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[19]\, 
        C => \line1[51]_net_1\, D => \line0[51]_net_1\, Y => 
        N_938);
    
    \line4_RNII6GB1[28]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[28]_net_1\, B => \line4[28]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[28]\);
    
    \line4[49]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[49]_net_1\);
    
    \line0[61]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[61]_net_1\);
    
    \line4[58]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[58]_net_1\);
    
    \line3[25]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[25]_net_1\);
    
    \line2_or[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line2_0_62, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line2_or[0]_net_1\);
    
    \line3[60]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[60]_net_1\);
    
    \line6[51]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[51]_net_1\);
    
    \line6_RNILEN61[44]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[12]\, C => \line7[44]_net_1\, D => 
        \line6[44]_net_1\, Y => N_1635);
    
    \line4[39]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[39]_net_1\);
    
    \line2[39]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[39]_net_1\);
    
    \line2_RNIS05I[23]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[23]_net_1\, B => \line2[23]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[23]\);
    
    \line6_RNI0VCD1[51]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[19]\, C => \line7[51]_net_1\, D => 
        \line6[51]_net_1\, Y => N_1642);
    
    \line4[60]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[60]_net_1\);
    
    \line0[45]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[45]_net_1\);
    
    \line2_RNILS551[54]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[22]\, C => \line3[54]_net_1\, D => 
        \line2[54]_net_1\, Y => N_1165);
    
    \line4_or[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line4_0_62, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line4_or[0]_net_1\);
    
    \line4_RNIR6SE2[60]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[28]\, C => \line5[60]_net_1\, D => 
        \line4[60]_net_1\, Y => N_1427);
    
    \line4_RNI18UB[2]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[2]_net_1\, B => \line5[2]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[2]\);
    
    \line1[50]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[50]_net_1\);
    
    \line3[30]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[30]_net_1\);
    
    \raddr_pos_RNI03HV6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1637, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[14]\, D => N_1413, Y => N_1701);
    
    \line1[27]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[27]_net_1\);
    
    \line7[38]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[38]_net_1\);
    
    \line0[50]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[50]_net_1\);
    
    \line0[19]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[19]_net_1\);
    
    \line6[33]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[33]_net_1\);
    
    \line6[12]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[12]_net_1\);
    
    \line3[56]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[56]_net_1\);
    
    \line1[62]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[62]_net_1\);
    
    \line0_RNIF6652[36]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[4]\, 
        C => \line1[36]_net_1\, D => \line0[36]_net_1\, Y => 
        N_923);
    
    \line2_RNI253I[17]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[17]_net_1\, B => \line2[17]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[17]\);
    
    \data_out_ready\ : SLE
      port map(D => \data_out_ready_1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => data_out_ready_net_1);
    
    \line4[4]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[4]_net_1\);
    
    \raddr_pos[3]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(3), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos[3]_net_1\);
    
    \line8[31]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line8_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        reg_17x32_0_last_word(3));
    
    \line6_RNI30AP[11]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[11]_net_1\, B => \line6[11]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[11]\);
    
    \line2_RNIDMGE1[4]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[4]_net_1\, B => \line2[4]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[4]\);
    
    m44 : CFG4
      generic map(INIT => x"20A8")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_39, D => CertificationSystem_sb_0_GPIO_9_M2F, Y => 
        line6_0);
    
    \line4[23]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[23]_net_1\);
    
    \line2_RNIEADT[44]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[12]\, C => \line3[44]_net_1\, D => 
        \line2[44]_net_1\, Y => N_1155);
    
    \line5[53]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[53]_net_1\);
    
    \line6[4]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[4]_net_1\);
    
    \line7[22]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[22]_net_1\);
    
    \line3[54]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[54]_net_1\);
    
    \line2_RNIJUAQ1[35]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[3]\, 
        C => \line3[35]_net_1\, D => \line2[35]_net_1\, Y => 
        N_1146);
    
    \line7[42]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[42]_net_1\);
    
    \line6_RNI37DG1[60]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[28]\, C => \line7[60]_net_1\, D => 
        \line6[60]_net_1\, Y => N_1651);
    
    \line4_RNIAITB2[52]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[20]\, C => \line5[52]_net_1\, D => 
        \line4[52]_net_1\, Y => N_1419);
    
    \line2_RNIHO551[53]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[21]\, C => \line3[53]_net_1\, D => 
        \line2[53]_net_1\, Y => N_1164);
    
    \line0[37]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[37]_net_1\);
    
    \line1[45]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[45]_net_1\);
    
    \line3[51]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[51]_net_1\);
    
    \line5[61]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[61]_net_1\);
    
    \line1[36]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[36]_net_1\);
    
    \raddr_pos_RNI1A488[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1651, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[28]\, D => N_1427, Y => N_1715);
    
    \line8[0]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line8_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => first_block);
    
    \line2[10]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[10]_net_1\);
    
    \line7_or[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line7_0_62, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line7_or[0]_net_1\);
    
    \raddr_pos_RNIUL3C7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1627, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[4]\, D => N_1403, Y => N_1691);
    
    \line0_RNI6EA32[34]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[2]\, 
        C => \line1[34]_net_1\, D => \line0[34]_net_1\, Y => 
        N_921);
    
    \line6_RNI9OAG[4]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[4]_net_1\, B => \line7[4]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[4]\);
    
    \line6_or[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line6_0_62, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line6_or[0]_net_1\);
    
    \line7[3]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[3]_net_1\);
    
    \line2_RNI3BVT[45]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[13]\, C => \line3[45]_net_1\, D => 
        \line2[45]_net_1\, Y => N_1156);
    
    \line6_RNI5RM41[40]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_29_1_1[8]\, 
        C => \line7[40]_net_1\, D => \line6[40]_net_1\, Y => 
        N_1631);
    
    \line7[17]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[17]_net_1\);
    
    \line5[27]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[27]_net_1\);
    
    \line3[45]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[45]_net_1\);
    
    \line6[38]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[38]_net_1\);
    
    \line4_RNI6OH81[15]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[15]_net_1\, B => \line4[15]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[15]\);
    
    \line6_RNI3IAG[1]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[1]_net_1\, B => \line7[1]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[1]\);
    
    \line1[34]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[34]_net_1\);
    
    \line3[19]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[19]_net_1\);
    
    \line2_RNIAA7P[21]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[21]_net_1\, B => \line2[21]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[21]\);
    
    \line7[57]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[57]_net_1\);
    
    \line4[28]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[28]_net_1\);
    
    \line1[31]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[31]_net_1\);
    
    \line5[58]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[58]_net_1\);
    
    \line4[10]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[10]_net_1\);
    
    \line4_RNIG4GB1[27]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[27]_net_1\, B => \line4[27]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[27]\);
    
    \line2[56]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[56]_net_1\);
    
    \line5[47]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[47]_net_1\);
    
    \line0_RNIVP271[24]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line1[24]_net_1\, B => \line0[24]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_7_1_1[24]\);
    
    \line4[3]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[3]_net_1\);
    
    \line2_RNI7UGH[12]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[12]_net_1\, B => \line2[12]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[12]\);
    
    \line2_RNIV56K[30]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line2[30]_net_1\, B => \line3[30]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_14_1_1[30]\);
    
    raddr_pos_0_rep1 : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_0_rep1\);
    
    \line6[26]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[26]_net_1\);
    
    \line5_or[32]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line5_0, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line5_or[32]_net_1\);
    
    \line0[26]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[26]_net_1\);
    
    \line0_RNINES82[59]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[27]\, C => \line1[59]_net_1\, D => 
        \line0[59]_net_1\, Y => N_946);
    
    \line1[15]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[15]_net_1\);
    
    \line6[49]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[49]_net_1\);
    
    \line6[13]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[13]_net_1\);
    
    \line1[63]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[63]_net_1\);
    
    \line2_RNI9IGE1[2]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[2]_net_1\, B => \line2[2]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[2]\);
    
    \line6_RNIB8AP[15]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[15]_net_1\, B => \line6[15]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[15]\);
    
    \line4_RNIG84F1[35]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[3]\, C => \line5[35]_net_1\, D => 
        \line4[35]_net_1\, Y => N_1402);
    
    \line2[54]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[54]_net_1\);
    
    \line2[26]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[26]_net_1\);
    
    \line6_RNI5VN61[48]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[16]\, C => \line7[48]_net_1\, D => 
        \line6[48]_net_1\, Y => N_1639);
    
    \line2_RNI3ARN[24]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line3[24]_net_1\, B => \line2[24]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_14_1_1[24]\);
    
    \line4[47]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[47]_net_1\);
    
    \line6[24]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[24]_net_1\);
    
    \line0_RNI2AA32[33]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[1]\, 
        C => \line1[33]_net_1\, D => \line0[33]_net_1\, Y => 
        N_920);
    
    data_available : SLE
      port map(D => N_12_0_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \SHA256_Module_0_data_available\);
    
    \line0[24]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[24]_net_1\);
    
    \line4_RNI7EUB[5]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[5]_net_1\, B => \line5[5]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[5]\);
    
    \line2[51]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[51]_net_1\);
    
    \line7[23]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[23]_net_1\);
    
    \raddr_pos_RNIHR1A3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_930, D => N_1154, Y => 
        \data_out_31_1_1[11]\);
    
    \line6[21]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[21]_net_1\);
    
    \line4[37]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[37]_net_1\);
    
    \line2[37]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[37]_net_1\);
    
    \line0_RNIIMSR1[47]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[15]\, 
        C => \line1[47]_net_1\, D => \line0[47]_net_1\, Y => 
        N_934);
    
    \raddr_pos_RNIK96D7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1643, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[20]\, D => N_1419, Y => N_1707);
    
    \line4[56]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[56]_net_1\);
    
    \line2[24]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[24]_net_1\);
    
    \line0[21]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[21]_net_1\);
    
    \line7[9]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[9]_net_1\);
    
    \line7[43]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[43]_net_1\);
    
    \line0_RNIRAES1[45]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[13]\, 
        C => \line1[45]_net_1\, D => \line0[45]_net_1\, Y => 
        N_932);
    
    \line6_RNI5KAG[2]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[2]_net_1\, B => \line7[2]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[2]\);
    
    \line6[59]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[59]_net_1\);
    
    \line0_RNIJA652[37]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_7_1_1[5]\, 
        C => \line1[37]_net_1\, D => \line0[37]_net_1\, Y => 
        N_924);
    
    \line5[12]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[12]_net_1\);
    
    \line0_RNI9OK32[53]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[21]\, 
        C => \line1[53]_net_1\, D => \line0[53]_net_1\, Y => 
        N_940);
    
    \line2_RNIR6BQ1[37]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[5]\, 
        C => \line3[37]_net_1\, D => \line2[37]_net_1\, Y => 
        N_1148);
    
    \line2_or[32]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line2_0, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line2_or[32]_net_1\);
    
    \line6_RNIHJBG1[59]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[27]\, C => \line7[59]_net_1\, D => 
        \line6[59]_net_1\, Y => N_1650);
    
    \raddr_pos_RNI367B3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_936, D => N_1160, Y => 
        \data_out_31_1_1[17]\);
    
    \line2[21]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[21]_net_1\);
    
    \line0[17]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[17]_net_1\);
    
    \line2_RNII2DA1[56]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[24]\, C => \line3[56]_net_1\, D => 
        \line2[56]_net_1\, Y => N_1167);
    
    \line1[55]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[55]_net_1\);
    
    \line3[35]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[35]_net_1\);
    
    \line6_RNIC6N61[42]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[10]\, C => \line7[42]_net_1\, D => 
        \line6[42]_net_1\, Y => N_1633);
    
    \line6_RNIQUID1[63]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[31]\, C => \line7[63]_net_1\, D => 
        \line6[63]_net_1\, Y => N_1654);
    
    \line4[54]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[54]_net_1\);
    
    \line0[55]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[55]_net_1\);
    
    \line5[3]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[3]_net_1\);
    
    \line7[36]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[36]_net_1\);
    
    \line6[18]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[18]_net_1\);
    
    raddr_pos_1_rep1 : SLE
      port map(D => sha256_controller_0_read_addr_0(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_1_rep1\);
    
    \line6_RNIPIN61[45]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[13]\, C => \line7[45]_net_1\, D => 
        \line6[45]_net_1\, Y => N_1636);
    
    \line6_RNIEE8S[24]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[24]_net_1\, B => \line6[24]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[24]\);
    
    \line4[51]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[51]_net_1\);
    
    \raddr_pos_RNIR8AG4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_925, D => N_1149, Y => 
        \data_out_31_1_1[6]\);
    
    \line4_RNIJM852[50]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[18]\, C => \line5[50]_net_1\, D => 
        \line4[50]_net_1\, Y => N_1417);
    
    \raddr_pos_fast_fast[0]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_fast_fast[0]_net_1\);
    
    \line5[30]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[30]_net_1\);
    
    \line2_RNIJRVT[49]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[17]\, C => \line3[49]_net_1\, D => 
        \line2[49]_net_1\, Y => N_1160);
    
    \line7[34]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[34]_net_1\);
    
    \line7[28]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[28]_net_1\);
    
    \line4_RNI1BQE2[57]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[25]\, C => \line5[57]_net_1\, D => 
        \line4[57]_net_1\, Y => N_1424);
    
    \line6[61]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[61]_net_1\);
    
    \line4_RNIIU1C2[63]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[31]\, C => \line5[63]_net_1\, D => 
        \line4[63]_net_1\, Y => N_1430);
    
    \line2_RNI5SGH[11]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[11]_net_1\, B => \line2[11]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[11]\);
    
    \raddr_pos[0]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos[0]_net_1\);
    
    \line7[48]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[48]_net_1\);
    
    \line2_RNISU2I[14]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[14]_net_1\, B => \line2[14]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[14]\);
    
    \line3[59]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[59]_net_1\);
    
    \line7[31]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[31]_net_1\);
    
    \line2[15]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[15]_net_1\);
    
    \line4_RNI5CUB[4]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[4]_net_1\, B => \line5[4]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[4]\);
    
    \line2[42]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[42]_net_1\);
    
    \line4_RNIVFH81[11]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[11]_net_1\, B => \line4[11]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[11]\);
    
    \raddr_pos_RNIRGT34[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_927, D => N_1151, Y => 
        \data_out_31_1_1[8]\);
    
    \line4_RNIC44F1[34]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[2]\, C => \line5[34]_net_1\, D => 
        \line4[34]_net_1\, Y => N_1401);
    
    \line2_RNI62DT[42]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[10]\, C => \line3[42]_net_1\, D => 
        \line2[42]_net_1\, Y => N_1153);
    
    \line1_or[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line1_0_62, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line1_or[0]_net_1\);
    
    \line3[22]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[22]_net_1\);
    
    \line0_RNIMCA11[13]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[13]_net_1\, B => \line0[13]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[13]\);
    
    \line5[0]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[0]_net_1\);
    
    \line4_RNI3KH81[13]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[13]_net_1\, B => \line4[13]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[13]\);
    
    \line6_RNITMN61[46]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[14]\, C => \line7[46]_net_1\, D => 
        \line6[46]_net_1\, Y => N_1637);
    
    \line4_RNIVASE2[61]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[29]\, C => \line5[61]_net_1\, D => 
        \line4[61]_net_1\, Y => N_1428);
    
    \line3[17]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[17]_net_1\);
    
    \line6_RNIS8941[36]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[4]\, C => \line7[36]_net_1\, D => 
        \line6[36]_net_1\, Y => N_1627);
    
    \line4_RNI13752[49]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[17]\, C => \line5[49]_net_1\, D => 
        \line4[49]_net_1\, Y => N_1416);
    
    \line4_RNI4S3F1[32]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[0]\, C => \line5[32]_net_1\, D => 
        \line4[32]_net_1\, Y => N_1399);
    
    \line6[36]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[36]_net_1\);
    
    \line0[42]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[42]_net_1\);
    
    \line4_RNIEMTB2[53]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[21]\, C => \line5[53]_net_1\, D => 
        \line4[53]_net_1\, Y => N_1420);
    
    \line2[5]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[5]_net_1\);
    
    \line1[39]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[39]_net_1\);
    
    \line5[13]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[13]_net_1\);
    
    \line6_RNITM9N[8]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line7[8]_net_1\, B => \line6[8]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_29_1_1[8]\);
    
    \line4[26]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[26]_net_1\);
    
    \line4[15]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[15]_net_1\);
    
    m35 : CFG4
      generic map(INIT => x"20A8")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_30, D => CertificationSystem_sb_0_GPIO_9_M2F, Y => 
        line0_0);
    
    \line2_RNIM6O61[61]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[29]\, C => \line3[61]_net_1\, D => 
        \line2[61]_net_1\, Y => N_1172);
    
    \line4_RNILM652[46]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[14]\, C => \line5[46]_net_1\, D => 
        \line4[46]_net_1\, Y => N_1413);
    
    \line5[56]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[56]_net_1\);
    
    \line6_RNI4H941[38]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[6]\, C => \line7[38]_net_1\, D => 
        \line6[38]_net_1\, Y => N_1629);
    
    \line6[47]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[47]_net_1\);
    
    \line6[34]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[34]_net_1\);
    
    \line2[62]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[62]_net_1\);
    
    \line0_RNI0NA11[18]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[18]_net_1\, B => \line0[18]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[18]\);
    
    m38 : CFG4
      generic map(INIT => x"80F7")

      port map(A => waddr_in_net_0(2), B => waddr_in_net_0(3), C
         => N_13_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => N_39);
    
    m1 : CFG2
      generic map(INIT => x"8")

      port map(A => CertificationSystem_sb_0_GPIO_1_M2F, B => 
        CertificationSystem_sb_0_GPIO_9_M2F, Y => 
        data_out_ready_0_sqmuxa);
    
    \line4_RNIDE652[44]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[12]\, C => \line5[44]_net_1\, D => 
        \line4[44]_net_1\, Y => N_1411);
    
    \raddr_pos_RNI9J1A3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_929, D => N_1153, Y => 
        \data_out_31_1_1[10]\);
    
    \line1[1]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[1]_net_1\);
    
    \line6[31]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[31]_net_1\);
    
    \line4[24]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[24]_net_1\);
    
    \line6_RNI1RN61[47]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[15]\, C => \line7[47]_net_1\, D => 
        \line6[47]_net_1\, Y => N_1638);
    
    \line5[54]\ : SLE
      port map(D => N_152_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[54]_net_1\);
    
    \line6_RNIDSAG[6]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[6]_net_1\, B => \line7[6]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[6]\);
    
    \line1[20]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[20]_net_1\);
    
    \line1[42]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[42]_net_1\);
    
    \line4[21]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[21]_net_1\);
    
    \line2[59]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[59]_net_1\);
    
    \raddr_pos_fast[0]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_fast[0]_net_1\);
    
    \line5[51]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[51]_net_1\);
    
    \line4_RNIIQTB2[54]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[22]\, C => \line5[54]_net_1\, D => 
        \line4[54]_net_1\, Y => N_1421);
    
    \line6[57]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[57]_net_1\);
    
    \line7[8]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[8]_net_1\);
    
    \raddr_pos_RNIRT6B3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_935, D => N_1159, Y => 
        \data_out_31_1_1[16]\);
    
    \line2_RNIFK4K[29]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line2[29]_net_1\, B => \line3[29]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_14_1_1[29]\);
    
    \line0[3]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[3]_net_1\);
    
    \line6[29]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[29]_net_1\);
    
    \raddr_pos_RNILSDB3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_939, D => N_1163, Y => 
        \data_out_31_1_1[20]\);
    
    \line0[29]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[29]_net_1\);
    
    \line3[42]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[42]_net_1\);
    
    \line5[18]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[18]_net_1\);
    
    \line0_RNIU1SR1[42]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[10]\, 
        C => \line1[42]_net_1\, D => \line0[42]_net_1\, Y => 
        N_929);
    
    \raddr_pos_RNI9SNS3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_948, D => N_1172, Y => 
        \data_out_31_1_1[29]\);
    
    \line4_RNI9GUB[6]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[6]_net_1\, B => \line5[6]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[6]\);
    
    \line2[43]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[43]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line2[29]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[29]_net_1\);
    
    \line6_RNI7MAG[3]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line6[3]_net_1\, B => \line7[3]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_29_1_1[3]\);
    
    \line0[30]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[30]_net_1\);
    
    \line3[23]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[23]_net_1\);
    
    \line7[62]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[62]_net_1\);
    
    \line1[5]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[5]_net_1\);
    
    \line4_RNI13IF1[41]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_22_1_1[9]\, 
        C => \line5[41]_net_1\, D => \line4[41]_net_1\, Y => 
        N_1408);
    
    \raddr_pos_RNI1K144[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_943, D => N_1167, Y => 
        \data_out_31_1_1[24]\);
    
    \line6[16]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[16]_net_1\);
    
    \line0[9]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[9]_net_1\);
    
    \line6_RNI8AAS[30]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[30]_net_1\, B => \line6[30]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_29_1_1[30]\);
    
    \line0[4]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[4]_net_1\);
    
    \line0[43]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[43]_net_1\);
    
    \line5[2]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[2]_net_1\);
    
    \line4[59]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[59]_net_1\);
    
    \raddr_pos_RNIP6C67[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1641, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[18]\, D => N_1417, Y => N_1705);
    
    raddr_pos_0_rep2 : SLE
      port map(D => sha256_controller_0_read_addr_0(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_0_rep2\);
    
    \line3_or[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line3_0_62, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line3_or[0]_net_1\);
    
    m25 : CFG4
      generic map(INIT => x"80A2")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_23_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => line3_0);
    
    \line7[10]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[10]_net_1\);
    
    \line5[20]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[20]_net_1\);
    
    \line6_RNIJGAP[19]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[19]_net_1\, B => \line6[19]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[19]\);
    
    \line1[12]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[12]_net_1\);
    
    \line6_RNIGS841[33]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[1]\, C => \line7[33]_net_1\, D => 
        \line6[33]_net_1\, Y => N_1624);
    
    \line5[35]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[35]_net_1\);
    
    \raddr_pos[1]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos[1]_net_1\);
    
    \line3[57]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[57]_net_1\);
    
    \line6[3]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[3]_net_1\);
    
    \raddr_pos_RNISCB04[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_946, D => N_1170, Y => 
        \data_out_31_1_1[27]\);
    
    \line0[5]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[5]_net_1\);
    
    m28 : CFG4
      generic map(INIT => x"20A8")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_23_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => line2_0);
    
    \line4_RNIOURB2[51]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[19]\, C => \line5[51]_net_1\, D => 
        \line4[51]_net_1\, Y => N_1418);
    
    \line7[26]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[26]_net_1\);
    
    \line6[14]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[14]_net_1\);
    
    \line2[63]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[63]_net_1\);
    
    \line2_RNIN2BQ1[36]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[4]\, 
        C => \line3[36]_net_1\, D => \line2[36]_net_1\, Y => 
        N_1147);
    
    \line2_RNI60LC1[1]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[1]_net_1\, B => \line2[1]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[1]\);
    
    \line0[2]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[2]_net_1\);
    
    \line7[50]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[50]_net_1\);
    
    \line2_RNI62FO1[32]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[0]\, 
        C => \line3[32]_net_1\, D => \line2[32]_net_1\, Y => 
        N_1143);
    
    \line7[46]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[46]_net_1\);
    
    \line7[39]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[39]_net_1\);
    
    \line0_RNI8UG81[31]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[31]_net_1\, B => \line0[31]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[31]\);
    
    \line0_RNIRLD31[30]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line0[30]_net_1\, B => \line1[30]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_7_1_1[30]\);
    
    \line6[11]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[11]_net_1\);
    
    \line1[61]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[61]_net_1\);
    
    \line5[40]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[40]_net_1\);
    
    \line2[48]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[48]_net_1\);
    
    \raddr_pos_RNIQNDE4[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_921, D => N_1145, Y => 
        \data_out_31_1_1[2]\);
    
    \line3[62]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[62]_net_1\);
    
    \line7[24]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[24]_net_1\);
    
    \line3[28]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[28]_net_1\);
    
    \line0_RNIK6IS1[52]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[20]\, 
        C => \line1[52]_net_1\, D => \line0[52]_net_1\, Y => 
        N_939);
    
    \line1[43]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[43]_net_1\);
    
    \line7[44]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[44]_net_1\);
    
    \line4[62]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[62]_net_1\);
    
    \line1[37]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[37]_net_1\);
    
    \raddr_pos_RNI3PT34[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_928, D => N_1152, Y => 
        \data_out_31_1_1[9]\);
    
    \line6_RNICO841[32]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[0]\, C => \line7[32]_net_1\, D => 
        \line6[32]_net_1\, Y => N_1623);
    
    \line7[21]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[21]_net_1\);
    
    \line0[48]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[48]_net_1\);
    
    \line0_RNIF6S82[57]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_7_1_1[25]\, C => \line1[57]_net_1\, D => 
        \line0[57]_net_1\, Y => N_944);
    
    \raddr_pos_RNI78JP3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_941, D => N_1165, Y => 
        \data_out_31_1_1[22]\);
    
    \line1[52]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[52]_net_1\);
    
    \line4[40]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[40]_net_1\);
    
    \line3[32]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[32]_net_1\);
    
    \line7[41]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[41]_net_1\);
    
    \line4_RNIAUFB1[24]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[24]_net_1\, B => \line4[24]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[24]\);
    
    \line0[52]\ : SLE
      port map(D => N_97_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[52]_net_1\);
    
    \line4_or[32]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line4_0, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line4_or[32]_net_1\);
    
    \line2_RNIS63U[52]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[20]\, C => \line3[52]_net_1\, D => 
        \line2[52]_net_1\, Y => N_1163);
    
    \line3[43]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[43]_net_1\);
    
    \line4_RNIE2GB1[26]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[26]_net_1\, B => \line4[26]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[26]\);
    
    raddr_pos_1_rep2 : SLE
      port map(D => sha256_controller_0_read_addr_0(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos_1_rep2\);
    
    \line0_RNIB4C31[29]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line0[29]_net_1\, B => \line1[29]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_7_1_1[29]\);
    
    \line4[30]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[30]_net_1\);
    
    \raddr_pos_RNI7DAB3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_937, D => N_1161, Y => 
        \data_out_31_1_1[18]\);
    
    \line2[30]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[30]_net_1\);
    
    \raddr_pos_RNIGKIV6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1640, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[17]\, D => N_1416, Y => N_1704);
    
    \line1[6]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[6]_net_1\);
    
    \raddr_pos_RNIGIGV6[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1636, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[13]\, D => N_1412, Y => N_1700);
    
    \line2_RNID4HH[15]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[15]_net_1\, B => \line2[15]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[15]\);
    
    \line0_RNI3EO01[12]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[12]_net_1\, B => \line0[12]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[12]\);
    
    \line7[63]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[63]_net_1\);
    
    \line4_RNIPATI[8]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line5[8]_net_1\, B => \line4[8]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_22_1_1[8]\);
    
    \line4_RNITU652[48]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_22_1_1[16]\, C => \line5[48]_net_1\, D => 
        \line4[48]_net_1\, Y => N_1415);
    
    \line6[39]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[39]_net_1\);
    
    \line0[10]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[10]_net_1\);
    
    \line4[5]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[5]_net_1\);
    
    \line2_RNI3QGH[10]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[10]_net_1\, B => \line2[10]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[10]\);
    
    \line2[57]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[57]_net_1\);
    
    \line2[0]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[0]_net_1\);
    
    \line1[25]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[25]_net_1\);
    
    \line4[2]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[2]_net_1\);
    
    \line6[27]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[27]_net_1\);
    
    \line4[29]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[29]_net_1\);
    
    \line1[48]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[48]_net_1\);
    
    \line1[13]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[13]_net_1\);
    
    \line2[12]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[12]_net_1\);
    
    \line0[27]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[27]_net_1\);
    
    \line5[59]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[59]_net_1\);
    
    \line0_RNI1CO01[11]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[11]_net_1\, B => \line0[11]_net_1\, C
         => \raddr_pos_fast_fast[0]_net_1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[11]\);
    
    m31 : CFG4
      generic map(INIT => x"4051")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_30, D => CertificationSystem_sb_0_GPIO_9_M2F, Y => 
        line1_0_62);
    
    \line2_RNI033I[16]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[16]_net_1\, B => \line2[16]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_14_1_1[16]\);
    
    \raddr_pos_RNIIQD48[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1652, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[29]\, D => N_1428, Y => N_1716);
    
    m17 : CFG4
      generic map(INIT => x"80A2")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_15_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => line5_0);
    
    \line2[27]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[27]_net_1\);
    
    \line2_RNIVABQ1[38]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[6]\, 
        C => \line3[38]_net_1\, D => \line2[38]_net_1\, Y => 
        N_1149);
    
    \raddr_pos_RNIPRT78[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1650, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[27]\, D => N_1426, Y => N_1714);
    
    \line2_RNI3FBQ1[39]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[7]\, 
        C => \line3[39]_net_1\, D => \line2[39]_net_1\, Y => 
        N_1150);
    
    \line3[48]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[48]_net_1\);
    
    \line6[7]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[7]_net_1\);
    
    \raddr_pos_RNI356B3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_932, D => N_1156, Y => 
        \data_out_31_1_1[13]\);
    
    \line5[16]\ : SLE
      port map(D => N_140_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[16]_net_1\);
    
    \line3_or[32]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line3_0, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line3_or[32]_net_1\);
    
    \raddr_pos_RNIBRVC7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1642, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[19]\, D => N_1418, Y => N_1706);
    
    \line0[35]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[35]_net_1\);
    
    \line0_RNIBRES1[49]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[17]\, 
        C => \line1[49]_net_1\, D => \line0[49]_net_1\, Y => 
        N_936);
    
    \line3[63]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[63]_net_1\);
    
    \line4[57]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[57]_net_1\);
    
    \line2_RNII2O61[60]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[28]\, C => \line3[60]_net_1\, D => 
        \line2[60]_net_1\, Y => N_1171);
    
    \line0_RNIOEA11[14]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[14]_net_1\, B => \line0[14]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[14]\);
    
    \line4[12]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[12]_net_1\);
    
    \line0_or[32]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line0_0, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line0_or[32]_net_1\);
    
    \line4[63]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[63]_net_1\);
    
    \raddr_pos_RNIOQJB8[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1648, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[25]\, D => N_1424, Y => N_1712);
    
    \line5[14]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[14]_net_1\);
    
    \raddr_pos_RNIP32A3[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_931, D => N_1155, Y => 
        \data_out_31_1_1[12]\);
    
    \line1[53]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[53]_net_1\);
    
    \line7[15]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[15]_net_1\);
    
    \line4_RNI3AUB[3]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \line4[3]_net_1\, B => \line5[3]_net_1\, C
         => \raddr_pos_0_rep2\, D => \raddr_pos[1]_net_1\, Y => 
        \data_out_22_1_1[3]\);
    
    \line3[33]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[33]_net_1\);
    
    \line5[25]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[25]_net_1\);
    
    \line0_or[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => line0_0_62, B => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, Y => 
        \line0_or[0]_net_1\);
    
    \line3[10]\ : SLE
      port map(D => N_77_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[10]_net_1\);
    
    \line0[53]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[53]_net_1\);
    
    \line7[2]\ : SLE
      port map(D => N_110_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[2]_net_1\);
    
    \line1[18]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[18]_net_1\);
    
    \line5[11]\ : SLE
      port map(D => N_83_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[11]_net_1\);
    
    \raddr_pos_RNIUM4C7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1629, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[6]\, D => N_1405, Y => N_1693);
    
    \raddr_pos_RNIM5CR7[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1645, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[22]\, D => N_1421, Y => N_1709);
    
    \raddr_pos_RNIJ4244[2]\ : CFG4
      generic map(INIT => x"2367")

      port map(A => \raddr_pos[3]_net_1\, B => 
        \raddr_pos[2]_net_1\, C => N_945, D => N_1169, Y => 
        \data_out_31_1_1[26]\);
    
    \line7[37]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[37]_net_1\);
    
    \line6_RNIDFBG1[58]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_29_1_1[26]\, C => \line7[58]_net_1\, D => 
        \line6[58]_net_1\, Y => N_1649);
    
    \line6_RNI98CP[23]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[23]_net_1\, B => \line6[23]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[23]\);
    
    \line7[55]\ : SLE
      port map(D => N_101_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[55]_net_1\);
    
    \line8[28]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line8_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        reg_17x32_0_last_word(0));
    
    \raddr_pos_RNISJA87[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1623, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[0]\, D => N_1399, Y => N_1687);
    
    \line1[3]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[3]_net_1\);
    
    \line5[45]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[45]_net_1\);
    
    \line6[19]\ : SLE
      port map(D => N_95_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[19]_net_1\);
    
    \line6[40]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[40]_net_1\);
    
    \line2[46]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[46]_net_1\);
    
    \line0_RNIBC4A1[5]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[5]_net_1\, B => \line0[5]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[5]\);
    
    \raddr_pos[2]\ : SLE
      port map(D => sha256_controller_0_read_addr_0(2), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_3_0, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => 
        CertificationSystem_sb_0_GPIO_9_M2F, SD => GND_net_1, LAT
         => GND_net_1, Q => \raddr_pos[2]_net_1\);
    
    \line4_RNI3OL81[31]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[31]_net_1\, B => \line4[31]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[31]\);
    
    \line0_RNISIA11[16]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[16]_net_1\, B => \line0[16]_net_1\, C
         => \raddr_pos_fast_0_rep1\, D => 
        \raddr_pos_fast[1]_net_1\, Y => \data_out_7_1_1[16]\);
    
    \line4_RNI1IH81[12]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[12]_net_1\, B => \line4[12]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_22_1_1[12]\);
    
    \line3[3]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[3]_net_1\);
    
    \line3[26]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[26]_net_1\);
    
    \line6_RNI93O61[49]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => 
        \data_out_29_1_1[17]\, C => \line7[49]_net_1\, D => 
        \line6[49]_net_1\, Y => N_1640);
    
    m9 : CFG4
      generic map(INIT => x"7555")

      port map(A => CertificationSystem_sb_0_GPIO_9_M2F, B => 
        CertificationSystem_sb_0_GPIO_1_M2F, C => 
        AHB_slave_dummy_0_write_en, D => N_49, Y => N_49_mux);
    
    \line6_RNI96AP[14]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[14]_net_1\, B => \line6[14]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[14]\);
    
    \line2[13]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[13]_net_1\);
    
    \line7[29]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[29]_net_1\);
    
    \line4[45]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[45]_net_1\);
    
    \line1[58]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[58]_net_1\);
    
    \line0[46]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[46]_net_1\);
    
    \line0[60]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[60]_net_1\);
    
    \line3[38]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[38]_net_1\);
    
    \line2[44]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[44]_net_1\);
    
    \line6_RNI76CP[22]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[22]_net_1\, B => \line6[22]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[22]\);
    
    \line7[49]\ : SLE
      port map(D => N_91_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line7_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line7[49]_net_1\);
    
    \line0[58]\ : SLE
      port map(D => N_103_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[58]_net_1\);
    
    \line4_RNIC0GB1[25]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[25]_net_1\, B => \line4[25]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[25]\);
    
    \line0[7]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[7]_net_1\);
    
    \line6[50]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[50]_net_1\);
    
    \line3[24]\ : SLE
      port map(D => N_156_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[24]_net_1\);
    
    \line2_RNIN6DA1[57]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_14_1_1[25]\, C => \line3[57]_net_1\, D => 
        \line2[57]_net_1\, Y => N_1168);
    
    \line4[35]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[35]_net_1\);
    
    \line6[9]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[9]_net_1\);
    
    \line2[41]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[41]_net_1\);
    
    \line2[35]\ : SLE
      port map(D => N_112_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[35]_net_1\);
    
    \line0_RNI7NES1[48]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[16]\, 
        C => \line1[48]_net_1\, D => \line0[48]_net_1\, Y => 
        N_935);
    
    \line6[37]\ : SLE
      port map(D => N_116_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[37]_net_1\);
    
    \raddr_pos_RNI0JI07[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1631, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[8]\, D => N_1407, Y => N_1695);
    
    \line0[44]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[44]_net_1\);
    
    \line3[21]\ : SLE
      port map(D => N_99_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[21]_net_1\);
    
    \line4_RNI804F1[33]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos[0]_net_1\, B => 
        \data_out_22_1_1[1]\, C => \line5[33]_net_1\, D => 
        \line4[33]_net_1\, Y => N_1400);
    
    \line5[32]\ : SLE
      port map(D => N_65_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[32]_net_1\);
    
    \line4[13]\ : SLE
      port map(D => N_133_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[13]_net_1\);
    
    \line2_RNIVU4K1[40]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_fast[0]_net_1\, B => 
        \data_out_14_1_1[8]\, C => \line3[40]_net_1\, D => 
        \line2[40]_net_1\, Y => N_1151);
    
    \line0[15]\ : SLE
      port map(D => N_89_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[15]_net_1\);
    
    \line2_RNIA6FO1[33]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_14_1_1[1]\, 
        C => \line3[33]_net_1\, D => \line2[33]_net_1\, Y => 
        N_1144);
    
    \line2_RNIA6DT[43]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[11]\, C => \line3[43]_net_1\, D => 
        \line2[43]_net_1\, Y => N_1154);
    
    \line4[27]\ : SLE
      port map(D => N_105_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[27]_net_1\);
    
    data_out_ready_1 : CFG4
      generic map(INIT => x"CDCC")

      port map(A => N_3_0, B => data_out_ready_0_sqmuxa, C => 
        AHB_slave_dummy_0_write_en, D => data_out_ready_net_1, Y
         => \data_out_ready_1\);
    
    \line5[6]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[6]_net_1\);
    
    \line5[57]\ : SLE
      port map(D => N_158_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[57]_net_1\);
    
    \line0[41]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[41]_net_1\);
    
    \line3[6]\ : SLE
      port map(D => N_69_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[6]_net_1\);
    
    \line0_RNI0I881[0]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line1[0]_net_1\, B => \line0[0]_net_1\, C
         => \raddr_pos_fast_0_rep2\, D => \raddr_pos_1_rep1\, Y
         => \data_out_7_1_1[0]\);
    
    \line6_RNI0U9P[10]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[10]_net_1\, B => \line6[10]_net_1\, C
         => \raddr_pos_1_rep1\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[10]\);
    
    \line8[30]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line8_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        reg_17x32_0_last_word(2));
    
    \raddr_pos_RNI1DBT6[3]\ : CFG4
      generic map(INIT => x"E323")

      port map(A => N_1632, B => \data_out_31_1_1[9]\, C => 
        \raddr_pos[3]_net_1\, D => N_1408, Y => N_1696);
    
    \line2[18]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[18]_net_1\);
    
    \raddr_pos_RNIQ8K48[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_1653, B => \raddr_pos[3]_net_1\, C => 
        \data_out_31_1_1[30]\, D => N_1429, Y => N_1717);
    
    \line1[46]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[46]_net_1\);
    
    m41 : CFG4
      generic map(INIT => x"80A2")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_39, D => CertificationSystem_sb_0_GPIO_9_M2F, Y => 
        line7_0);
    
    m12 : CFG4
      generic map(INIT => x"5755")

      port map(A => CertificationSystem_sb_0_GPIO_9_M2F, B => 
        CertificationSystem_sb_0_GPIO_1_M2F, C => 
        waddr_in_net_0(4), D => AHB_slave_dummy_0_write_en, Y => 
        N_13_0);
    
    m19 : CFG4
      generic map(INIT => x"1054")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_15_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => line4_0_62);
    
    \line2[61]\ : SLE
      port map(D => N_168_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[61]_net_1\);
    
    \line5[7]\ : SLE
      port map(D => N_71_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[7]_net_1\);
    
    \line6[8]\ : SLE
      port map(D => N_73_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line6_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line6[8]_net_1\);
    
    \line2_RNIFOGE1[5]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[5]_net_1\, B => \line2[5]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[5]\);
    
    \line2[9]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line2_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line2[9]_net_1\);
    
    \line0[1]\ : SLE
      port map(D => N_67_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line0_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line0[1]_net_1\);
    
    \line3[50]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[50]_net_1\);
    
    \line3[46]\ : SLE
      port map(D => N_87_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[46]_net_1\);
    
    \line5[60]\ : SLE
      port map(D => N_107_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line5_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line5[60]_net_1\);
    
    \line1[44]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[44]_net_1\);
    
    \line6_RNI78EP[31]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line7[31]_net_1\, B => \line6[31]_net_1\, C
         => \raddr_pos_1_rep2\, D => \raddr_pos_0_rep1\, Y => 
        \data_out_29_1_1[31]\);
    
    \line4_RNI4QHB1[30]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \line5[30]_net_1\, B => \line4[30]_net_1\, C
         => \raddr_pos[1]_net_1\, D => \raddr_pos[0]_net_1\, Y
         => \data_out_22_1_1[30]\);
    
    \line0_RNITEGS1[50]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => \data_out_7_1_1[18]\, 
        C => \line1[50]_net_1\, D => \line0[50]_net_1\, Y => 
        N_937);
    
    \line6_RNIQ8F11[41]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep2\, B => \data_out_29_1_1[9]\, 
        C => \line7[41]_net_1\, D => \line6[41]_net_1\, Y => 
        N_1632);
    
    \line2_RNIAJ1U[51]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => \raddr_pos_0_rep1\, B => 
        \data_out_14_1_1[19]\, C => \line3[51]_net_1\, D => 
        \line2[51]_net_1\, Y => N_1162);
    
    \line1[41]\ : SLE
      port map(D => N_75_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[41]_net_1\);
    
    \line4[18]\ : SLE
      port map(D => N_93_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line4_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line4[18]_net_1\);
    
    m20 : CFG4
      generic map(INIT => x"20A8")

      port map(A => waddr_in_net_0(0), B => waddr_in_net_0(1), C
         => N_15_0, D => CertificationSystem_sb_0_GPIO_9_M2F, Y
         => line4_0);
    
    \line2_RNIBKGE1[3]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \line3[3]_net_1\, B => \line2[3]_net_1\, C
         => \raddr_pos_fast[0]_net_1\, D => \raddr_pos_1_rep1\, Y
         => \data_out_14_1_1[3]\);
    
    data_available_RNO : CFG4
      generic map(INIT => x"BAFE")

      port map(A => \SHA256_Module_0_data_available\, B => 
        waddr_in_net_0(0), C => N_49_mux, D => 
        CertificationSystem_sb_0_GPIO_9_M2F, Y => N_12_0_i_0);
    
    \line3[44]\ : SLE
      port map(D => N_85_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line3_or[32]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line3[44]_net_1\);
    
    \line1[4]\ : SLE
      port map(D => N_114_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \line1_or[0]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => CertificationSystem_sb_0_GPIO_9_M2F, SD => 
        GND_net_1, LAT => GND_net_1, Q => \line1[4]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity SHA256_BLOCK is

    port( SHA256_BLOCK_0_H0_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o                       : out   std_logic_vector(31 downto 0);
          waddr_in_net_0                            : in    std_logic_vector(4 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0      : in    std_logic;
          SHA256_Module_0_di_req_o                  : out   std_logic;
          SHA256_BLOCK_0_do_valid_o                 : out   std_logic;
          SHA256_Module_0_waiting_data              : out   std_logic;
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic;
          SHA256_Module_0_error_o                   : out   std_logic;
          SHA256_BLOCK_0_start_o                    : out   std_logic;
          data_out_ready                            : out   std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F       : in    std_logic;
          SHA256_Module_0_data_available            : out   std_logic;
          N_111_i_0                                 : in    std_logic;
          N_109_i_0                                 : in    std_logic;
          N_168_i_0                                 : in    std_logic;
          N_107_i_0                                 : in    std_logic;
          N_99_i_0                                  : in    std_logic;
          N_97_i_0                                  : in    std_logic;
          N_67_i_0                                  : in    std_logic;
          N_65_i_0                                  : in    std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F_i_0   : in    std_logic;
          N_105_i_0                                 : in    std_logic;
          N_103_i_0                                 : in    std_logic;
          N_158_i_0                                 : in    std_logic;
          N_156_i_0                                 : in    std_logic;
          N_101_i_0                                 : in    std_logic;
          N_152_i_0                                 : in    std_logic;
          N_95_i_0                                  : in    std_logic;
          N_93_i_0                                  : in    std_logic;
          N_91_i_0                                  : in    std_logic;
          N_140_i_0                                 : in    std_logic;
          N_89_i_0                                  : in    std_logic;
          N_87_i_0                                  : in    std_logic;
          N_133_i_0                                 : in    std_logic;
          N_85_i_0                                  : in    std_logic;
          N_83_i_0                                  : in    std_logic;
          N_77_i_0                                  : in    std_logic;
          N_75_i_0                                  : in    std_logic;
          N_73_i_0                                  : in    std_logic;
          N_71_i_0                                  : in    std_logic;
          N_69_i_0                                  : in    std_logic;
          N_116_i_0                                 : in    std_logic;
          N_114_i_0                                 : in    std_logic;
          N_112_i_0                                 : in    std_logic;
          N_110_i_0                                 : in    std_logic;
          CertificationSystem_sb_0_GPIO_1_M2F       : in    std_logic;
          AHB_slave_dummy_0_write_en                : in    std_logic
        );

end SHA256_BLOCK;

architecture DEF_ARCH of SHA256_BLOCK is 

  component sha256_controller
    port( sha256_controller_0_read_addr_0      : out   std_logic_vector(3 downto 0);
          reg_17x32_0_last_word                : in    std_logic_vector(3 downto 0) := (others => 'U');
          di_o_0                               : in    std_logic_vector(1 to 1) := (others => 'U');
          state_1                              : out   std_logic;
          state_4                              : out   std_logic;
          state_3                              : out   std_logic;
          sha256_controller_0_di_o_5           : out   std_logic;
          sha256_controller_0_di_o_3           : out   std_logic;
          sha256_controller_0_di_o_0           : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          CertificationSystem_sb_0_GPIO_9_M2F  : in    std_logic := 'U';
          SHA256_Module_0_waiting_data         : out   std_logic;
          bytes_sel                            : out   std_logic;
          N_484                                : out   std_logic;
          data_out_ready                       : in    std_logic := 'U';
          prev_sig                             : in    std_logic := 'U';
          prev_sig_0                           : in    std_logic := 'U';
          first_block                          : in    std_logic := 'U';
          SHA256_Module_0_di_req_o             : in    std_logic := 'U';
          SHA256_BLOCK_0_do_valid_o            : in    std_logic := 'U';
          N_1705                               : in    std_logic := 'U';
          N_1703                               : in    std_logic := 'U';
          N_1700                               : in    std_logic := 'U';
          SHA256_BLOCK_0_start_o               : out   std_logic
        );
  end component;

  component gv_sha256
    port( reg_17x32_0_valid_bytes_0                 : in    std_logic_vector(1 downto 0) := (others => 'U');
          di_o_0                                    : out   std_logic_vector(1 to 1);
          SHA256_BLOCK_0_H0_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o                       : out   std_logic_vector(31 downto 0);
          state_0                                   : in    std_logic := 'U';
          state_2                                   : in    std_logic := 'U';
          state_3                                   : in    std_logic := 'U';
          sha256_controller_0_di_o_3                : in    std_logic := 'U';
          sha256_controller_0_di_o_5                : in    std_logic := 'U';
          sha256_controller_0_di_o_0                : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0      : in    std_logic := 'U';
          SHA256_Module_0_di_req_o                  : out   std_logic;
          SHA256_BLOCK_0_do_valid_o                 : out   std_logic;
          SHA256_Module_0_waiting_data              : in    std_logic := 'U';
          SHA256_Module_0_data_available_lastbank_8 : in    std_logic := 'U';
          N_484                                     : in    std_logic := 'U';
          bytes_sel                                 : in    std_logic := 'U';
          SHA256_Module_0_error_o                   : out   std_logic;
          SHA256_BLOCK_0_start_o                    : in    std_logic := 'U';
          N_1702                                    : in    std_logic := 'U';
          N_1710                                    : in    std_logic := 'U';
          ren_pos                                   : in    std_logic := 'U';
          N_1690                                    : in    std_logic := 'U';
          N_1691                                    : in    std_logic := 'U';
          N_1693                                    : in    std_logic := 'U';
          N_1692                                    : in    std_logic := 'U';
          N_1718                                    : in    std_logic := 'U';
          N_1694                                    : in    std_logic := 'U';
          N_1698                                    : in    std_logic := 'U';
          N_1701                                    : in    std_logic := 'U';
          N_1696                                    : in    std_logic := 'U';
          N_1697                                    : in    std_logic := 'U';
          N_1695                                    : in    std_logic := 'U';
          N_1699                                    : in    std_logic := 'U';
          N_1707                                    : in    std_logic := 'U';
          N_1708                                    : in    std_logic := 'U';
          N_1709                                    : in    std_logic := 'U';
          N_1706                                    : in    std_logic := 'U';
          N_1704                                    : in    std_logic := 'U';
          N_1688                                    : in    std_logic := 'U';
          N_1687                                    : in    std_logic := 'U';
          N_1689                                    : in    std_logic := 'U';
          N_1713                                    : in    std_logic := 'U';
          N_1716                                    : in    std_logic := 'U';
          N_1712                                    : in    std_logic := 'U';
          N_1717                                    : in    std_logic := 'U';
          N_1715                                    : in    std_logic := 'U';
          N_1711                                    : in    std_logic := 'U';
          N_1714                                    : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component limiter_1cycle
    port( prev_sig                             : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          first_block                          : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component limiter_1cycle_0
    port( prev_sig                             : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          data_out_ready                       : in    std_logic := 'U'
        );
  end component;

  component reg_17x32
    port( reg_17x32_0_last_word                     : out   std_logic_vector(3 downto 0);
          reg_17x32_0_valid_bytes_0                 : out   std_logic_vector(1 downto 0);
          sha256_controller_0_read_addr_0           : in    std_logic_vector(3 downto 0) := (others => 'U');
          waddr_in_net_0                            : in    std_logic_vector(4 downto 0) := (others => 'U');
          data_out_ready                            : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0      : in    std_logic := 'U';
          CertificationSystem_sb_0_GPIO_9_M2F       : in    std_logic := 'U';
          SHA256_Module_0_data_available            : out   std_logic;
          ren_pos                                   : out   std_logic;
          N_111_i_0                                 : in    std_logic := 'U';
          N_109_i_0                                 : in    std_logic := 'U';
          N_168_i_0                                 : in    std_logic := 'U';
          N_107_i_0                                 : in    std_logic := 'U';
          N_99_i_0                                  : in    std_logic := 'U';
          N_97_i_0                                  : in    std_logic := 'U';
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic;
          N_67_i_0                                  : in    std_logic := 'U';
          first_block                               : out   std_logic;
          N_65_i_0                                  : in    std_logic := 'U';
          CertificationSystem_sb_0_GPIO_9_M2F_i_0   : in    std_logic := 'U';
          N_105_i_0                                 : in    std_logic := 'U';
          N_103_i_0                                 : in    std_logic := 'U';
          N_158_i_0                                 : in    std_logic := 'U';
          N_156_i_0                                 : in    std_logic := 'U';
          N_101_i_0                                 : in    std_logic := 'U';
          N_152_i_0                                 : in    std_logic := 'U';
          N_95_i_0                                  : in    std_logic := 'U';
          N_93_i_0                                  : in    std_logic := 'U';
          N_91_i_0                                  : in    std_logic := 'U';
          N_140_i_0                                 : in    std_logic := 'U';
          N_89_i_0                                  : in    std_logic := 'U';
          N_87_i_0                                  : in    std_logic := 'U';
          N_133_i_0                                 : in    std_logic := 'U';
          N_85_i_0                                  : in    std_logic := 'U';
          N_83_i_0                                  : in    std_logic := 'U';
          N_77_i_0                                  : in    std_logic := 'U';
          N_75_i_0                                  : in    std_logic := 'U';
          N_73_i_0                                  : in    std_logic := 'U';
          N_71_i_0                                  : in    std_logic := 'U';
          N_69_i_0                                  : in    std_logic := 'U';
          N_116_i_0                                 : in    std_logic := 'U';
          N_114_i_0                                 : in    std_logic := 'U';
          N_112_i_0                                 : in    std_logic := 'U';
          N_110_i_0                                 : in    std_logic := 'U';
          N_1687                                    : out   std_logic;
          N_1717                                    : out   std_logic;
          N_1690                                    : out   std_logic;
          N_1689                                    : out   std_logic;
          N_1688                                    : out   std_logic;
          N_1715                                    : out   std_logic;
          N_1713                                    : out   std_logic;
          N_1710                                    : out   std_logic;
          N_1701                                    : out   std_logic;
          N_1714                                    : out   std_logic;
          N_1712                                    : out   std_logic;
          N_1716                                    : out   std_logic;
          N_1700                                    : out   std_logic;
          N_1698                                    : out   std_logic;
          N_1697                                    : out   std_logic;
          N_1692                                    : out   std_logic;
          N_1691                                    : out   std_logic;
          N_1704                                    : out   std_logic;
          N_1694                                    : out   std_logic;
          N_1709                                    : out   std_logic;
          N_1708                                    : out   std_logic;
          N_1707                                    : out   std_logic;
          N_1718                                    : out   std_logic;
          N_1703                                    : out   std_logic;
          N_1696                                    : out   std_logic;
          N_1699                                    : out   std_logic;
          N_1705                                    : out   std_logic;
          N_1695                                    : out   std_logic;
          N_1693                                    : out   std_logic;
          N_1706                                    : out   std_logic;
          N_1702                                    : out   std_logic;
          N_1711                                    : out   std_logic;
          CertificationSystem_sb_0_GPIO_1_M2F       : in    std_logic := 'U';
          AHB_slave_dummy_0_write_en                : in    std_logic := 'U'
        );
  end component;

    signal \reg_17x32_0_valid_bytes_0[0]\, 
        \reg_17x32_0_valid_bytes_0[1]\, \di_o_0[1]\, \state[1]\, 
        \state[3]\, \state[4]\, \sha256_controller_0_di_o[16]\, 
        \sha256_controller_0_di_o[18]\, 
        \sha256_controller_0_di_o[13]\, 
        \SHA256_Module_0_di_req_o\, \SHA256_BLOCK_0_do_valid_o\, 
        \SHA256_Module_0_waiting_data\, 
        \SHA256_Module_0_data_available_lastbank_8\, N_484, 
        bytes_sel, \SHA256_BLOCK_0_start_o\, N_1702, N_1710, 
        ren_pos, N_1690, N_1691, N_1693, N_1692, N_1718, N_1694, 
        N_1698, N_1701, N_1696, N_1697, N_1695, N_1699, N_1707, 
        N_1708, N_1709, N_1706, N_1704, N_1688, N_1687, N_1689, 
        N_1713, N_1716, N_1712, N_1717, N_1715, N_1711, N_1714, 
        prev_sig, first_block, prev_sig_0, \data_out_ready\, 
        \reg_17x32_0_last_word[0]\, \reg_17x32_0_last_word[1]\, 
        \reg_17x32_0_last_word[2]\, \reg_17x32_0_last_word[3]\, 
        \sha256_controller_0_read_addr_0[0]\, 
        \sha256_controller_0_read_addr_0[1]\, 
        \sha256_controller_0_read_addr_0[2]\, 
        \sha256_controller_0_read_addr_0[3]\, N_1700, N_1703, 
        N_1705, GND_net_1, VCC_net_1 : std_logic;

    for all : sha256_controller
	Use entity work.sha256_controller(DEF_ARCH);
    for all : gv_sha256
	Use entity work.gv_sha256(DEF_ARCH);
    for all : limiter_1cycle
	Use entity work.limiter_1cycle(DEF_ARCH);
    for all : limiter_1cycle_0
	Use entity work.limiter_1cycle_0(DEF_ARCH);
    for all : reg_17x32
	Use entity work.reg_17x32(DEF_ARCH);
begin 

    SHA256_Module_0_di_req_o <= \SHA256_Module_0_di_req_o\;
    SHA256_BLOCK_0_do_valid_o <= \SHA256_BLOCK_0_do_valid_o\;
    SHA256_Module_0_waiting_data <= 
        \SHA256_Module_0_waiting_data\;
    SHA256_Module_0_data_available_lastbank_8 <= 
        \SHA256_Module_0_data_available_lastbank_8\;
    SHA256_BLOCK_0_start_o <= \SHA256_BLOCK_0_start_o\;
    data_out_ready <= \data_out_ready\;

    sha256_controller_0 : sha256_controller
      port map(sha256_controller_0_read_addr_0(3) => 
        \sha256_controller_0_read_addr_0[3]\, 
        sha256_controller_0_read_addr_0(2) => 
        \sha256_controller_0_read_addr_0[2]\, 
        sha256_controller_0_read_addr_0(1) => 
        \sha256_controller_0_read_addr_0[1]\, 
        sha256_controller_0_read_addr_0(0) => 
        \sha256_controller_0_read_addr_0[0]\, 
        reg_17x32_0_last_word(3) => \reg_17x32_0_last_word[3]\, 
        reg_17x32_0_last_word(2) => \reg_17x32_0_last_word[2]\, 
        reg_17x32_0_last_word(1) => \reg_17x32_0_last_word[1]\, 
        reg_17x32_0_last_word(0) => \reg_17x32_0_last_word[0]\, 
        di_o_0(1) => \di_o_0[1]\, state_1 => \state[1]\, state_4
         => \state[4]\, state_3 => \state[3]\, 
        sha256_controller_0_di_o_5 => 
        \sha256_controller_0_di_o[18]\, 
        sha256_controller_0_di_o_3 => 
        \sha256_controller_0_di_o[16]\, 
        sha256_controller_0_di_o_0 => 
        \sha256_controller_0_di_o[13]\, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, 
        CertificationSystem_sb_0_GPIO_9_M2F => 
        CertificationSystem_sb_0_GPIO_9_M2F, 
        SHA256_Module_0_waiting_data => 
        \SHA256_Module_0_waiting_data\, bytes_sel => bytes_sel, 
        N_484 => N_484, data_out_ready => \data_out_ready\, 
        prev_sig => prev_sig_0, prev_sig_0 => prev_sig, 
        first_block => first_block, SHA256_Module_0_di_req_o => 
        \SHA256_Module_0_di_req_o\, SHA256_BLOCK_0_do_valid_o => 
        \SHA256_BLOCK_0_do_valid_o\, N_1705 => N_1705, N_1703 => 
        N_1703, N_1700 => N_1700, SHA256_BLOCK_0_start_o => 
        \SHA256_BLOCK_0_start_o\);
    
    gv_sha256_0 : gv_sha256
      port map(reg_17x32_0_valid_bytes_0(1) => 
        \reg_17x32_0_valid_bytes_0[1]\, 
        reg_17x32_0_valid_bytes_0(0) => 
        \reg_17x32_0_valid_bytes_0[0]\, di_o_0(1) => \di_o_0[1]\, 
        SHA256_BLOCK_0_H0_o(31) => SHA256_BLOCK_0_H0_o(31), 
        SHA256_BLOCK_0_H0_o(30) => SHA256_BLOCK_0_H0_o(30), 
        SHA256_BLOCK_0_H0_o(29) => SHA256_BLOCK_0_H0_o(29), 
        SHA256_BLOCK_0_H0_o(28) => SHA256_BLOCK_0_H0_o(28), 
        SHA256_BLOCK_0_H0_o(27) => SHA256_BLOCK_0_H0_o(27), 
        SHA256_BLOCK_0_H0_o(26) => SHA256_BLOCK_0_H0_o(26), 
        SHA256_BLOCK_0_H0_o(25) => SHA256_BLOCK_0_H0_o(25), 
        SHA256_BLOCK_0_H0_o(24) => SHA256_BLOCK_0_H0_o(24), 
        SHA256_BLOCK_0_H0_o(23) => SHA256_BLOCK_0_H0_o(23), 
        SHA256_BLOCK_0_H0_o(22) => SHA256_BLOCK_0_H0_o(22), 
        SHA256_BLOCK_0_H0_o(21) => SHA256_BLOCK_0_H0_o(21), 
        SHA256_BLOCK_0_H0_o(20) => SHA256_BLOCK_0_H0_o(20), 
        SHA256_BLOCK_0_H0_o(19) => SHA256_BLOCK_0_H0_o(19), 
        SHA256_BLOCK_0_H0_o(18) => SHA256_BLOCK_0_H0_o(18), 
        SHA256_BLOCK_0_H0_o(17) => SHA256_BLOCK_0_H0_o(17), 
        SHA256_BLOCK_0_H0_o(16) => SHA256_BLOCK_0_H0_o(16), 
        SHA256_BLOCK_0_H0_o(15) => SHA256_BLOCK_0_H0_o(15), 
        SHA256_BLOCK_0_H0_o(14) => SHA256_BLOCK_0_H0_o(14), 
        SHA256_BLOCK_0_H0_o(13) => SHA256_BLOCK_0_H0_o(13), 
        SHA256_BLOCK_0_H0_o(12) => SHA256_BLOCK_0_H0_o(12), 
        SHA256_BLOCK_0_H0_o(11) => SHA256_BLOCK_0_H0_o(11), 
        SHA256_BLOCK_0_H0_o(10) => SHA256_BLOCK_0_H0_o(10), 
        SHA256_BLOCK_0_H0_o(9) => SHA256_BLOCK_0_H0_o(9), 
        SHA256_BLOCK_0_H0_o(8) => SHA256_BLOCK_0_H0_o(8), 
        SHA256_BLOCK_0_H0_o(7) => SHA256_BLOCK_0_H0_o(7), 
        SHA256_BLOCK_0_H0_o(6) => SHA256_BLOCK_0_H0_o(6), 
        SHA256_BLOCK_0_H0_o(5) => SHA256_BLOCK_0_H0_o(5), 
        SHA256_BLOCK_0_H0_o(4) => SHA256_BLOCK_0_H0_o(4), 
        SHA256_BLOCK_0_H0_o(3) => SHA256_BLOCK_0_H0_o(3), 
        SHA256_BLOCK_0_H0_o(2) => SHA256_BLOCK_0_H0_o(2), 
        SHA256_BLOCK_0_H0_o(1) => SHA256_BLOCK_0_H0_o(1), 
        SHA256_BLOCK_0_H0_o(0) => SHA256_BLOCK_0_H0_o(0), 
        SHA256_BLOCK_0_H1_o(31) => SHA256_BLOCK_0_H1_o(31), 
        SHA256_BLOCK_0_H1_o(30) => SHA256_BLOCK_0_H1_o(30), 
        SHA256_BLOCK_0_H1_o(29) => SHA256_BLOCK_0_H1_o(29), 
        SHA256_BLOCK_0_H1_o(28) => SHA256_BLOCK_0_H1_o(28), 
        SHA256_BLOCK_0_H1_o(27) => SHA256_BLOCK_0_H1_o(27), 
        SHA256_BLOCK_0_H1_o(26) => SHA256_BLOCK_0_H1_o(26), 
        SHA256_BLOCK_0_H1_o(25) => SHA256_BLOCK_0_H1_o(25), 
        SHA256_BLOCK_0_H1_o(24) => SHA256_BLOCK_0_H1_o(24), 
        SHA256_BLOCK_0_H1_o(23) => SHA256_BLOCK_0_H1_o(23), 
        SHA256_BLOCK_0_H1_o(22) => SHA256_BLOCK_0_H1_o(22), 
        SHA256_BLOCK_0_H1_o(21) => SHA256_BLOCK_0_H1_o(21), 
        SHA256_BLOCK_0_H1_o(20) => SHA256_BLOCK_0_H1_o(20), 
        SHA256_BLOCK_0_H1_o(19) => SHA256_BLOCK_0_H1_o(19), 
        SHA256_BLOCK_0_H1_o(18) => SHA256_BLOCK_0_H1_o(18), 
        SHA256_BLOCK_0_H1_o(17) => SHA256_BLOCK_0_H1_o(17), 
        SHA256_BLOCK_0_H1_o(16) => SHA256_BLOCK_0_H1_o(16), 
        SHA256_BLOCK_0_H1_o(15) => SHA256_BLOCK_0_H1_o(15), 
        SHA256_BLOCK_0_H1_o(14) => SHA256_BLOCK_0_H1_o(14), 
        SHA256_BLOCK_0_H1_o(13) => SHA256_BLOCK_0_H1_o(13), 
        SHA256_BLOCK_0_H1_o(12) => SHA256_BLOCK_0_H1_o(12), 
        SHA256_BLOCK_0_H1_o(11) => SHA256_BLOCK_0_H1_o(11), 
        SHA256_BLOCK_0_H1_o(10) => SHA256_BLOCK_0_H1_o(10), 
        SHA256_BLOCK_0_H1_o(9) => SHA256_BLOCK_0_H1_o(9), 
        SHA256_BLOCK_0_H1_o(8) => SHA256_BLOCK_0_H1_o(8), 
        SHA256_BLOCK_0_H1_o(7) => SHA256_BLOCK_0_H1_o(7), 
        SHA256_BLOCK_0_H1_o(6) => SHA256_BLOCK_0_H1_o(6), 
        SHA256_BLOCK_0_H1_o(5) => SHA256_BLOCK_0_H1_o(5), 
        SHA256_BLOCK_0_H1_o(4) => SHA256_BLOCK_0_H1_o(4), 
        SHA256_BLOCK_0_H1_o(3) => SHA256_BLOCK_0_H1_o(3), 
        SHA256_BLOCK_0_H1_o(2) => SHA256_BLOCK_0_H1_o(2), 
        SHA256_BLOCK_0_H1_o(1) => SHA256_BLOCK_0_H1_o(1), 
        SHA256_BLOCK_0_H1_o(0) => SHA256_BLOCK_0_H1_o(0), 
        SHA256_BLOCK_0_H2_o(31) => SHA256_BLOCK_0_H2_o(31), 
        SHA256_BLOCK_0_H2_o(30) => SHA256_BLOCK_0_H2_o(30), 
        SHA256_BLOCK_0_H2_o(29) => SHA256_BLOCK_0_H2_o(29), 
        SHA256_BLOCK_0_H2_o(28) => SHA256_BLOCK_0_H2_o(28), 
        SHA256_BLOCK_0_H2_o(27) => SHA256_BLOCK_0_H2_o(27), 
        SHA256_BLOCK_0_H2_o(26) => SHA256_BLOCK_0_H2_o(26), 
        SHA256_BLOCK_0_H2_o(25) => SHA256_BLOCK_0_H2_o(25), 
        SHA256_BLOCK_0_H2_o(24) => SHA256_BLOCK_0_H2_o(24), 
        SHA256_BLOCK_0_H2_o(23) => SHA256_BLOCK_0_H2_o(23), 
        SHA256_BLOCK_0_H2_o(22) => SHA256_BLOCK_0_H2_o(22), 
        SHA256_BLOCK_0_H2_o(21) => SHA256_BLOCK_0_H2_o(21), 
        SHA256_BLOCK_0_H2_o(20) => SHA256_BLOCK_0_H2_o(20), 
        SHA256_BLOCK_0_H2_o(19) => SHA256_BLOCK_0_H2_o(19), 
        SHA256_BLOCK_0_H2_o(18) => SHA256_BLOCK_0_H2_o(18), 
        SHA256_BLOCK_0_H2_o(17) => SHA256_BLOCK_0_H2_o(17), 
        SHA256_BLOCK_0_H2_o(16) => SHA256_BLOCK_0_H2_o(16), 
        SHA256_BLOCK_0_H2_o(15) => SHA256_BLOCK_0_H2_o(15), 
        SHA256_BLOCK_0_H2_o(14) => SHA256_BLOCK_0_H2_o(14), 
        SHA256_BLOCK_0_H2_o(13) => SHA256_BLOCK_0_H2_o(13), 
        SHA256_BLOCK_0_H2_o(12) => SHA256_BLOCK_0_H2_o(12), 
        SHA256_BLOCK_0_H2_o(11) => SHA256_BLOCK_0_H2_o(11), 
        SHA256_BLOCK_0_H2_o(10) => SHA256_BLOCK_0_H2_o(10), 
        SHA256_BLOCK_0_H2_o(9) => SHA256_BLOCK_0_H2_o(9), 
        SHA256_BLOCK_0_H2_o(8) => SHA256_BLOCK_0_H2_o(8), 
        SHA256_BLOCK_0_H2_o(7) => SHA256_BLOCK_0_H2_o(7), 
        SHA256_BLOCK_0_H2_o(6) => SHA256_BLOCK_0_H2_o(6), 
        SHA256_BLOCK_0_H2_o(5) => SHA256_BLOCK_0_H2_o(5), 
        SHA256_BLOCK_0_H2_o(4) => SHA256_BLOCK_0_H2_o(4), 
        SHA256_BLOCK_0_H2_o(3) => SHA256_BLOCK_0_H2_o(3), 
        SHA256_BLOCK_0_H2_o(2) => SHA256_BLOCK_0_H2_o(2), 
        SHA256_BLOCK_0_H2_o(1) => SHA256_BLOCK_0_H2_o(1), 
        SHA256_BLOCK_0_H2_o(0) => SHA256_BLOCK_0_H2_o(0), 
        SHA256_BLOCK_0_H3_o(31) => SHA256_BLOCK_0_H3_o(31), 
        SHA256_BLOCK_0_H3_o(30) => SHA256_BLOCK_0_H3_o(30), 
        SHA256_BLOCK_0_H3_o(29) => SHA256_BLOCK_0_H3_o(29), 
        SHA256_BLOCK_0_H3_o(28) => SHA256_BLOCK_0_H3_o(28), 
        SHA256_BLOCK_0_H3_o(27) => SHA256_BLOCK_0_H3_o(27), 
        SHA256_BLOCK_0_H3_o(26) => SHA256_BLOCK_0_H3_o(26), 
        SHA256_BLOCK_0_H3_o(25) => SHA256_BLOCK_0_H3_o(25), 
        SHA256_BLOCK_0_H3_o(24) => SHA256_BLOCK_0_H3_o(24), 
        SHA256_BLOCK_0_H3_o(23) => SHA256_BLOCK_0_H3_o(23), 
        SHA256_BLOCK_0_H3_o(22) => SHA256_BLOCK_0_H3_o(22), 
        SHA256_BLOCK_0_H3_o(21) => SHA256_BLOCK_0_H3_o(21), 
        SHA256_BLOCK_0_H3_o(20) => SHA256_BLOCK_0_H3_o(20), 
        SHA256_BLOCK_0_H3_o(19) => SHA256_BLOCK_0_H3_o(19), 
        SHA256_BLOCK_0_H3_o(18) => SHA256_BLOCK_0_H3_o(18), 
        SHA256_BLOCK_0_H3_o(17) => SHA256_BLOCK_0_H3_o(17), 
        SHA256_BLOCK_0_H3_o(16) => SHA256_BLOCK_0_H3_o(16), 
        SHA256_BLOCK_0_H3_o(15) => SHA256_BLOCK_0_H3_o(15), 
        SHA256_BLOCK_0_H3_o(14) => SHA256_BLOCK_0_H3_o(14), 
        SHA256_BLOCK_0_H3_o(13) => SHA256_BLOCK_0_H3_o(13), 
        SHA256_BLOCK_0_H3_o(12) => SHA256_BLOCK_0_H3_o(12), 
        SHA256_BLOCK_0_H3_o(11) => SHA256_BLOCK_0_H3_o(11), 
        SHA256_BLOCK_0_H3_o(10) => SHA256_BLOCK_0_H3_o(10), 
        SHA256_BLOCK_0_H3_o(9) => SHA256_BLOCK_0_H3_o(9), 
        SHA256_BLOCK_0_H3_o(8) => SHA256_BLOCK_0_H3_o(8), 
        SHA256_BLOCK_0_H3_o(7) => SHA256_BLOCK_0_H3_o(7), 
        SHA256_BLOCK_0_H3_o(6) => SHA256_BLOCK_0_H3_o(6), 
        SHA256_BLOCK_0_H3_o(5) => SHA256_BLOCK_0_H3_o(5), 
        SHA256_BLOCK_0_H3_o(4) => SHA256_BLOCK_0_H3_o(4), 
        SHA256_BLOCK_0_H3_o(3) => SHA256_BLOCK_0_H3_o(3), 
        SHA256_BLOCK_0_H3_o(2) => SHA256_BLOCK_0_H3_o(2), 
        SHA256_BLOCK_0_H3_o(1) => SHA256_BLOCK_0_H3_o(1), 
        SHA256_BLOCK_0_H3_o(0) => SHA256_BLOCK_0_H3_o(0), 
        SHA256_BLOCK_0_H4_o(31) => SHA256_BLOCK_0_H4_o(31), 
        SHA256_BLOCK_0_H4_o(30) => SHA256_BLOCK_0_H4_o(30), 
        SHA256_BLOCK_0_H4_o(29) => SHA256_BLOCK_0_H4_o(29), 
        SHA256_BLOCK_0_H4_o(28) => SHA256_BLOCK_0_H4_o(28), 
        SHA256_BLOCK_0_H4_o(27) => SHA256_BLOCK_0_H4_o(27), 
        SHA256_BLOCK_0_H4_o(26) => SHA256_BLOCK_0_H4_o(26), 
        SHA256_BLOCK_0_H4_o(25) => SHA256_BLOCK_0_H4_o(25), 
        SHA256_BLOCK_0_H4_o(24) => SHA256_BLOCK_0_H4_o(24), 
        SHA256_BLOCK_0_H4_o(23) => SHA256_BLOCK_0_H4_o(23), 
        SHA256_BLOCK_0_H4_o(22) => SHA256_BLOCK_0_H4_o(22), 
        SHA256_BLOCK_0_H4_o(21) => SHA256_BLOCK_0_H4_o(21), 
        SHA256_BLOCK_0_H4_o(20) => SHA256_BLOCK_0_H4_o(20), 
        SHA256_BLOCK_0_H4_o(19) => SHA256_BLOCK_0_H4_o(19), 
        SHA256_BLOCK_0_H4_o(18) => SHA256_BLOCK_0_H4_o(18), 
        SHA256_BLOCK_0_H4_o(17) => SHA256_BLOCK_0_H4_o(17), 
        SHA256_BLOCK_0_H4_o(16) => SHA256_BLOCK_0_H4_o(16), 
        SHA256_BLOCK_0_H4_o(15) => SHA256_BLOCK_0_H4_o(15), 
        SHA256_BLOCK_0_H4_o(14) => SHA256_BLOCK_0_H4_o(14), 
        SHA256_BLOCK_0_H4_o(13) => SHA256_BLOCK_0_H4_o(13), 
        SHA256_BLOCK_0_H4_o(12) => SHA256_BLOCK_0_H4_o(12), 
        SHA256_BLOCK_0_H4_o(11) => SHA256_BLOCK_0_H4_o(11), 
        SHA256_BLOCK_0_H4_o(10) => SHA256_BLOCK_0_H4_o(10), 
        SHA256_BLOCK_0_H4_o(9) => SHA256_BLOCK_0_H4_o(9), 
        SHA256_BLOCK_0_H4_o(8) => SHA256_BLOCK_0_H4_o(8), 
        SHA256_BLOCK_0_H4_o(7) => SHA256_BLOCK_0_H4_o(7), 
        SHA256_BLOCK_0_H4_o(6) => SHA256_BLOCK_0_H4_o(6), 
        SHA256_BLOCK_0_H4_o(5) => SHA256_BLOCK_0_H4_o(5), 
        SHA256_BLOCK_0_H4_o(4) => SHA256_BLOCK_0_H4_o(4), 
        SHA256_BLOCK_0_H4_o(3) => SHA256_BLOCK_0_H4_o(3), 
        SHA256_BLOCK_0_H4_o(2) => SHA256_BLOCK_0_H4_o(2), 
        SHA256_BLOCK_0_H4_o(1) => SHA256_BLOCK_0_H4_o(1), 
        SHA256_BLOCK_0_H4_o(0) => SHA256_BLOCK_0_H4_o(0), 
        SHA256_BLOCK_0_H5_o(31) => SHA256_BLOCK_0_H5_o(31), 
        SHA256_BLOCK_0_H5_o(30) => SHA256_BLOCK_0_H5_o(30), 
        SHA256_BLOCK_0_H5_o(29) => SHA256_BLOCK_0_H5_o(29), 
        SHA256_BLOCK_0_H5_o(28) => SHA256_BLOCK_0_H5_o(28), 
        SHA256_BLOCK_0_H5_o(27) => SHA256_BLOCK_0_H5_o(27), 
        SHA256_BLOCK_0_H5_o(26) => SHA256_BLOCK_0_H5_o(26), 
        SHA256_BLOCK_0_H5_o(25) => SHA256_BLOCK_0_H5_o(25), 
        SHA256_BLOCK_0_H5_o(24) => SHA256_BLOCK_0_H5_o(24), 
        SHA256_BLOCK_0_H5_o(23) => SHA256_BLOCK_0_H5_o(23), 
        SHA256_BLOCK_0_H5_o(22) => SHA256_BLOCK_0_H5_o(22), 
        SHA256_BLOCK_0_H5_o(21) => SHA256_BLOCK_0_H5_o(21), 
        SHA256_BLOCK_0_H5_o(20) => SHA256_BLOCK_0_H5_o(20), 
        SHA256_BLOCK_0_H5_o(19) => SHA256_BLOCK_0_H5_o(19), 
        SHA256_BLOCK_0_H5_o(18) => SHA256_BLOCK_0_H5_o(18), 
        SHA256_BLOCK_0_H5_o(17) => SHA256_BLOCK_0_H5_o(17), 
        SHA256_BLOCK_0_H5_o(16) => SHA256_BLOCK_0_H5_o(16), 
        SHA256_BLOCK_0_H5_o(15) => SHA256_BLOCK_0_H5_o(15), 
        SHA256_BLOCK_0_H5_o(14) => SHA256_BLOCK_0_H5_o(14), 
        SHA256_BLOCK_0_H5_o(13) => SHA256_BLOCK_0_H5_o(13), 
        SHA256_BLOCK_0_H5_o(12) => SHA256_BLOCK_0_H5_o(12), 
        SHA256_BLOCK_0_H5_o(11) => SHA256_BLOCK_0_H5_o(11), 
        SHA256_BLOCK_0_H5_o(10) => SHA256_BLOCK_0_H5_o(10), 
        SHA256_BLOCK_0_H5_o(9) => SHA256_BLOCK_0_H5_o(9), 
        SHA256_BLOCK_0_H5_o(8) => SHA256_BLOCK_0_H5_o(8), 
        SHA256_BLOCK_0_H5_o(7) => SHA256_BLOCK_0_H5_o(7), 
        SHA256_BLOCK_0_H5_o(6) => SHA256_BLOCK_0_H5_o(6), 
        SHA256_BLOCK_0_H5_o(5) => SHA256_BLOCK_0_H5_o(5), 
        SHA256_BLOCK_0_H5_o(4) => SHA256_BLOCK_0_H5_o(4), 
        SHA256_BLOCK_0_H5_o(3) => SHA256_BLOCK_0_H5_o(3), 
        SHA256_BLOCK_0_H5_o(2) => SHA256_BLOCK_0_H5_o(2), 
        SHA256_BLOCK_0_H5_o(1) => SHA256_BLOCK_0_H5_o(1), 
        SHA256_BLOCK_0_H5_o(0) => SHA256_BLOCK_0_H5_o(0), 
        SHA256_BLOCK_0_H6_o(31) => SHA256_BLOCK_0_H6_o(31), 
        SHA256_BLOCK_0_H6_o(30) => SHA256_BLOCK_0_H6_o(30), 
        SHA256_BLOCK_0_H6_o(29) => SHA256_BLOCK_0_H6_o(29), 
        SHA256_BLOCK_0_H6_o(28) => SHA256_BLOCK_0_H6_o(28), 
        SHA256_BLOCK_0_H6_o(27) => SHA256_BLOCK_0_H6_o(27), 
        SHA256_BLOCK_0_H6_o(26) => SHA256_BLOCK_0_H6_o(26), 
        SHA256_BLOCK_0_H6_o(25) => SHA256_BLOCK_0_H6_o(25), 
        SHA256_BLOCK_0_H6_o(24) => SHA256_BLOCK_0_H6_o(24), 
        SHA256_BLOCK_0_H6_o(23) => SHA256_BLOCK_0_H6_o(23), 
        SHA256_BLOCK_0_H6_o(22) => SHA256_BLOCK_0_H6_o(22), 
        SHA256_BLOCK_0_H6_o(21) => SHA256_BLOCK_0_H6_o(21), 
        SHA256_BLOCK_0_H6_o(20) => SHA256_BLOCK_0_H6_o(20), 
        SHA256_BLOCK_0_H6_o(19) => SHA256_BLOCK_0_H6_o(19), 
        SHA256_BLOCK_0_H6_o(18) => SHA256_BLOCK_0_H6_o(18), 
        SHA256_BLOCK_0_H6_o(17) => SHA256_BLOCK_0_H6_o(17), 
        SHA256_BLOCK_0_H6_o(16) => SHA256_BLOCK_0_H6_o(16), 
        SHA256_BLOCK_0_H6_o(15) => SHA256_BLOCK_0_H6_o(15), 
        SHA256_BLOCK_0_H6_o(14) => SHA256_BLOCK_0_H6_o(14), 
        SHA256_BLOCK_0_H6_o(13) => SHA256_BLOCK_0_H6_o(13), 
        SHA256_BLOCK_0_H6_o(12) => SHA256_BLOCK_0_H6_o(12), 
        SHA256_BLOCK_0_H6_o(11) => SHA256_BLOCK_0_H6_o(11), 
        SHA256_BLOCK_0_H6_o(10) => SHA256_BLOCK_0_H6_o(10), 
        SHA256_BLOCK_0_H6_o(9) => SHA256_BLOCK_0_H6_o(9), 
        SHA256_BLOCK_0_H6_o(8) => SHA256_BLOCK_0_H6_o(8), 
        SHA256_BLOCK_0_H6_o(7) => SHA256_BLOCK_0_H6_o(7), 
        SHA256_BLOCK_0_H6_o(6) => SHA256_BLOCK_0_H6_o(6), 
        SHA256_BLOCK_0_H6_o(5) => SHA256_BLOCK_0_H6_o(5), 
        SHA256_BLOCK_0_H6_o(4) => SHA256_BLOCK_0_H6_o(4), 
        SHA256_BLOCK_0_H6_o(3) => SHA256_BLOCK_0_H6_o(3), 
        SHA256_BLOCK_0_H6_o(2) => SHA256_BLOCK_0_H6_o(2), 
        SHA256_BLOCK_0_H6_o(1) => SHA256_BLOCK_0_H6_o(1), 
        SHA256_BLOCK_0_H6_o(0) => SHA256_BLOCK_0_H6_o(0), 
        SHA256_BLOCK_0_H7_o(31) => SHA256_BLOCK_0_H7_o(31), 
        SHA256_BLOCK_0_H7_o(30) => SHA256_BLOCK_0_H7_o(30), 
        SHA256_BLOCK_0_H7_o(29) => SHA256_BLOCK_0_H7_o(29), 
        SHA256_BLOCK_0_H7_o(28) => SHA256_BLOCK_0_H7_o(28), 
        SHA256_BLOCK_0_H7_o(27) => SHA256_BLOCK_0_H7_o(27), 
        SHA256_BLOCK_0_H7_o(26) => SHA256_BLOCK_0_H7_o(26), 
        SHA256_BLOCK_0_H7_o(25) => SHA256_BLOCK_0_H7_o(25), 
        SHA256_BLOCK_0_H7_o(24) => SHA256_BLOCK_0_H7_o(24), 
        SHA256_BLOCK_0_H7_o(23) => SHA256_BLOCK_0_H7_o(23), 
        SHA256_BLOCK_0_H7_o(22) => SHA256_BLOCK_0_H7_o(22), 
        SHA256_BLOCK_0_H7_o(21) => SHA256_BLOCK_0_H7_o(21), 
        SHA256_BLOCK_0_H7_o(20) => SHA256_BLOCK_0_H7_o(20), 
        SHA256_BLOCK_0_H7_o(19) => SHA256_BLOCK_0_H7_o(19), 
        SHA256_BLOCK_0_H7_o(18) => SHA256_BLOCK_0_H7_o(18), 
        SHA256_BLOCK_0_H7_o(17) => SHA256_BLOCK_0_H7_o(17), 
        SHA256_BLOCK_0_H7_o(16) => SHA256_BLOCK_0_H7_o(16), 
        SHA256_BLOCK_0_H7_o(15) => SHA256_BLOCK_0_H7_o(15), 
        SHA256_BLOCK_0_H7_o(14) => SHA256_BLOCK_0_H7_o(14), 
        SHA256_BLOCK_0_H7_o(13) => SHA256_BLOCK_0_H7_o(13), 
        SHA256_BLOCK_0_H7_o(12) => SHA256_BLOCK_0_H7_o(12), 
        SHA256_BLOCK_0_H7_o(11) => SHA256_BLOCK_0_H7_o(11), 
        SHA256_BLOCK_0_H7_o(10) => SHA256_BLOCK_0_H7_o(10), 
        SHA256_BLOCK_0_H7_o(9) => SHA256_BLOCK_0_H7_o(9), 
        SHA256_BLOCK_0_H7_o(8) => SHA256_BLOCK_0_H7_o(8), 
        SHA256_BLOCK_0_H7_o(7) => SHA256_BLOCK_0_H7_o(7), 
        SHA256_BLOCK_0_H7_o(6) => SHA256_BLOCK_0_H7_o(6), 
        SHA256_BLOCK_0_H7_o(5) => SHA256_BLOCK_0_H7_o(5), 
        SHA256_BLOCK_0_H7_o(4) => SHA256_BLOCK_0_H7_o(4), 
        SHA256_BLOCK_0_H7_o(3) => SHA256_BLOCK_0_H7_o(3), 
        SHA256_BLOCK_0_H7_o(2) => SHA256_BLOCK_0_H7_o(2), 
        SHA256_BLOCK_0_H7_o(1) => SHA256_BLOCK_0_H7_o(1), 
        SHA256_BLOCK_0_H7_o(0) => SHA256_BLOCK_0_H7_o(0), state_0
         => \state[1]\, state_2 => \state[3]\, state_3 => 
        \state[4]\, sha256_controller_0_di_o_3 => 
        \sha256_controller_0_di_o[16]\, 
        sha256_controller_0_di_o_5 => 
        \sha256_controller_0_di_o[18]\, 
        sha256_controller_0_di_o_0 => 
        \sha256_controller_0_di_o[13]\, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, 
        SHA256_Module_0_di_req_o => \SHA256_Module_0_di_req_o\, 
        SHA256_BLOCK_0_do_valid_o => \SHA256_BLOCK_0_do_valid_o\, 
        SHA256_Module_0_waiting_data => 
        \SHA256_Module_0_waiting_data\, 
        SHA256_Module_0_data_available_lastbank_8 => 
        \SHA256_Module_0_data_available_lastbank_8\, N_484 => 
        N_484, bytes_sel => bytes_sel, SHA256_Module_0_error_o
         => SHA256_Module_0_error_o, SHA256_BLOCK_0_start_o => 
        \SHA256_BLOCK_0_start_o\, N_1702 => N_1702, N_1710 => 
        N_1710, ren_pos => ren_pos, N_1690 => N_1690, N_1691 => 
        N_1691, N_1693 => N_1693, N_1692 => N_1692, N_1718 => 
        N_1718, N_1694 => N_1694, N_1698 => N_1698, N_1701 => 
        N_1701, N_1696 => N_1696, N_1697 => N_1697, N_1695 => 
        N_1695, N_1699 => N_1699, N_1707 => N_1707, N_1708 => 
        N_1708, N_1709 => N_1709, N_1706 => N_1706, N_1704 => 
        N_1704, N_1688 => N_1688, N_1687 => N_1687, N_1689 => 
        N_1689, N_1713 => N_1713, N_1716 => N_1716, N_1712 => 
        N_1712, N_1717 => N_1717, N_1715 => N_1715, N_1711 => 
        N_1711, N_1714 => N_1714);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    limiter_1cycle_first : limiter_1cycle
      port map(prev_sig => prev_sig, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, first_block => 
        first_block);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    limiter_1cycle_ready : limiter_1cycle_0
      port map(prev_sig => prev_sig_0, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, data_out_ready => 
        \data_out_ready\);
    
    reg_17x32_0 : reg_17x32
      port map(reg_17x32_0_last_word(3) => 
        \reg_17x32_0_last_word[3]\, reg_17x32_0_last_word(2) => 
        \reg_17x32_0_last_word[2]\, reg_17x32_0_last_word(1) => 
        \reg_17x32_0_last_word[1]\, reg_17x32_0_last_word(0) => 
        \reg_17x32_0_last_word[0]\, reg_17x32_0_valid_bytes_0(1)
         => \reg_17x32_0_valid_bytes_0[1]\, 
        reg_17x32_0_valid_bytes_0(0) => 
        \reg_17x32_0_valid_bytes_0[0]\, 
        sha256_controller_0_read_addr_0(3) => 
        \sha256_controller_0_read_addr_0[3]\, 
        sha256_controller_0_read_addr_0(2) => 
        \sha256_controller_0_read_addr_0[2]\, 
        sha256_controller_0_read_addr_0(1) => 
        \sha256_controller_0_read_addr_0[1]\, 
        sha256_controller_0_read_addr_0(0) => 
        \sha256_controller_0_read_addr_0[0]\, waddr_in_net_0(4)
         => waddr_in_net_0(4), waddr_in_net_0(3) => 
        waddr_in_net_0(3), waddr_in_net_0(2) => waddr_in_net_0(2), 
        waddr_in_net_0(1) => waddr_in_net_0(1), waddr_in_net_0(0)
         => waddr_in_net_0(0), data_out_ready => \data_out_ready\, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, 
        CertificationSystem_sb_0_GPIO_9_M2F => 
        CertificationSystem_sb_0_GPIO_9_M2F, 
        SHA256_Module_0_data_available => 
        SHA256_Module_0_data_available, ren_pos => ren_pos, 
        N_111_i_0 => N_111_i_0, N_109_i_0 => N_109_i_0, N_168_i_0
         => N_168_i_0, N_107_i_0 => N_107_i_0, N_99_i_0 => 
        N_99_i_0, N_97_i_0 => N_97_i_0, 
        SHA256_Module_0_data_available_lastbank_8 => 
        \SHA256_Module_0_data_available_lastbank_8\, N_67_i_0 => 
        N_67_i_0, first_block => first_block, N_65_i_0 => 
        N_65_i_0, CertificationSystem_sb_0_GPIO_9_M2F_i_0 => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, N_105_i_0 => 
        N_105_i_0, N_103_i_0 => N_103_i_0, N_158_i_0 => N_158_i_0, 
        N_156_i_0 => N_156_i_0, N_101_i_0 => N_101_i_0, N_152_i_0
         => N_152_i_0, N_95_i_0 => N_95_i_0, N_93_i_0 => N_93_i_0, 
        N_91_i_0 => N_91_i_0, N_140_i_0 => N_140_i_0, N_89_i_0
         => N_89_i_0, N_87_i_0 => N_87_i_0, N_133_i_0 => 
        N_133_i_0, N_85_i_0 => N_85_i_0, N_83_i_0 => N_83_i_0, 
        N_77_i_0 => N_77_i_0, N_75_i_0 => N_75_i_0, N_73_i_0 => 
        N_73_i_0, N_71_i_0 => N_71_i_0, N_69_i_0 => N_69_i_0, 
        N_116_i_0 => N_116_i_0, N_114_i_0 => N_114_i_0, N_112_i_0
         => N_112_i_0, N_110_i_0 => N_110_i_0, N_1687 => N_1687, 
        N_1717 => N_1717, N_1690 => N_1690, N_1689 => N_1689, 
        N_1688 => N_1688, N_1715 => N_1715, N_1713 => N_1713, 
        N_1710 => N_1710, N_1701 => N_1701, N_1714 => N_1714, 
        N_1712 => N_1712, N_1716 => N_1716, N_1700 => N_1700, 
        N_1698 => N_1698, N_1697 => N_1697, N_1692 => N_1692, 
        N_1691 => N_1691, N_1704 => N_1704, N_1694 => N_1694, 
        N_1709 => N_1709, N_1708 => N_1708, N_1707 => N_1707, 
        N_1718 => N_1718, N_1703 => N_1703, N_1696 => N_1696, 
        N_1699 => N_1699, N_1705 => N_1705, N_1695 => N_1695, 
        N_1693 => N_1693, N_1706 => N_1706, N_1702 => N_1702, 
        N_1711 => N_1711, CertificationSystem_sb_0_GPIO_1_M2F => 
        CertificationSystem_sb_0_GPIO_1_M2F, 
        AHB_slave_dummy_0_write_en => AHB_slave_dummy_0_write_en);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_1 is

    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o                  : in    std_logic_vector(31 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          wen_or_i_3_i_0                       : in    std_logic;
          data_out_ready                       : in    std_logic
        );

end reg_1x32_1;

architecture DEF_ARCH of reg_1x32_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(12), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(3), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(23), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(10), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(26), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(31), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(15), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(19), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(14), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(5), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(22), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(20), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(17), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(2), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(18), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(4), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(25), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(30), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(29), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(11), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(24), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(9), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(13), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(27), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(16), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(8), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(28), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(7), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(21), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H1_o(6), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity mux_9_1 is

    port( line_7                      : in    std_logic_vector(0 to 0);
          result_addr_net_0           : in    std_logic_vector(3 downto 0);
          line_31                     : in    std_logic;
          line_28                     : in    std_logic;
          line_5_d0                   : in    std_logic;
          line_23                     : in    std_logic;
          line_8                      : in    std_logic;
          line_13                     : in    std_logic;
          line_0_d0                   : in    std_logic;
          line_12                     : in    std_logic;
          line_0_31                   : in    std_logic;
          line_0_28                   : in    std_logic;
          line_0_5                    : in    std_logic;
          line_0_23                   : in    std_logic;
          line_0_8                    : in    std_logic;
          line_0_13                   : in    std_logic;
          line_0_0                    : in    std_logic;
          line_0_12                   : in    std_logic;
          line_1_31                   : in    std_logic;
          line_1_28                   : in    std_logic;
          line_1_5                    : in    std_logic;
          line_1_23                   : in    std_logic;
          line_1_8                    : in    std_logic;
          line_1_13                   : in    std_logic;
          line_1_0                    : in    std_logic;
          line_1_12                   : in    std_logic;
          line_2_31                   : in    std_logic;
          line_2_28                   : in    std_logic;
          line_2_5                    : in    std_logic;
          line_2_23                   : in    std_logic;
          line_2_8                    : in    std_logic;
          line_2_13                   : in    std_logic;
          line_2_0                    : in    std_logic;
          line_2_12                   : in    std_logic;
          line_3_5                    : in    std_logic;
          line_3_13                   : in    std_logic;
          line_3_12                   : in    std_logic;
          line_3_0                    : in    std_logic;
          line_3_8                    : in    std_logic;
          line_3_23                   : in    std_logic;
          line_4_5                    : in    std_logic;
          line_4_13                   : in    std_logic;
          line_4_12                   : in    std_logic;
          line_4_0                    : in    std_logic;
          line_4_8                    : in    std_logic;
          line_4_23                   : in    std_logic;
          line_5_5                    : in    std_logic;
          line_5_13                   : in    std_logic;
          line_5_12                   : in    std_logic;
          line_5_0                    : in    std_logic;
          line_5_8                    : in    std_logic;
          line_5_23                   : in    std_logic;
          line_6_5                    : in    std_logic;
          line_6_13                   : in    std_logic;
          line_6_12                   : in    std_logic;
          line_6_0                    : in    std_logic;
          line_6_8                    : in    std_logic;
          line_6_23                   : in    std_logic;
          SHA256_Module_0_data_out_5  : out   std_logic;
          SHA256_Module_0_data_out_13 : out   std_logic;
          SHA256_Module_0_data_out_12 : out   std_logic;
          SHA256_Module_0_data_out_23 : out   std_logic;
          SHA256_Module_0_data_out_8  : out   std_logic;
          SHA256_Module_0_data_out_0  : out   std_logic;
          N_507                       : out   std_logic;
          N_508                       : out   std_logic;
          ren_pos                     : in    std_logic
        );

end mux_9_1;

architecture DEF_ARCH of mux_9_1 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \data_out_5_i_m3_i_m3_1_1[31]_net_1\, 
        \data_out_6_i_m2_i_m3_1_1[28]_net_1\, 
        \data_out_5_bm[23]_net_1\, \data_out_5_am[23]_net_1\, 
        N_551, \data_out_4_bm[8]_net_1\, \data_out_4_am[8]_net_1\, 
        N_504, \data_out_5_bm[0]_net_1\, \data_out_5_am[0]_net_1\, 
        N_528, \data_out_4_bm[12]_net_1\, 
        \data_out_4_am[12]_net_1\, N_508_0, 
        \data_out_5_bm[12]_net_1\, \data_out_5_am[12]_net_1\, 
        N_540, \data_out_4_bm[0]_net_1\, \data_out_4_am[0]_net_1\, 
        N_496, \data_out_5_bm[13]_net_1\, 
        \data_out_5_am[13]_net_1\, N_541, 
        \data_out_4_bm[13]_net_1\, \data_out_4_am[13]_net_1\, 
        N_509, \data_out_5_bm[8]_net_1\, \data_out_5_am[8]_net_1\, 
        N_536, \data_out_5_bm[5]_net_1\, \data_out_5_am[5]_net_1\, 
        N_533, \data_out_4_bm[23]_net_1\, 
        \data_out_4_am[23]_net_1\, N_519, 
        \data_out_4_bm[5]_net_1\, \data_out_4_am[5]_net_1\, N_501, 
        N_562, GND_net_1, VCC_net_1 : std_logic;

begin 


    \data_out_5_bm[13]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_13, B => line_4_13, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[13]_net_1\);
    
    \data_out_5_am[0]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_0, B => line_6_0, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[0]_net_1\);
    
    \data_out_4_ns[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[0]_net_1\, C => \data_out_4_am[0]_net_1\, 
        Y => N_496);
    
    \data_out_5_ns[23]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_5_bm[23]_net_1\, C => \data_out_5_am[23]_net_1\, 
        Y => N_551);
    
    \data_out_5_bm[23]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_23, B => line_4_23, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[23]_net_1\);
    
    \data_out_4_ns[23]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[23]_net_1\, C => \data_out_4_am[23]_net_1\, 
        Y => N_519);
    
    \data_out[8]\ : CFG4
      generic map(INIT => x"DC10")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(0), C => N_536, D => N_504, Y => 
        SHA256_Module_0_data_out_8);
    
    \data_out_6_i_m2_i_m3[28]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => result_addr_net_0(1), B => 
        \data_out_6_i_m2_i_m3_1_1[28]_net_1\, C => line_28, D => 
        line_0_28, Y => N_508);
    
    \data_out_5_bm[12]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_12, B => line_0_12, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[12]_net_1\);
    
    \data_out_5_am[12]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_12, B => line_2_12, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[12]_net_1\);
    
    \data_out_5_ns[5]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_5_bm[5]_net_1\, C => \data_out_5_am[5]_net_1\, 
        Y => N_533);
    
    \data_out_5_am[5]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_5, B => line_6_5, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[5]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \data_out_4_am[13]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_13, B => line_2_13, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[13]_net_1\);
    
    \data_out_4_am[0]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_0, B => line_2_0, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[0]_net_1\);
    
    \data_out_4_am[23]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_23, B => line_2_23, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[23]_net_1\);
    
    \data_out[13]\ : CFG4
      generic map(INIT => x"DC10")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(0), C => N_541, D => N_509, Y => 
        SHA256_Module_0_data_out_13);
    
    \data_out_5_ns[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_5_bm[0]_net_1\, C => \data_out_5_am[0]_net_1\, 
        Y => N_528);
    
    \data_out_5_am[8]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_8, B => line_2_8, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[8]_net_1\);
    
    \data_out_4_bm[13]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_13, B => line_0_13, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[13]_net_1\);
    
    \data_out_4_am[5]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_1_5, B => line_2_5, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[5]_net_1\);
    
    \data_out_4_bm[12]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_12, B => line_4_12, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[12]_net_1\);
    
    \data_out_4_bm[23]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_23, B => line_0_23, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[23]_net_1\);
    
    \data_out_6_i_m2_i_m3_1_1[28]\ : CFG4
      generic map(INIT => x"350F")

      port map(A => line_1_28, B => line_2_28, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \data_out_6_i_m2_i_m3_1_1[28]_net_1\);
    
    \data_out[12]\ : CFG4
      generic map(INIT => x"DC10")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(0), C => N_540, D => N_508_0, Y => 
        SHA256_Module_0_data_out_12);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \data_out_5_ns[13]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_5_bm[13]_net_1\, C => \data_out_5_am[13]_net_1\, 
        Y => N_541);
    
    \data_out_5_bm[0]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_0, B => line_4_0, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[0]_net_1\);
    
    \data_out_5_am[13]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_13, B => line_6_13, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[13]_net_1\);
    
    \data_out_4_ns[13]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[13]_net_1\, C => \data_out_4_am[13]_net_1\, 
        Y => N_509);
    
    \data_out_5_i_m3_i_m3[31]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => result_addr_net_0(1), B => 
        \data_out_5_i_m3_i_m3_1_1[31]_net_1\, C => line_31, D => 
        line_0_31, Y => N_507);
    
    \data_out_5_am[23]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_23, B => line_6_23, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_am[23]_net_1\);
    
    \data_out[5]\ : CFG4
      generic map(INIT => x"DC10")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(0), C => N_533, D => N_501, Y => 
        SHA256_Module_0_data_out_5);
    
    \data_out_4_ns[8]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[8]_net_1\, C => \data_out_4_am[8]_net_1\, 
        Y => N_504);
    
    \data_out_4_am[8]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_8, B => line_6_8, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[8]_net_1\);
    
    \data_out_5_bm[5]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_5, B => line_4_5, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[5]_net_1\);
    
    \data_out[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_562, B => result_addr_net_0(0), C => N_496, 
        Y => SHA256_Module_0_data_out_0);
    
    \data_out_4_bm[0]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_0_d0, B => line_0_0, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[0]_net_1\);
    
    \data_out[23]\ : CFG4
      generic map(INIT => x"DC10")

      port map(A => result_addr_net_0(3), B => 
        result_addr_net_0(0), C => N_551, D => N_519, Y => 
        SHA256_Module_0_data_out_23);
    
    \data_out_5_i_m3_i_m3_1_1[31]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_31, B => line_2_31, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \data_out_5_i_m3_i_m3_1_1[31]_net_1\);
    
    \data_out_4_am[12]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_12, B => line_6_12, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_am[12]_net_1\);
    
    \data_out_5_bm[8]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_8, B => line_0_8, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_5_bm[8]_net_1\);
    
    \data_out_4_bm[5]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_5_d0, B => line_0_5, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[5]_net_1\);
    
    \data_out_5_ns[8]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_5_bm[8]_net_1\, C => \data_out_5_am[8]_net_1\, 
        Y => N_536);
    
    \data_out_6[0]\ : CFG4
      generic map(INIT => x"D850")

      port map(A => result_addr_net_0(3), B => line_7(0), C => 
        N_528, D => ren_pos, Y => N_562);
    
    \data_out_4_ns[5]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[5]_net_1\, C => \data_out_4_am[5]_net_1\, 
        Y => N_501);
    
    \data_out_5_ns[12]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_5_bm[12]_net_1\, C => \data_out_5_am[12]_net_1\, 
        Y => N_540);
    
    \data_out_4_bm[8]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => line_3_8, B => line_4_8, C => 
        result_addr_net_0(2), D => ren_pos, Y => 
        \data_out_4_bm[8]_net_1\);
    
    \data_out_4_ns[12]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => result_addr_net_0(1), B => 
        \data_out_4_bm[12]_net_1\, C => \data_out_4_am[12]_net_1\, 
        Y => N_508_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32 is

    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H0_o                  : in    std_logic_vector(31 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          wen_or_i_3_i_0                       : out   std_logic;
          data_out_ready                       : in    std_logic;
          ren_pos                              : out   std_logic;
          AHB_slave_dummy_0_read_en            : in    std_logic;
          start_wen                            : in    std_logic
        );

end reg_1x32;

architecture DEF_ARCH of reg_1x32 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \wen_or_i_3_i_0\, GND_net_1, ren_pos_0
         : std_logic;

begin 

    wen_or_i_3_i_0 <= \wen_or_i_3_i_0\;

    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(12), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(3), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(23), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(10), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(26), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(31), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(15), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(19), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(14), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(5), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(22), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(20), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(17), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(2), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(18), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(18));
    
    \ren_pos\ : SLE
      port map(D => ren_pos_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => ren_pos);
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(4), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(25), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(30), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(29), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(11), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(24), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(9), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(13), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(27), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(16), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(16));
    
    wen_or_i_3_i : CFG2
      generic map(INIT => x"D")

      port map(A => data_out_ready, B => start_wen, Y => 
        \wen_or_i_3_i_0\);
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(8), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(28), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(7), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(7));
    
    ren_pos_r : CFG2
      generic map(INIT => x"8")

      port map(A => data_out_ready, B => 
        AHB_slave_dummy_0_read_en, Y => ren_pos_0);
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(21), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H0_o(6), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \wen_or_i_3_i_0\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_7 is

    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o                  : in    std_logic_vector(31 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          wen_or_i_3_i_0                       : in    std_logic;
          data_out_ready                       : in    std_logic
        );

end reg_1x32_7;

architecture DEF_ARCH of reg_1x32_7 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(12), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(3), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(23), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(10), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(26), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(31), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(15), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(19), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(14), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(5), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(22), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(20), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(17), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(2), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(18), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(4), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(25), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(30), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(29), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(11), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(24), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(9), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(13), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(27), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(16), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(8), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(28), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(7), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(21), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H7_o(6), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_6 is

    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o                  : in    std_logic_vector(31 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          wen_or_i_3_i_0                       : in    std_logic;
          data_out_ready                       : in    std_logic
        );

end reg_1x32_6;

architecture DEF_ARCH of reg_1x32_6 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(12), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(3), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(23), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(10), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(26), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(31), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(15), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(19), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(14), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(5), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(22), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(20), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(17), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(2), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(18), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(4), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(25), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(30), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(29), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(11), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(24), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(9), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(13), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(27), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(16), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(8), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(28), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(7), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(21), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H6_o(6), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_5 is

    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o                  : in    std_logic_vector(31 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          wen_or_i_3_i_0                       : in    std_logic;
          data_out_ready                       : in    std_logic
        );

end reg_1x32_5;

architecture DEF_ARCH of reg_1x32_5 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(12), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(3), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(23), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(10), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(26), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(31), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(15), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(19), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(14), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(5), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(22), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(20), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(17), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(2), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(18), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(4), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(25), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(30), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(29), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(11), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(24), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(9), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(13), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(27), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(16), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(8), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(28), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(7), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(21), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H5_o(6), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_2 is

    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o                  : in    std_logic_vector(31 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          wen_or_i_3_i_0                       : in    std_logic;
          data_out_ready                       : in    std_logic
        );

end reg_1x32_2;

architecture DEF_ARCH of reg_1x32_2 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(12), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(3), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(23), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(10), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(26), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(31), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(15), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(19), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(14), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(5), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(22), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(20), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(17), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(2), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(18), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(4), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(25), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(30), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(29), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(11), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(24), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(9), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(13), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(27), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(16), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(8), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(28), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(7), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(21), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H2_o(6), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_8 is

    port( line                                 : out   std_logic_vector(2 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          SHA256_Module_0_error_o              : in    std_logic;
          wen_or_i_3_i_0                       : in    std_logic;
          data_out_ready                       : in    std_logic;
          SHA256_Module_0_di_req_o             : in    std_logic;
          SHA256_Module_0_do_valid_o           : in    std_logic
        );

end reg_1x32_8;

architecture DEF_ARCH of reg_1x32_8 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_Module_0_error_o, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(2));
    
    \line[1]\ : SLE
      port map(D => SHA256_Module_0_di_req_o, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(1));
    
    \line[0]\ : SLE
      port map(D => SHA256_Module_0_do_valid_o, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(0));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_3 is

    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o                  : in    std_logic_vector(31 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          wen_or_i_3_i_0                       : in    std_logic;
          data_out_ready                       : in    std_logic
        );

end reg_1x32_3;

architecture DEF_ARCH of reg_1x32_3 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(12), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(3), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(23), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(10), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(26), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(31), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(15), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(19), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(14), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(5), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(22), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(20), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(17), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(2), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(18), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(4), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(25), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(30), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(29), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(11), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(24), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(9), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(13), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(27), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(16), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(8), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(28), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(7), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(21), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H3_o(6), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg_1x32_4 is

    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o                  : in    std_logic_vector(31 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          wen_or_i_3_i_0                       : in    std_logic;
          data_out_ready                       : in    std_logic
        );

end reg_1x32_4;

architecture DEF_ARCH of reg_1x32_4 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \line[12]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(12), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(12));
    
    \line[3]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(3), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(3));
    
    \line[23]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(23), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(23));
    
    \line[10]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(10), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(10));
    
    \line[26]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(26), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(26));
    
    \line[31]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(31), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(31));
    
    \line[15]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(15), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \line[19]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(19), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(19));
    
    \line[14]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(14), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(14));
    
    \line[5]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(5), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(5));
    
    \line[22]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(22), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(22));
    
    \line[20]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(20), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(20));
    
    \line[17]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(17), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(17));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \line[2]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(2), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(2));
    
    \line[18]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(18), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(18));
    
    \line[4]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(4), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(4));
    
    \line[25]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(25), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(25));
    
    \line[30]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(30), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(30));
    
    \line[29]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(29), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(29));
    
    \line[11]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(11), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(11));
    
    \line[24]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(24), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(24));
    
    \line[9]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(9), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(9));
    
    \line[1]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(1), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(1));
    
    \line[13]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(13), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(13));
    
    \line[27]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(27), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(27));
    
    \line[16]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(16), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(16));
    
    \line[8]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(8), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(8));
    
    \line[28]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(28), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(28));
    
    \line[0]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(0), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(0));
    
    \line[7]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(7), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(7));
    
    \line[21]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(21), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(21));
    
    \line[6]\ : SLE
      port map(D => SHA256_BLOCK_0_H4_o(6), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        wen_or_i_3_i_0, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => data_out_ready, SD => GND_net_1, LAT => GND_net_1, Q
         => line(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg9_1x32 is

    port( result_addr_net_0                    : in    std_logic_vector(3 downto 0);
          SHA256_BLOCK_0_H0_o                  : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o                  : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o                  : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o                  : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o                  : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o                  : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o                  : in    std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o                  : in    std_logic_vector(31 downto 0);
          SHA256_Module_0_data_out_5           : out   std_logic;
          SHA256_Module_0_data_out_13          : out   std_logic;
          SHA256_Module_0_data_out_12          : out   std_logic;
          SHA256_Module_0_data_out_23          : out   std_logic;
          SHA256_Module_0_data_out_8           : out   std_logic;
          SHA256_Module_0_data_out_0           : out   std_logic;
          line_1_d0                            : out   std_logic;
          line_2_d0                            : out   std_logic;
          line_3_d0                            : out   std_logic;
          line_4_d0                            : out   std_logic;
          line_6_d0                            : out   std_logic;
          line_7_d0                            : out   std_logic;
          line_9                               : out   std_logic;
          line_10                              : out   std_logic;
          line_11                              : out   std_logic;
          line_14                              : out   std_logic;
          line_15                              : out   std_logic;
          line_16                              : out   std_logic;
          line_17                              : out   std_logic;
          line_18                              : out   std_logic;
          line_19                              : out   std_logic;
          line_20                              : out   std_logic;
          line_21                              : out   std_logic;
          line_22                              : out   std_logic;
          line_24                              : out   std_logic;
          line_25                              : out   std_logic;
          line_26                              : out   std_logic;
          line_27                              : out   std_logic;
          line_29                              : out   std_logic;
          line_30                              : out   std_logic;
          line_0_1                             : out   std_logic;
          line_0_2                             : out   std_logic;
          line_0_3                             : out   std_logic;
          line_0_4                             : out   std_logic;
          line_0_6                             : out   std_logic;
          line_0_7                             : out   std_logic;
          line_0_9                             : out   std_logic;
          line_0_10                            : out   std_logic;
          line_0_11                            : out   std_logic;
          line_0_14                            : out   std_logic;
          line_0_15                            : out   std_logic;
          line_0_16                            : out   std_logic;
          line_0_17                            : out   std_logic;
          line_0_18                            : out   std_logic;
          line_0_19                            : out   std_logic;
          line_0_20                            : out   std_logic;
          line_0_21                            : out   std_logic;
          line_0_22                            : out   std_logic;
          line_0_24                            : out   std_logic;
          line_0_25                            : out   std_logic;
          line_0_26                            : out   std_logic;
          line_0_27                            : out   std_logic;
          line_0_29                            : out   std_logic;
          line_0_30                            : out   std_logic;
          line_1_1                             : out   std_logic;
          line_1_2                             : out   std_logic;
          line_1_3                             : out   std_logic;
          line_1_4                             : out   std_logic;
          line_1_6                             : out   std_logic;
          line_1_7                             : out   std_logic;
          line_1_9                             : out   std_logic;
          line_1_10                            : out   std_logic;
          line_1_11                            : out   std_logic;
          line_1_14                            : out   std_logic;
          line_1_15                            : out   std_logic;
          line_1_16                            : out   std_logic;
          line_1_17                            : out   std_logic;
          line_1_18                            : out   std_logic;
          line_1_19                            : out   std_logic;
          line_1_20                            : out   std_logic;
          line_1_21                            : out   std_logic;
          line_1_22                            : out   std_logic;
          line_1_24                            : out   std_logic;
          line_1_25                            : out   std_logic;
          line_1_26                            : out   std_logic;
          line_1_27                            : out   std_logic;
          line_1_29                            : out   std_logic;
          line_1_30                            : out   std_logic;
          line_2_1                             : out   std_logic;
          line_2_2                             : out   std_logic;
          line_2_3                             : out   std_logic;
          line_2_4                             : out   std_logic;
          line_2_6                             : out   std_logic;
          line_2_7                             : out   std_logic;
          line_2_9                             : out   std_logic;
          line_2_10                            : out   std_logic;
          line_2_11                            : out   std_logic;
          line_2_14                            : out   std_logic;
          line_2_15                            : out   std_logic;
          line_2_16                            : out   std_logic;
          line_2_17                            : out   std_logic;
          line_2_18                            : out   std_logic;
          line_2_19                            : out   std_logic;
          line_2_20                            : out   std_logic;
          line_2_21                            : out   std_logic;
          line_2_22                            : out   std_logic;
          line_2_24                            : out   std_logic;
          line_2_25                            : out   std_logic;
          line_2_26                            : out   std_logic;
          line_2_27                            : out   std_logic;
          line_2_29                            : out   std_logic;
          line_2_30                            : out   std_logic;
          line_3_28                            : out   std_logic;
          line_3_31                            : out   std_logic;
          line_3_1                             : out   std_logic;
          line_3_2                             : out   std_logic;
          line_3_3                             : out   std_logic;
          line_3_4                             : out   std_logic;
          line_3_6                             : out   std_logic;
          line_3_7                             : out   std_logic;
          line_3_9                             : out   std_logic;
          line_3_10                            : out   std_logic;
          line_3_11                            : out   std_logic;
          line_3_14                            : out   std_logic;
          line_3_15                            : out   std_logic;
          line_3_16                            : out   std_logic;
          line_3_17                            : out   std_logic;
          line_3_18                            : out   std_logic;
          line_3_19                            : out   std_logic;
          line_3_20                            : out   std_logic;
          line_3_21                            : out   std_logic;
          line_3_22                            : out   std_logic;
          line_3_24                            : out   std_logic;
          line_3_25                            : out   std_logic;
          line_3_26                            : out   std_logic;
          line_3_27                            : out   std_logic;
          line_3_29                            : out   std_logic;
          line_3_30                            : out   std_logic;
          line_4_28                            : out   std_logic;
          line_4_31                            : out   std_logic;
          line_4_1                             : out   std_logic;
          line_4_2                             : out   std_logic;
          line_4_3                             : out   std_logic;
          line_4_4                             : out   std_logic;
          line_4_6                             : out   std_logic;
          line_4_7                             : out   std_logic;
          line_4_9                             : out   std_logic;
          line_4_10                            : out   std_logic;
          line_4_11                            : out   std_logic;
          line_4_14                            : out   std_logic;
          line_4_15                            : out   std_logic;
          line_4_16                            : out   std_logic;
          line_4_17                            : out   std_logic;
          line_4_18                            : out   std_logic;
          line_4_19                            : out   std_logic;
          line_4_20                            : out   std_logic;
          line_4_21                            : out   std_logic;
          line_4_22                            : out   std_logic;
          line_4_24                            : out   std_logic;
          line_4_25                            : out   std_logic;
          line_4_26                            : out   std_logic;
          line_4_27                            : out   std_logic;
          line_4_29                            : out   std_logic;
          line_4_30                            : out   std_logic;
          line_5_28                            : out   std_logic;
          line_5_31                            : out   std_logic;
          line_5_1                             : out   std_logic;
          line_5_2                             : out   std_logic;
          line_5_3                             : out   std_logic;
          line_5_4                             : out   std_logic;
          line_5_6                             : out   std_logic;
          line_5_7                             : out   std_logic;
          line_5_9                             : out   std_logic;
          line_5_10                            : out   std_logic;
          line_5_11                            : out   std_logic;
          line_5_14                            : out   std_logic;
          line_5_15                            : out   std_logic;
          line_5_16                            : out   std_logic;
          line_5_17                            : out   std_logic;
          line_5_18                            : out   std_logic;
          line_5_19                            : out   std_logic;
          line_5_20                            : out   std_logic;
          line_5_21                            : out   std_logic;
          line_5_22                            : out   std_logic;
          line_5_24                            : out   std_logic;
          line_5_25                            : out   std_logic;
          line_5_26                            : out   std_logic;
          line_5_27                            : out   std_logic;
          line_5_29                            : out   std_logic;
          line_5_30                            : out   std_logic;
          line_6_1                             : out   std_logic;
          line_6_2                             : out   std_logic;
          line_6_3                             : out   std_logic;
          line_6_4                             : out   std_logic;
          line_6_6                             : out   std_logic;
          line_6_7                             : out   std_logic;
          line_6_9                             : out   std_logic;
          line_6_10                            : out   std_logic;
          line_6_11                            : out   std_logic;
          line_6_14                            : out   std_logic;
          line_6_15                            : out   std_logic;
          line_6_16                            : out   std_logic;
          line_6_17                            : out   std_logic;
          line_6_18                            : out   std_logic;
          line_6_19                            : out   std_logic;
          line_6_20                            : out   std_logic;
          line_6_21                            : out   std_logic;
          line_6_22                            : out   std_logic;
          line_6_24                            : out   std_logic;
          line_6_25                            : out   std_logic;
          line_6_26                            : out   std_logic;
          line_6_27                            : out   std_logic;
          line_6_28                            : out   std_logic;
          line_6_29                            : out   std_logic;
          line_6_30                            : out   std_logic;
          line_6_31                            : out   std_logic;
          line_7_1                             : out   std_logic;
          line_7_2                             : out   std_logic;
          N_507                                : out   std_logic;
          N_508                                : out   std_logic;
          ren_pos                              : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          data_out_ready                       : in    std_logic;
          AHB_slave_dummy_0_read_en            : in    std_logic;
          start_wen                            : in    std_logic;
          SHA256_Module_0_error_o              : in    std_logic;
          SHA256_Module_0_di_req_o             : in    std_logic;
          SHA256_Module_0_do_valid_o           : in    std_logic
        );

end reg9_1x32;

architecture DEF_ARCH of reg9_1x32 is 

  component reg_1x32_1
    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          wen_or_i_3_i_0                       : in    std_logic := 'U';
          data_out_ready                       : in    std_logic := 'U'
        );
  end component;

  component mux_9_1
    port( line_7                      : in    std_logic_vector(0 to 0) := (others => 'U');
          result_addr_net_0           : in    std_logic_vector(3 downto 0) := (others => 'U');
          line_31                     : in    std_logic := 'U';
          line_28                     : in    std_logic := 'U';
          line_5_d0                   : in    std_logic := 'U';
          line_23                     : in    std_logic := 'U';
          line_8                      : in    std_logic := 'U';
          line_13                     : in    std_logic := 'U';
          line_0_d0                   : in    std_logic := 'U';
          line_12                     : in    std_logic := 'U';
          line_0_31                   : in    std_logic := 'U';
          line_0_28                   : in    std_logic := 'U';
          line_0_5                    : in    std_logic := 'U';
          line_0_23                   : in    std_logic := 'U';
          line_0_8                    : in    std_logic := 'U';
          line_0_13                   : in    std_logic := 'U';
          line_0_0                    : in    std_logic := 'U';
          line_0_12                   : in    std_logic := 'U';
          line_1_31                   : in    std_logic := 'U';
          line_1_28                   : in    std_logic := 'U';
          line_1_5                    : in    std_logic := 'U';
          line_1_23                   : in    std_logic := 'U';
          line_1_8                    : in    std_logic := 'U';
          line_1_13                   : in    std_logic := 'U';
          line_1_0                    : in    std_logic := 'U';
          line_1_12                   : in    std_logic := 'U';
          line_2_31                   : in    std_logic := 'U';
          line_2_28                   : in    std_logic := 'U';
          line_2_5                    : in    std_logic := 'U';
          line_2_23                   : in    std_logic := 'U';
          line_2_8                    : in    std_logic := 'U';
          line_2_13                   : in    std_logic := 'U';
          line_2_0                    : in    std_logic := 'U';
          line_2_12                   : in    std_logic := 'U';
          line_3_5                    : in    std_logic := 'U';
          line_3_13                   : in    std_logic := 'U';
          line_3_12                   : in    std_logic := 'U';
          line_3_0                    : in    std_logic := 'U';
          line_3_8                    : in    std_logic := 'U';
          line_3_23                   : in    std_logic := 'U';
          line_4_5                    : in    std_logic := 'U';
          line_4_13                   : in    std_logic := 'U';
          line_4_12                   : in    std_logic := 'U';
          line_4_0                    : in    std_logic := 'U';
          line_4_8                    : in    std_logic := 'U';
          line_4_23                   : in    std_logic := 'U';
          line_5_5                    : in    std_logic := 'U';
          line_5_13                   : in    std_logic := 'U';
          line_5_12                   : in    std_logic := 'U';
          line_5_0                    : in    std_logic := 'U';
          line_5_8                    : in    std_logic := 'U';
          line_5_23                   : in    std_logic := 'U';
          line_6_5                    : in    std_logic := 'U';
          line_6_13                   : in    std_logic := 'U';
          line_6_12                   : in    std_logic := 'U';
          line_6_0                    : in    std_logic := 'U';
          line_6_8                    : in    std_logic := 'U';
          line_6_23                   : in    std_logic := 'U';
          SHA256_Module_0_data_out_5  : out   std_logic;
          SHA256_Module_0_data_out_13 : out   std_logic;
          SHA256_Module_0_data_out_12 : out   std_logic;
          SHA256_Module_0_data_out_23 : out   std_logic;
          SHA256_Module_0_data_out_8  : out   std_logic;
          SHA256_Module_0_data_out_0  : out   std_logic;
          N_507                       : out   std_logic;
          N_508                       : out   std_logic;
          ren_pos                     : in    std_logic := 'U'
        );
  end component;

  component reg_1x32
    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H0_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          wen_or_i_3_i_0                       : out   std_logic;
          data_out_ready                       : in    std_logic := 'U';
          ren_pos                              : out   std_logic;
          AHB_slave_dummy_0_read_en            : in    std_logic := 'U';
          start_wen                            : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_7
    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          wen_or_i_3_i_0                       : in    std_logic := 'U';
          data_out_ready                       : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_6
    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          wen_or_i_3_i_0                       : in    std_logic := 'U';
          data_out_ready                       : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component reg_1x32_5
    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          wen_or_i_3_i_0                       : in    std_logic := 'U';
          data_out_ready                       : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_2
    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          wen_or_i_3_i_0                       : in    std_logic := 'U';
          data_out_ready                       : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_8
    port( line                                 : out   std_logic_vector(2 downto 0);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          SHA256_Module_0_error_o              : in    std_logic := 'U';
          wen_or_i_3_i_0                       : in    std_logic := 'U';
          data_out_ready                       : in    std_logic := 'U';
          SHA256_Module_0_di_req_o             : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o           : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_3
    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          wen_or_i_3_i_0                       : in    std_logic := 'U';
          data_out_ready                       : in    std_logic := 'U'
        );
  end component;

  component reg_1x32_4
    port( line                                 : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          wen_or_i_3_i_0                       : in    std_logic := 'U';
          data_out_ready                       : in    std_logic := 'U'
        );
  end component;

    signal \line[31]\, \line[28]\, \line[5]\, \line[23]\, 
        \line[8]\, \line[13]\, \line[0]\, \line[12]\, 
        \line_0[31]\, \line_0[28]\, \line_0[5]\, \line_0[23]\, 
        \line_0[8]\, \line_0[13]\, \line_0[0]\, \line_0[12]\, 
        \line_1[31]\, \line_1[28]\, \line_1[5]\, \line_1[23]\, 
        \line_1[8]\, \line_1[13]\, \line_1[0]\, \line_1[12]\, 
        \line_2[31]\, \line_2[28]\, \line_2[5]\, \line_2[23]\, 
        \line_2[8]\, \line_2[13]\, \line_2[0]\, \line_2[12]\, 
        \line_3[5]\, \line_3[13]\, \line_3[12]\, \line_3[0]\, 
        \line_3[8]\, \line_3[23]\, \line_4[5]\, \line_4[13]\, 
        \line_4[12]\, \line_4[0]\, \line_4[8]\, \line_4[23]\, 
        \line_5[5]\, \line_5[13]\, \line_5[12]\, \line_5[0]\, 
        \line_5[8]\, \line_5[23]\, \line_6[5]\, \line_6[13]\, 
        \line_6[12]\, \line_6[0]\, \line_6[8]\, \line_6[23]\, 
        \line_7[0]\, \ren_pos\, wen_or_i_3_i_0, GND_net_1, 
        VCC_net_1 : std_logic;

    for all : reg_1x32_1
	Use entity work.reg_1x32_1(DEF_ARCH);
    for all : mux_9_1
	Use entity work.mux_9_1(DEF_ARCH);
    for all : reg_1x32
	Use entity work.reg_1x32(DEF_ARCH);
    for all : reg_1x32_7
	Use entity work.reg_1x32_7(DEF_ARCH);
    for all : reg_1x32_6
	Use entity work.reg_1x32_6(DEF_ARCH);
    for all : reg_1x32_5
	Use entity work.reg_1x32_5(DEF_ARCH);
    for all : reg_1x32_2
	Use entity work.reg_1x32_2(DEF_ARCH);
    for all : reg_1x32_8
	Use entity work.reg_1x32_8(DEF_ARCH);
    for all : reg_1x32_3
	Use entity work.reg_1x32_3(DEF_ARCH);
    for all : reg_1x32_4
	Use entity work.reg_1x32_4(DEF_ARCH);
begin 

    ren_pos <= \ren_pos\;

    \reg_1x32_1\ : reg_1x32_1
      port map(line(31) => line_3_31, line(30) => line_0_30, 
        line(29) => line_0_29, line(28) => line_3_28, line(27)
         => line_0_27, line(26) => line_0_26, line(25) => 
        line_0_25, line(24) => line_0_24, line(23) => 
        \line_1[23]\, line(22) => line_0_22, line(21) => 
        line_0_21, line(20) => line_0_20, line(19) => line_0_19, 
        line(18) => line_0_18, line(17) => line_0_17, line(16)
         => line_0_16, line(15) => line_0_15, line(14) => 
        line_0_14, line(13) => \line_1[13]\, line(12) => 
        \line_5[12]\, line(11) => line_0_11, line(10) => 
        line_0_10, line(9) => line_0_9, line(8) => \line_5[8]\, 
        line(7) => line_0_7, line(6) => line_0_6, line(5) => 
        \line_1[5]\, line(4) => line_0_4, line(3) => line_0_3, 
        line(2) => line_0_2, line(1) => line_0_1, line(0) => 
        \line_1[0]\, SHA256_BLOCK_0_H1_o(31) => 
        SHA256_BLOCK_0_H1_o(31), SHA256_BLOCK_0_H1_o(30) => 
        SHA256_BLOCK_0_H1_o(30), SHA256_BLOCK_0_H1_o(29) => 
        SHA256_BLOCK_0_H1_o(29), SHA256_BLOCK_0_H1_o(28) => 
        SHA256_BLOCK_0_H1_o(28), SHA256_BLOCK_0_H1_o(27) => 
        SHA256_BLOCK_0_H1_o(27), SHA256_BLOCK_0_H1_o(26) => 
        SHA256_BLOCK_0_H1_o(26), SHA256_BLOCK_0_H1_o(25) => 
        SHA256_BLOCK_0_H1_o(25), SHA256_BLOCK_0_H1_o(24) => 
        SHA256_BLOCK_0_H1_o(24), SHA256_BLOCK_0_H1_o(23) => 
        SHA256_BLOCK_0_H1_o(23), SHA256_BLOCK_0_H1_o(22) => 
        SHA256_BLOCK_0_H1_o(22), SHA256_BLOCK_0_H1_o(21) => 
        SHA256_BLOCK_0_H1_o(21), SHA256_BLOCK_0_H1_o(20) => 
        SHA256_BLOCK_0_H1_o(20), SHA256_BLOCK_0_H1_o(19) => 
        SHA256_BLOCK_0_H1_o(19), SHA256_BLOCK_0_H1_o(18) => 
        SHA256_BLOCK_0_H1_o(18), SHA256_BLOCK_0_H1_o(17) => 
        SHA256_BLOCK_0_H1_o(17), SHA256_BLOCK_0_H1_o(16) => 
        SHA256_BLOCK_0_H1_o(16), SHA256_BLOCK_0_H1_o(15) => 
        SHA256_BLOCK_0_H1_o(15), SHA256_BLOCK_0_H1_o(14) => 
        SHA256_BLOCK_0_H1_o(14), SHA256_BLOCK_0_H1_o(13) => 
        SHA256_BLOCK_0_H1_o(13), SHA256_BLOCK_0_H1_o(12) => 
        SHA256_BLOCK_0_H1_o(12), SHA256_BLOCK_0_H1_o(11) => 
        SHA256_BLOCK_0_H1_o(11), SHA256_BLOCK_0_H1_o(10) => 
        SHA256_BLOCK_0_H1_o(10), SHA256_BLOCK_0_H1_o(9) => 
        SHA256_BLOCK_0_H1_o(9), SHA256_BLOCK_0_H1_o(8) => 
        SHA256_BLOCK_0_H1_o(8), SHA256_BLOCK_0_H1_o(7) => 
        SHA256_BLOCK_0_H1_o(7), SHA256_BLOCK_0_H1_o(6) => 
        SHA256_BLOCK_0_H1_o(6), SHA256_BLOCK_0_H1_o(5) => 
        SHA256_BLOCK_0_H1_o(5), SHA256_BLOCK_0_H1_o(4) => 
        SHA256_BLOCK_0_H1_o(4), SHA256_BLOCK_0_H1_o(3) => 
        SHA256_BLOCK_0_H1_o(3), SHA256_BLOCK_0_H1_o(2) => 
        SHA256_BLOCK_0_H1_o(2), SHA256_BLOCK_0_H1_o(1) => 
        SHA256_BLOCK_0_H1_o(1), SHA256_BLOCK_0_H1_o(0) => 
        SHA256_BLOCK_0_H1_o(0), 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, wen_or_i_3_i_0 => 
        wen_or_i_3_i_0, data_out_ready => data_out_ready);
    
    mux_9_1_0 : mux_9_1
      port map(line_7(0) => \line_7[0]\, result_addr_net_0(3) => 
        result_addr_net_0(3), result_addr_net_0(2) => 
        result_addr_net_0(2), result_addr_net_0(1) => 
        result_addr_net_0(1), result_addr_net_0(0) => 
        result_addr_net_0(0), line_31 => \line[31]\, line_28 => 
        \line[28]\, line_5_d0 => \line[5]\, line_23 => \line[23]\, 
        line_8 => \line[8]\, line_13 => \line[13]\, line_0_d0 => 
        \line[0]\, line_12 => \line[12]\, line_0_31 => 
        \line_0[31]\, line_0_28 => \line_0[28]\, line_0_5 => 
        \line_0[5]\, line_0_23 => \line_0[23]\, line_0_8 => 
        \line_0[8]\, line_0_13 => \line_0[13]\, line_0_0 => 
        \line_0[0]\, line_0_12 => \line_0[12]\, line_1_31 => 
        \line_1[31]\, line_1_28 => \line_1[28]\, line_1_5 => 
        \line_1[5]\, line_1_23 => \line_1[23]\, line_1_8 => 
        \line_1[8]\, line_1_13 => \line_1[13]\, line_1_0 => 
        \line_1[0]\, line_1_12 => \line_1[12]\, line_2_31 => 
        \line_2[31]\, line_2_28 => \line_2[28]\, line_2_5 => 
        \line_2[5]\, line_2_23 => \line_2[23]\, line_2_8 => 
        \line_2[8]\, line_2_13 => \line_2[13]\, line_2_0 => 
        \line_2[0]\, line_2_12 => \line_2[12]\, line_3_5 => 
        \line_3[5]\, line_3_13 => \line_3[13]\, line_3_12 => 
        \line_3[12]\, line_3_0 => \line_3[0]\, line_3_8 => 
        \line_3[8]\, line_3_23 => \line_3[23]\, line_4_5 => 
        \line_4[5]\, line_4_13 => \line_4[13]\, line_4_12 => 
        \line_4[12]\, line_4_0 => \line_4[0]\, line_4_8 => 
        \line_4[8]\, line_4_23 => \line_4[23]\, line_5_5 => 
        \line_5[5]\, line_5_13 => \line_5[13]\, line_5_12 => 
        \line_5[12]\, line_5_0 => \line_5[0]\, line_5_8 => 
        \line_5[8]\, line_5_23 => \line_5[23]\, line_6_5 => 
        \line_6[5]\, line_6_13 => \line_6[13]\, line_6_12 => 
        \line_6[12]\, line_6_0 => \line_6[0]\, line_6_8 => 
        \line_6[8]\, line_6_23 => \line_6[23]\, 
        SHA256_Module_0_data_out_5 => SHA256_Module_0_data_out_5, 
        SHA256_Module_0_data_out_13 => 
        SHA256_Module_0_data_out_13, SHA256_Module_0_data_out_12
         => SHA256_Module_0_data_out_12, 
        SHA256_Module_0_data_out_23 => 
        SHA256_Module_0_data_out_23, SHA256_Module_0_data_out_8
         => SHA256_Module_0_data_out_8, 
        SHA256_Module_0_data_out_0 => SHA256_Module_0_data_out_0, 
        N_507 => N_507, N_508 => N_508, ren_pos => \ren_pos\);
    
    reg_1x32_0 : reg_1x32
      port map(line(31) => \line_1[31]\, line(30) => line_30, 
        line(29) => line_29, line(28) => \line_0[28]\, line(27)
         => line_27, line(26) => line_26, line(25) => line_25, 
        line(24) => line_24, line(23) => \line_5[23]\, line(22)
         => line_22, line(21) => line_21, line(20) => line_20, 
        line(19) => line_19, line(18) => line_18, line(17) => 
        line_17, line(16) => line_16, line(15) => line_15, 
        line(14) => line_14, line(13) => \line_5[13]\, line(12)
         => \line_1[12]\, line(11) => line_11, line(10) => 
        line_10, line(9) => line_9, line(8) => \line_1[8]\, 
        line(7) => line_7_d0, line(6) => line_6_d0, line(5) => 
        \line_5[5]\, line(4) => line_4_d0, line(3) => line_3_d0, 
        line(2) => line_2_d0, line(1) => line_1_d0, line(0) => 
        \line_5[0]\, SHA256_BLOCK_0_H0_o(31) => 
        SHA256_BLOCK_0_H0_o(31), SHA256_BLOCK_0_H0_o(30) => 
        SHA256_BLOCK_0_H0_o(30), SHA256_BLOCK_0_H0_o(29) => 
        SHA256_BLOCK_0_H0_o(29), SHA256_BLOCK_0_H0_o(28) => 
        SHA256_BLOCK_0_H0_o(28), SHA256_BLOCK_0_H0_o(27) => 
        SHA256_BLOCK_0_H0_o(27), SHA256_BLOCK_0_H0_o(26) => 
        SHA256_BLOCK_0_H0_o(26), SHA256_BLOCK_0_H0_o(25) => 
        SHA256_BLOCK_0_H0_o(25), SHA256_BLOCK_0_H0_o(24) => 
        SHA256_BLOCK_0_H0_o(24), SHA256_BLOCK_0_H0_o(23) => 
        SHA256_BLOCK_0_H0_o(23), SHA256_BLOCK_0_H0_o(22) => 
        SHA256_BLOCK_0_H0_o(22), SHA256_BLOCK_0_H0_o(21) => 
        SHA256_BLOCK_0_H0_o(21), SHA256_BLOCK_0_H0_o(20) => 
        SHA256_BLOCK_0_H0_o(20), SHA256_BLOCK_0_H0_o(19) => 
        SHA256_BLOCK_0_H0_o(19), SHA256_BLOCK_0_H0_o(18) => 
        SHA256_BLOCK_0_H0_o(18), SHA256_BLOCK_0_H0_o(17) => 
        SHA256_BLOCK_0_H0_o(17), SHA256_BLOCK_0_H0_o(16) => 
        SHA256_BLOCK_0_H0_o(16), SHA256_BLOCK_0_H0_o(15) => 
        SHA256_BLOCK_0_H0_o(15), SHA256_BLOCK_0_H0_o(14) => 
        SHA256_BLOCK_0_H0_o(14), SHA256_BLOCK_0_H0_o(13) => 
        SHA256_BLOCK_0_H0_o(13), SHA256_BLOCK_0_H0_o(12) => 
        SHA256_BLOCK_0_H0_o(12), SHA256_BLOCK_0_H0_o(11) => 
        SHA256_BLOCK_0_H0_o(11), SHA256_BLOCK_0_H0_o(10) => 
        SHA256_BLOCK_0_H0_o(10), SHA256_BLOCK_0_H0_o(9) => 
        SHA256_BLOCK_0_H0_o(9), SHA256_BLOCK_0_H0_o(8) => 
        SHA256_BLOCK_0_H0_o(8), SHA256_BLOCK_0_H0_o(7) => 
        SHA256_BLOCK_0_H0_o(7), SHA256_BLOCK_0_H0_o(6) => 
        SHA256_BLOCK_0_H0_o(6), SHA256_BLOCK_0_H0_o(5) => 
        SHA256_BLOCK_0_H0_o(5), SHA256_BLOCK_0_H0_o(4) => 
        SHA256_BLOCK_0_H0_o(4), SHA256_BLOCK_0_H0_o(3) => 
        SHA256_BLOCK_0_H0_o(3), SHA256_BLOCK_0_H0_o(2) => 
        SHA256_BLOCK_0_H0_o(2), SHA256_BLOCK_0_H0_o(1) => 
        SHA256_BLOCK_0_H0_o(1), SHA256_BLOCK_0_H0_o(0) => 
        SHA256_BLOCK_0_H0_o(0), 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, wen_or_i_3_i_0 => 
        wen_or_i_3_i_0, data_out_ready => data_out_ready, ren_pos
         => \ren_pos\, AHB_slave_dummy_0_read_en => 
        AHB_slave_dummy_0_read_en, start_wen => start_wen);
    
    \reg_1x32_7\ : reg_1x32_7
      port map(line(31) => line_6_31, line(30) => line_6_30, 
        line(29) => line_6_29, line(28) => line_6_28, line(27)
         => line_6_27, line(26) => line_6_26, line(25) => 
        line_6_25, line(24) => line_6_24, line(23) => 
        \line_0[23]\, line(22) => line_6_22, line(21) => 
        line_6_21, line(20) => line_6_20, line(19) => line_6_19, 
        line(18) => line_6_18, line(17) => line_6_17, line(16)
         => line_6_16, line(15) => line_6_15, line(14) => 
        line_6_14, line(13) => \line_0[13]\, line(12) => 
        \line_4[12]\, line(11) => line_6_11, line(10) => 
        line_6_10, line(9) => line_6_9, line(8) => \line_4[8]\, 
        line(7) => line_6_7, line(6) => line_6_6, line(5) => 
        \line_0[5]\, line(4) => line_6_4, line(3) => line_6_3, 
        line(2) => line_6_2, line(1) => line_6_1, line(0) => 
        \line_0[0]\, SHA256_BLOCK_0_H7_o(31) => 
        SHA256_BLOCK_0_H7_o(31), SHA256_BLOCK_0_H7_o(30) => 
        SHA256_BLOCK_0_H7_o(30), SHA256_BLOCK_0_H7_o(29) => 
        SHA256_BLOCK_0_H7_o(29), SHA256_BLOCK_0_H7_o(28) => 
        SHA256_BLOCK_0_H7_o(28), SHA256_BLOCK_0_H7_o(27) => 
        SHA256_BLOCK_0_H7_o(27), SHA256_BLOCK_0_H7_o(26) => 
        SHA256_BLOCK_0_H7_o(26), SHA256_BLOCK_0_H7_o(25) => 
        SHA256_BLOCK_0_H7_o(25), SHA256_BLOCK_0_H7_o(24) => 
        SHA256_BLOCK_0_H7_o(24), SHA256_BLOCK_0_H7_o(23) => 
        SHA256_BLOCK_0_H7_o(23), SHA256_BLOCK_0_H7_o(22) => 
        SHA256_BLOCK_0_H7_o(22), SHA256_BLOCK_0_H7_o(21) => 
        SHA256_BLOCK_0_H7_o(21), SHA256_BLOCK_0_H7_o(20) => 
        SHA256_BLOCK_0_H7_o(20), SHA256_BLOCK_0_H7_o(19) => 
        SHA256_BLOCK_0_H7_o(19), SHA256_BLOCK_0_H7_o(18) => 
        SHA256_BLOCK_0_H7_o(18), SHA256_BLOCK_0_H7_o(17) => 
        SHA256_BLOCK_0_H7_o(17), SHA256_BLOCK_0_H7_o(16) => 
        SHA256_BLOCK_0_H7_o(16), SHA256_BLOCK_0_H7_o(15) => 
        SHA256_BLOCK_0_H7_o(15), SHA256_BLOCK_0_H7_o(14) => 
        SHA256_BLOCK_0_H7_o(14), SHA256_BLOCK_0_H7_o(13) => 
        SHA256_BLOCK_0_H7_o(13), SHA256_BLOCK_0_H7_o(12) => 
        SHA256_BLOCK_0_H7_o(12), SHA256_BLOCK_0_H7_o(11) => 
        SHA256_BLOCK_0_H7_o(11), SHA256_BLOCK_0_H7_o(10) => 
        SHA256_BLOCK_0_H7_o(10), SHA256_BLOCK_0_H7_o(9) => 
        SHA256_BLOCK_0_H7_o(9), SHA256_BLOCK_0_H7_o(8) => 
        SHA256_BLOCK_0_H7_o(8), SHA256_BLOCK_0_H7_o(7) => 
        SHA256_BLOCK_0_H7_o(7), SHA256_BLOCK_0_H7_o(6) => 
        SHA256_BLOCK_0_H7_o(6), SHA256_BLOCK_0_H7_o(5) => 
        SHA256_BLOCK_0_H7_o(5), SHA256_BLOCK_0_H7_o(4) => 
        SHA256_BLOCK_0_H7_o(4), SHA256_BLOCK_0_H7_o(3) => 
        SHA256_BLOCK_0_H7_o(3), SHA256_BLOCK_0_H7_o(2) => 
        SHA256_BLOCK_0_H7_o(2), SHA256_BLOCK_0_H7_o(1) => 
        SHA256_BLOCK_0_H7_o(1), SHA256_BLOCK_0_H7_o(0) => 
        SHA256_BLOCK_0_H7_o(0), 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, wen_or_i_3_i_0 => 
        wen_or_i_3_i_0, data_out_ready => data_out_ready);
    
    \reg_1x32_6\ : reg_1x32_6
      port map(line(31) => \line[31]\, line(30) => line_5_30, 
        line(29) => line_5_29, line(28) => \line_2[28]\, line(27)
         => line_5_27, line(26) => line_5_26, line(25) => 
        line_5_25, line(24) => line_5_24, line(23) => 
        \line_4[23]\, line(22) => line_5_22, line(21) => 
        line_5_21, line(20) => line_5_20, line(19) => line_5_19, 
        line(18) => line_5_18, line(17) => line_5_17, line(16)
         => line_5_16, line(15) => line_5_15, line(14) => 
        line_5_14, line(13) => \line_4[13]\, line(12) => 
        \line_0[12]\, line(11) => line_5_11, line(10) => 
        line_5_10, line(9) => line_5_9, line(8) => \line_0[8]\, 
        line(7) => line_5_7, line(6) => line_5_6, line(5) => 
        \line_4[5]\, line(4) => line_5_4, line(3) => line_5_3, 
        line(2) => line_5_2, line(1) => line_5_1, line(0) => 
        \line_4[0]\, SHA256_BLOCK_0_H6_o(31) => 
        SHA256_BLOCK_0_H6_o(31), SHA256_BLOCK_0_H6_o(30) => 
        SHA256_BLOCK_0_H6_o(30), SHA256_BLOCK_0_H6_o(29) => 
        SHA256_BLOCK_0_H6_o(29), SHA256_BLOCK_0_H6_o(28) => 
        SHA256_BLOCK_0_H6_o(28), SHA256_BLOCK_0_H6_o(27) => 
        SHA256_BLOCK_0_H6_o(27), SHA256_BLOCK_0_H6_o(26) => 
        SHA256_BLOCK_0_H6_o(26), SHA256_BLOCK_0_H6_o(25) => 
        SHA256_BLOCK_0_H6_o(25), SHA256_BLOCK_0_H6_o(24) => 
        SHA256_BLOCK_0_H6_o(24), SHA256_BLOCK_0_H6_o(23) => 
        SHA256_BLOCK_0_H6_o(23), SHA256_BLOCK_0_H6_o(22) => 
        SHA256_BLOCK_0_H6_o(22), SHA256_BLOCK_0_H6_o(21) => 
        SHA256_BLOCK_0_H6_o(21), SHA256_BLOCK_0_H6_o(20) => 
        SHA256_BLOCK_0_H6_o(20), SHA256_BLOCK_0_H6_o(19) => 
        SHA256_BLOCK_0_H6_o(19), SHA256_BLOCK_0_H6_o(18) => 
        SHA256_BLOCK_0_H6_o(18), SHA256_BLOCK_0_H6_o(17) => 
        SHA256_BLOCK_0_H6_o(17), SHA256_BLOCK_0_H6_o(16) => 
        SHA256_BLOCK_0_H6_o(16), SHA256_BLOCK_0_H6_o(15) => 
        SHA256_BLOCK_0_H6_o(15), SHA256_BLOCK_0_H6_o(14) => 
        SHA256_BLOCK_0_H6_o(14), SHA256_BLOCK_0_H6_o(13) => 
        SHA256_BLOCK_0_H6_o(13), SHA256_BLOCK_0_H6_o(12) => 
        SHA256_BLOCK_0_H6_o(12), SHA256_BLOCK_0_H6_o(11) => 
        SHA256_BLOCK_0_H6_o(11), SHA256_BLOCK_0_H6_o(10) => 
        SHA256_BLOCK_0_H6_o(10), SHA256_BLOCK_0_H6_o(9) => 
        SHA256_BLOCK_0_H6_o(9), SHA256_BLOCK_0_H6_o(8) => 
        SHA256_BLOCK_0_H6_o(8), SHA256_BLOCK_0_H6_o(7) => 
        SHA256_BLOCK_0_H6_o(7), SHA256_BLOCK_0_H6_o(6) => 
        SHA256_BLOCK_0_H6_o(6), SHA256_BLOCK_0_H6_o(5) => 
        SHA256_BLOCK_0_H6_o(5), SHA256_BLOCK_0_H6_o(4) => 
        SHA256_BLOCK_0_H6_o(4), SHA256_BLOCK_0_H6_o(3) => 
        SHA256_BLOCK_0_H6_o(3), SHA256_BLOCK_0_H6_o(2) => 
        SHA256_BLOCK_0_H6_o(2), SHA256_BLOCK_0_H6_o(1) => 
        SHA256_BLOCK_0_H6_o(1), SHA256_BLOCK_0_H6_o(0) => 
        SHA256_BLOCK_0_H6_o(0), 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, wen_or_i_3_i_0 => 
        wen_or_i_3_i_0, data_out_ready => data_out_ready);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \reg_1x32_5\ : reg_1x32_5
      port map(line(31) => line_5_31, line(30) => line_4_30, 
        line(29) => line_4_29, line(28) => line_5_28, line(27)
         => line_4_27, line(26) => line_4_26, line(25) => 
        line_4_25, line(24) => line_4_24, line(23) => 
        \line_2[23]\, line(22) => line_4_22, line(21) => 
        line_4_21, line(20) => line_4_20, line(19) => line_4_19, 
        line(18) => line_4_18, line(17) => line_4_17, line(16)
         => line_4_16, line(15) => line_4_15, line(14) => 
        line_4_14, line(13) => \line_2[13]\, line(12) => 
        \line_6[12]\, line(11) => line_4_11, line(10) => 
        line_4_10, line(9) => line_4_9, line(8) => \line_6[8]\, 
        line(7) => line_4_7, line(6) => line_4_6, line(5) => 
        \line_2[5]\, line(4) => line_4_4, line(3) => line_4_3, 
        line(2) => line_4_2, line(1) => line_4_1, line(0) => 
        \line_2[0]\, SHA256_BLOCK_0_H5_o(31) => 
        SHA256_BLOCK_0_H5_o(31), SHA256_BLOCK_0_H5_o(30) => 
        SHA256_BLOCK_0_H5_o(30), SHA256_BLOCK_0_H5_o(29) => 
        SHA256_BLOCK_0_H5_o(29), SHA256_BLOCK_0_H5_o(28) => 
        SHA256_BLOCK_0_H5_o(28), SHA256_BLOCK_0_H5_o(27) => 
        SHA256_BLOCK_0_H5_o(27), SHA256_BLOCK_0_H5_o(26) => 
        SHA256_BLOCK_0_H5_o(26), SHA256_BLOCK_0_H5_o(25) => 
        SHA256_BLOCK_0_H5_o(25), SHA256_BLOCK_0_H5_o(24) => 
        SHA256_BLOCK_0_H5_o(24), SHA256_BLOCK_0_H5_o(23) => 
        SHA256_BLOCK_0_H5_o(23), SHA256_BLOCK_0_H5_o(22) => 
        SHA256_BLOCK_0_H5_o(22), SHA256_BLOCK_0_H5_o(21) => 
        SHA256_BLOCK_0_H5_o(21), SHA256_BLOCK_0_H5_o(20) => 
        SHA256_BLOCK_0_H5_o(20), SHA256_BLOCK_0_H5_o(19) => 
        SHA256_BLOCK_0_H5_o(19), SHA256_BLOCK_0_H5_o(18) => 
        SHA256_BLOCK_0_H5_o(18), SHA256_BLOCK_0_H5_o(17) => 
        SHA256_BLOCK_0_H5_o(17), SHA256_BLOCK_0_H5_o(16) => 
        SHA256_BLOCK_0_H5_o(16), SHA256_BLOCK_0_H5_o(15) => 
        SHA256_BLOCK_0_H5_o(15), SHA256_BLOCK_0_H5_o(14) => 
        SHA256_BLOCK_0_H5_o(14), SHA256_BLOCK_0_H5_o(13) => 
        SHA256_BLOCK_0_H5_o(13), SHA256_BLOCK_0_H5_o(12) => 
        SHA256_BLOCK_0_H5_o(12), SHA256_BLOCK_0_H5_o(11) => 
        SHA256_BLOCK_0_H5_o(11), SHA256_BLOCK_0_H5_o(10) => 
        SHA256_BLOCK_0_H5_o(10), SHA256_BLOCK_0_H5_o(9) => 
        SHA256_BLOCK_0_H5_o(9), SHA256_BLOCK_0_H5_o(8) => 
        SHA256_BLOCK_0_H5_o(8), SHA256_BLOCK_0_H5_o(7) => 
        SHA256_BLOCK_0_H5_o(7), SHA256_BLOCK_0_H5_o(6) => 
        SHA256_BLOCK_0_H5_o(6), SHA256_BLOCK_0_H5_o(5) => 
        SHA256_BLOCK_0_H5_o(5), SHA256_BLOCK_0_H5_o(4) => 
        SHA256_BLOCK_0_H5_o(4), SHA256_BLOCK_0_H5_o(3) => 
        SHA256_BLOCK_0_H5_o(3), SHA256_BLOCK_0_H5_o(2) => 
        SHA256_BLOCK_0_H5_o(2), SHA256_BLOCK_0_H5_o(1) => 
        SHA256_BLOCK_0_H5_o(1), SHA256_BLOCK_0_H5_o(0) => 
        SHA256_BLOCK_0_H5_o(0), 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, wen_or_i_3_i_0 => 
        wen_or_i_3_i_0, data_out_ready => data_out_ready);
    
    \reg_1x32_2\ : reg_1x32_2
      port map(line(31) => \line_0[31]\, line(30) => line_1_30, 
        line(29) => line_1_29, line(28) => \line_1[28]\, line(27)
         => line_1_27, line(26) => line_1_26, line(25) => 
        line_1_25, line(24) => line_1_24, line(23) => 
        \line_3[23]\, line(22) => line_1_22, line(21) => 
        line_1_21, line(20) => line_1_20, line(19) => line_1_19, 
        line(18) => line_1_18, line(17) => line_1_17, line(16)
         => line_1_16, line(15) => line_1_15, line(14) => 
        line_1_14, line(13) => \line_3[13]\, line(12) => 
        \line[12]\, line(11) => line_1_11, line(10) => line_1_10, 
        line(9) => line_1_9, line(8) => \line[8]\, line(7) => 
        line_1_7, line(6) => line_1_6, line(5) => \line_3[5]\, 
        line(4) => line_1_4, line(3) => line_1_3, line(2) => 
        line_1_2, line(1) => line_1_1, line(0) => \line_3[0]\, 
        SHA256_BLOCK_0_H2_o(31) => SHA256_BLOCK_0_H2_o(31), 
        SHA256_BLOCK_0_H2_o(30) => SHA256_BLOCK_0_H2_o(30), 
        SHA256_BLOCK_0_H2_o(29) => SHA256_BLOCK_0_H2_o(29), 
        SHA256_BLOCK_0_H2_o(28) => SHA256_BLOCK_0_H2_o(28), 
        SHA256_BLOCK_0_H2_o(27) => SHA256_BLOCK_0_H2_o(27), 
        SHA256_BLOCK_0_H2_o(26) => SHA256_BLOCK_0_H2_o(26), 
        SHA256_BLOCK_0_H2_o(25) => SHA256_BLOCK_0_H2_o(25), 
        SHA256_BLOCK_0_H2_o(24) => SHA256_BLOCK_0_H2_o(24), 
        SHA256_BLOCK_0_H2_o(23) => SHA256_BLOCK_0_H2_o(23), 
        SHA256_BLOCK_0_H2_o(22) => SHA256_BLOCK_0_H2_o(22), 
        SHA256_BLOCK_0_H2_o(21) => SHA256_BLOCK_0_H2_o(21), 
        SHA256_BLOCK_0_H2_o(20) => SHA256_BLOCK_0_H2_o(20), 
        SHA256_BLOCK_0_H2_o(19) => SHA256_BLOCK_0_H2_o(19), 
        SHA256_BLOCK_0_H2_o(18) => SHA256_BLOCK_0_H2_o(18), 
        SHA256_BLOCK_0_H2_o(17) => SHA256_BLOCK_0_H2_o(17), 
        SHA256_BLOCK_0_H2_o(16) => SHA256_BLOCK_0_H2_o(16), 
        SHA256_BLOCK_0_H2_o(15) => SHA256_BLOCK_0_H2_o(15), 
        SHA256_BLOCK_0_H2_o(14) => SHA256_BLOCK_0_H2_o(14), 
        SHA256_BLOCK_0_H2_o(13) => SHA256_BLOCK_0_H2_o(13), 
        SHA256_BLOCK_0_H2_o(12) => SHA256_BLOCK_0_H2_o(12), 
        SHA256_BLOCK_0_H2_o(11) => SHA256_BLOCK_0_H2_o(11), 
        SHA256_BLOCK_0_H2_o(10) => SHA256_BLOCK_0_H2_o(10), 
        SHA256_BLOCK_0_H2_o(9) => SHA256_BLOCK_0_H2_o(9), 
        SHA256_BLOCK_0_H2_o(8) => SHA256_BLOCK_0_H2_o(8), 
        SHA256_BLOCK_0_H2_o(7) => SHA256_BLOCK_0_H2_o(7), 
        SHA256_BLOCK_0_H2_o(6) => SHA256_BLOCK_0_H2_o(6), 
        SHA256_BLOCK_0_H2_o(5) => SHA256_BLOCK_0_H2_o(5), 
        SHA256_BLOCK_0_H2_o(4) => SHA256_BLOCK_0_H2_o(4), 
        SHA256_BLOCK_0_H2_o(3) => SHA256_BLOCK_0_H2_o(3), 
        SHA256_BLOCK_0_H2_o(2) => SHA256_BLOCK_0_H2_o(2), 
        SHA256_BLOCK_0_H2_o(1) => SHA256_BLOCK_0_H2_o(1), 
        SHA256_BLOCK_0_H2_o(0) => SHA256_BLOCK_0_H2_o(0), 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, wen_or_i_3_i_0 => 
        wen_or_i_3_i_0, data_out_ready => data_out_ready);
    
    \reg_1x32_8\ : reg_1x32_8
      port map(line(2) => line_7_2, line(1) => line_7_1, line(0)
         => \line_7[0]\, CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, 
        SHA256_Module_0_error_o => SHA256_Module_0_error_o, 
        wen_or_i_3_i_0 => wen_or_i_3_i_0, data_out_ready => 
        data_out_ready, SHA256_Module_0_di_req_o => 
        SHA256_Module_0_di_req_o, SHA256_Module_0_do_valid_o => 
        SHA256_Module_0_do_valid_o);
    
    \reg_1x32_3\ : reg_1x32_3
      port map(line(31) => line_4_31, line(30) => line_2_30, 
        line(29) => line_2_29, line(28) => line_4_28, line(27)
         => line_2_27, line(26) => line_2_26, line(25) => 
        line_2_25, line(24) => line_2_24, line(23) => \line[23]\, 
        line(22) => line_2_22, line(21) => line_2_21, line(20)
         => line_2_20, line(19) => line_2_19, line(18) => 
        line_2_18, line(17) => line_2_17, line(16) => line_2_16, 
        line(15) => line_2_15, line(14) => line_2_14, line(13)
         => \line[13]\, line(12) => \line_3[12]\, line(11) => 
        line_2_11, line(10) => line_2_10, line(9) => line_2_9, 
        line(8) => \line_3[8]\, line(7) => line_2_7, line(6) => 
        line_2_6, line(5) => \line[5]\, line(4) => line_2_4, 
        line(3) => line_2_3, line(2) => line_2_2, line(1) => 
        line_2_1, line(0) => \line[0]\, SHA256_BLOCK_0_H3_o(31)
         => SHA256_BLOCK_0_H3_o(31), SHA256_BLOCK_0_H3_o(30) => 
        SHA256_BLOCK_0_H3_o(30), SHA256_BLOCK_0_H3_o(29) => 
        SHA256_BLOCK_0_H3_o(29), SHA256_BLOCK_0_H3_o(28) => 
        SHA256_BLOCK_0_H3_o(28), SHA256_BLOCK_0_H3_o(27) => 
        SHA256_BLOCK_0_H3_o(27), SHA256_BLOCK_0_H3_o(26) => 
        SHA256_BLOCK_0_H3_o(26), SHA256_BLOCK_0_H3_o(25) => 
        SHA256_BLOCK_0_H3_o(25), SHA256_BLOCK_0_H3_o(24) => 
        SHA256_BLOCK_0_H3_o(24), SHA256_BLOCK_0_H3_o(23) => 
        SHA256_BLOCK_0_H3_o(23), SHA256_BLOCK_0_H3_o(22) => 
        SHA256_BLOCK_0_H3_o(22), SHA256_BLOCK_0_H3_o(21) => 
        SHA256_BLOCK_0_H3_o(21), SHA256_BLOCK_0_H3_o(20) => 
        SHA256_BLOCK_0_H3_o(20), SHA256_BLOCK_0_H3_o(19) => 
        SHA256_BLOCK_0_H3_o(19), SHA256_BLOCK_0_H3_o(18) => 
        SHA256_BLOCK_0_H3_o(18), SHA256_BLOCK_0_H3_o(17) => 
        SHA256_BLOCK_0_H3_o(17), SHA256_BLOCK_0_H3_o(16) => 
        SHA256_BLOCK_0_H3_o(16), SHA256_BLOCK_0_H3_o(15) => 
        SHA256_BLOCK_0_H3_o(15), SHA256_BLOCK_0_H3_o(14) => 
        SHA256_BLOCK_0_H3_o(14), SHA256_BLOCK_0_H3_o(13) => 
        SHA256_BLOCK_0_H3_o(13), SHA256_BLOCK_0_H3_o(12) => 
        SHA256_BLOCK_0_H3_o(12), SHA256_BLOCK_0_H3_o(11) => 
        SHA256_BLOCK_0_H3_o(11), SHA256_BLOCK_0_H3_o(10) => 
        SHA256_BLOCK_0_H3_o(10), SHA256_BLOCK_0_H3_o(9) => 
        SHA256_BLOCK_0_H3_o(9), SHA256_BLOCK_0_H3_o(8) => 
        SHA256_BLOCK_0_H3_o(8), SHA256_BLOCK_0_H3_o(7) => 
        SHA256_BLOCK_0_H3_o(7), SHA256_BLOCK_0_H3_o(6) => 
        SHA256_BLOCK_0_H3_o(6), SHA256_BLOCK_0_H3_o(5) => 
        SHA256_BLOCK_0_H3_o(5), SHA256_BLOCK_0_H3_o(4) => 
        SHA256_BLOCK_0_H3_o(4), SHA256_BLOCK_0_H3_o(3) => 
        SHA256_BLOCK_0_H3_o(3), SHA256_BLOCK_0_H3_o(2) => 
        SHA256_BLOCK_0_H3_o(2), SHA256_BLOCK_0_H3_o(1) => 
        SHA256_BLOCK_0_H3_o(1), SHA256_BLOCK_0_H3_o(0) => 
        SHA256_BLOCK_0_H3_o(0), 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, wen_or_i_3_i_0 => 
        wen_or_i_3_i_0, data_out_ready => data_out_ready);
    
    \reg_1x32_4\ : reg_1x32_4
      port map(line(31) => \line_2[31]\, line(30) => line_3_30, 
        line(29) => line_3_29, line(28) => \line[28]\, line(27)
         => line_3_27, line(26) => line_3_26, line(25) => 
        line_3_25, line(24) => line_3_24, line(23) => 
        \line_6[23]\, line(22) => line_3_22, line(21) => 
        line_3_21, line(20) => line_3_20, line(19) => line_3_19, 
        line(18) => line_3_18, line(17) => line_3_17, line(16)
         => line_3_16, line(15) => line_3_15, line(14) => 
        line_3_14, line(13) => \line_6[13]\, line(12) => 
        \line_2[12]\, line(11) => line_3_11, line(10) => 
        line_3_10, line(9) => line_3_9, line(8) => \line_2[8]\, 
        line(7) => line_3_7, line(6) => line_3_6, line(5) => 
        \line_6[5]\, line(4) => line_3_4, line(3) => line_3_3, 
        line(2) => line_3_2, line(1) => line_3_1, line(0) => 
        \line_6[0]\, SHA256_BLOCK_0_H4_o(31) => 
        SHA256_BLOCK_0_H4_o(31), SHA256_BLOCK_0_H4_o(30) => 
        SHA256_BLOCK_0_H4_o(30), SHA256_BLOCK_0_H4_o(29) => 
        SHA256_BLOCK_0_H4_o(29), SHA256_BLOCK_0_H4_o(28) => 
        SHA256_BLOCK_0_H4_o(28), SHA256_BLOCK_0_H4_o(27) => 
        SHA256_BLOCK_0_H4_o(27), SHA256_BLOCK_0_H4_o(26) => 
        SHA256_BLOCK_0_H4_o(26), SHA256_BLOCK_0_H4_o(25) => 
        SHA256_BLOCK_0_H4_o(25), SHA256_BLOCK_0_H4_o(24) => 
        SHA256_BLOCK_0_H4_o(24), SHA256_BLOCK_0_H4_o(23) => 
        SHA256_BLOCK_0_H4_o(23), SHA256_BLOCK_0_H4_o(22) => 
        SHA256_BLOCK_0_H4_o(22), SHA256_BLOCK_0_H4_o(21) => 
        SHA256_BLOCK_0_H4_o(21), SHA256_BLOCK_0_H4_o(20) => 
        SHA256_BLOCK_0_H4_o(20), SHA256_BLOCK_0_H4_o(19) => 
        SHA256_BLOCK_0_H4_o(19), SHA256_BLOCK_0_H4_o(18) => 
        SHA256_BLOCK_0_H4_o(18), SHA256_BLOCK_0_H4_o(17) => 
        SHA256_BLOCK_0_H4_o(17), SHA256_BLOCK_0_H4_o(16) => 
        SHA256_BLOCK_0_H4_o(16), SHA256_BLOCK_0_H4_o(15) => 
        SHA256_BLOCK_0_H4_o(15), SHA256_BLOCK_0_H4_o(14) => 
        SHA256_BLOCK_0_H4_o(14), SHA256_BLOCK_0_H4_o(13) => 
        SHA256_BLOCK_0_H4_o(13), SHA256_BLOCK_0_H4_o(12) => 
        SHA256_BLOCK_0_H4_o(12), SHA256_BLOCK_0_H4_o(11) => 
        SHA256_BLOCK_0_H4_o(11), SHA256_BLOCK_0_H4_o(10) => 
        SHA256_BLOCK_0_H4_o(10), SHA256_BLOCK_0_H4_o(9) => 
        SHA256_BLOCK_0_H4_o(9), SHA256_BLOCK_0_H4_o(8) => 
        SHA256_BLOCK_0_H4_o(8), SHA256_BLOCK_0_H4_o(7) => 
        SHA256_BLOCK_0_H4_o(7), SHA256_BLOCK_0_H4_o(6) => 
        SHA256_BLOCK_0_H4_o(6), SHA256_BLOCK_0_H4_o(5) => 
        SHA256_BLOCK_0_H4_o(5), SHA256_BLOCK_0_H4_o(4) => 
        SHA256_BLOCK_0_H4_o(4), SHA256_BLOCK_0_H4_o(3) => 
        SHA256_BLOCK_0_H4_o(3), SHA256_BLOCK_0_H4_o(2) => 
        SHA256_BLOCK_0_H4_o(2), SHA256_BLOCK_0_H4_o(1) => 
        SHA256_BLOCK_0_H4_o(1), SHA256_BLOCK_0_H4_o(0) => 
        SHA256_BLOCK_0_H4_o(0), 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, wen_or_i_3_i_0 => 
        wen_or_i_3_i_0, data_out_ready => data_out_ready);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity reg1_highonly is

    port( CertificationSystem_sb_0_GPIO_9_M2F     : in    std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F_i_0 : out   std_logic;
          start_wen                               : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0    : in    std_logic;
          SHA256_BLOCK_0_start_o                  : in    std_logic
        );

end reg1_highonly;

architecture DEF_ARCH of reg1_highonly is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal CertificationSystem_sb_0_GPIO_9_M2F_i_0_net_1, 
        \start_wen\, VCC_net_1, \data_2\, GND_net_1 : std_logic;

begin 

    CertificationSystem_sb_0_GPIO_9_M2F_i_0 <= 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0_net_1;
    start_wen <= \start_wen\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    data : SLE
      port map(D => \data_2\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \start_wen\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \CertificationSystem_sb_0_GPIO_9_M2F_i_0\ : CFG1
      generic map(INIT => "01")

      port map(A => CertificationSystem_sb_0_GPIO_9_M2F, Y => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0_net_1);
    
    data_2 : CFG4
      generic map(INIT => x"0E0A")

      port map(A => SHA256_BLOCK_0_start_o, B => \start_wen\, C
         => CertificationSystem_sb_0_GPIO_9_M2F_i_0_net_1, D => 
        CertificationSystem_sb_0_GPIO_9_M2F, Y => \data_2\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity SHA256_Module is

    port( result_addr_net_0                         : in    std_logic_vector(3 downto 0);
          line_7                                    : out   std_logic_vector(2 downto 1);
          waddr_in_net_0                            : in    std_logic_vector(4 downto 0);
          SHA256_Module_0_data_out_5                : out   std_logic;
          SHA256_Module_0_data_out_13               : out   std_logic;
          SHA256_Module_0_data_out_12               : out   std_logic;
          SHA256_Module_0_data_out_23               : out   std_logic;
          SHA256_Module_0_data_out_8                : out   std_logic;
          SHA256_Module_0_data_out_0                : out   std_logic;
          line_0_d0                                 : out   std_logic;
          line_1_d0                                 : out   std_logic;
          line_2_d0                                 : out   std_logic;
          line_3_d0                                 : out   std_logic;
          line_5_d0                                 : out   std_logic;
          line_6_d0                                 : out   std_logic;
          line_8                                    : out   std_logic;
          line_9                                    : out   std_logic;
          line_10                                   : out   std_logic;
          line_13                                   : out   std_logic;
          line_14                                   : out   std_logic;
          line_15                                   : out   std_logic;
          line_16                                   : out   std_logic;
          line_17                                   : out   std_logic;
          line_18                                   : out   std_logic;
          line_19                                   : out   std_logic;
          line_20                                   : out   std_logic;
          line_21                                   : out   std_logic;
          line_23                                   : out   std_logic;
          line_24                                   : out   std_logic;
          line_25                                   : out   std_logic;
          line_26                                   : out   std_logic;
          line_28                                   : out   std_logic;
          line_29                                   : out   std_logic;
          line_27                                   : out   std_logic;
          line_30                                   : out   std_logic;
          line_3_0                                  : out   std_logic;
          line_3_1                                  : out   std_logic;
          line_3_2                                  : out   std_logic;
          line_3_3                                  : out   std_logic;
          line_3_5                                  : out   std_logic;
          line_3_6                                  : out   std_logic;
          line_3_8                                  : out   std_logic;
          line_3_9                                  : out   std_logic;
          line_3_10                                 : out   std_logic;
          line_3_13                                 : out   std_logic;
          line_3_14                                 : out   std_logic;
          line_3_15                                 : out   std_logic;
          line_3_16                                 : out   std_logic;
          line_3_17                                 : out   std_logic;
          line_3_18                                 : out   std_logic;
          line_3_19                                 : out   std_logic;
          line_3_20                                 : out   std_logic;
          line_3_21                                 : out   std_logic;
          line_3_23                                 : out   std_logic;
          line_3_24                                 : out   std_logic;
          line_3_25                                 : out   std_logic;
          line_3_26                                 : out   std_logic;
          line_3_28                                 : out   std_logic;
          line_3_29                                 : out   std_logic;
          line_0_0                                  : out   std_logic;
          line_0_1                                  : out   std_logic;
          line_0_2                                  : out   std_logic;
          line_0_3                                  : out   std_logic;
          line_0_5                                  : out   std_logic;
          line_0_6                                  : out   std_logic;
          line_0_8                                  : out   std_logic;
          line_0_9                                  : out   std_logic;
          line_0_10                                 : out   std_logic;
          line_0_13                                 : out   std_logic;
          line_0_14                                 : out   std_logic;
          line_0_15                                 : out   std_logic;
          line_0_16                                 : out   std_logic;
          line_0_17                                 : out   std_logic;
          line_0_18                                 : out   std_logic;
          line_0_19                                 : out   std_logic;
          line_0_20                                 : out   std_logic;
          line_0_21                                 : out   std_logic;
          line_0_23                                 : out   std_logic;
          line_0_24                                 : out   std_logic;
          line_0_25                                 : out   std_logic;
          line_0_26                                 : out   std_logic;
          line_0_28                                 : out   std_logic;
          line_0_29                                 : out   std_logic;
          line_0_27                                 : out   std_logic;
          line_0_30                                 : out   std_logic;
          line_4_0                                  : out   std_logic;
          line_4_1                                  : out   std_logic;
          line_4_2                                  : out   std_logic;
          line_4_3                                  : out   std_logic;
          line_4_5                                  : out   std_logic;
          line_4_6                                  : out   std_logic;
          line_4_8                                  : out   std_logic;
          line_4_9                                  : out   std_logic;
          line_4_10                                 : out   std_logic;
          line_4_13                                 : out   std_logic;
          line_4_14                                 : out   std_logic;
          line_4_15                                 : out   std_logic;
          line_4_16                                 : out   std_logic;
          line_4_17                                 : out   std_logic;
          line_4_18                                 : out   std_logic;
          line_4_19                                 : out   std_logic;
          line_4_20                                 : out   std_logic;
          line_4_21                                 : out   std_logic;
          line_4_23                                 : out   std_logic;
          line_4_24                                 : out   std_logic;
          line_4_25                                 : out   std_logic;
          line_4_26                                 : out   std_logic;
          line_4_28                                 : out   std_logic;
          line_4_29                                 : out   std_logic;
          line_1_0                                  : out   std_logic;
          line_1_1                                  : out   std_logic;
          line_1_2                                  : out   std_logic;
          line_1_3                                  : out   std_logic;
          line_1_5                                  : out   std_logic;
          line_1_6                                  : out   std_logic;
          line_1_8                                  : out   std_logic;
          line_1_9                                  : out   std_logic;
          line_1_10                                 : out   std_logic;
          line_1_13                                 : out   std_logic;
          line_1_14                                 : out   std_logic;
          line_1_15                                 : out   std_logic;
          line_1_16                                 : out   std_logic;
          line_1_17                                 : out   std_logic;
          line_1_18                                 : out   std_logic;
          line_1_19                                 : out   std_logic;
          line_1_20                                 : out   std_logic;
          line_1_21                                 : out   std_logic;
          line_1_23                                 : out   std_logic;
          line_1_24                                 : out   std_logic;
          line_1_25                                 : out   std_logic;
          line_1_26                                 : out   std_logic;
          line_1_28                                 : out   std_logic;
          line_1_29                                 : out   std_logic;
          line_1_27                                 : out   std_logic;
          line_1_30                                 : out   std_logic;
          line_5_0                                  : out   std_logic;
          line_5_1                                  : out   std_logic;
          line_5_2                                  : out   std_logic;
          line_5_3                                  : out   std_logic;
          line_5_5                                  : out   std_logic;
          line_5_6                                  : out   std_logic;
          line_5_8                                  : out   std_logic;
          line_5_9                                  : out   std_logic;
          line_5_10                                 : out   std_logic;
          line_5_13                                 : out   std_logic;
          line_5_14                                 : out   std_logic;
          line_5_15                                 : out   std_logic;
          line_5_16                                 : out   std_logic;
          line_5_17                                 : out   std_logic;
          line_5_18                                 : out   std_logic;
          line_5_19                                 : out   std_logic;
          line_5_20                                 : out   std_logic;
          line_5_21                                 : out   std_logic;
          line_5_23                                 : out   std_logic;
          line_5_24                                 : out   std_logic;
          line_5_25                                 : out   std_logic;
          line_5_26                                 : out   std_logic;
          line_5_28                                 : out   std_logic;
          line_5_29                                 : out   std_logic;
          line_6_0                                  : out   std_logic;
          line_6_1                                  : out   std_logic;
          line_6_2                                  : out   std_logic;
          line_6_3                                  : out   std_logic;
          line_6_5                                  : out   std_logic;
          line_6_6                                  : out   std_logic;
          line_6_8                                  : out   std_logic;
          line_6_9                                  : out   std_logic;
          line_6_10                                 : out   std_logic;
          line_6_13                                 : out   std_logic;
          line_6_14                                 : out   std_logic;
          line_6_15                                 : out   std_logic;
          line_6_16                                 : out   std_logic;
          line_6_17                                 : out   std_logic;
          line_6_18                                 : out   std_logic;
          line_6_19                                 : out   std_logic;
          line_6_20                                 : out   std_logic;
          line_6_21                                 : out   std_logic;
          line_6_23                                 : out   std_logic;
          line_6_24                                 : out   std_logic;
          line_6_25                                 : out   std_logic;
          line_6_26                                 : out   std_logic;
          line_6_28                                 : out   std_logic;
          line_6_29                                 : out   std_logic;
          line_2_0                                  : out   std_logic;
          line_2_1                                  : out   std_logic;
          line_2_2                                  : out   std_logic;
          line_2_3                                  : out   std_logic;
          line_2_5                                  : out   std_logic;
          line_2_6                                  : out   std_logic;
          line_2_8                                  : out   std_logic;
          line_2_9                                  : out   std_logic;
          line_2_10                                 : out   std_logic;
          line_2_13                                 : out   std_logic;
          line_2_14                                 : out   std_logic;
          line_2_15                                 : out   std_logic;
          line_2_16                                 : out   std_logic;
          line_2_17                                 : out   std_logic;
          line_2_18                                 : out   std_logic;
          line_2_19                                 : out   std_logic;
          line_2_20                                 : out   std_logic;
          line_2_21                                 : out   std_logic;
          line_2_23                                 : out   std_logic;
          line_2_24                                 : out   std_logic;
          line_2_25                                 : out   std_logic;
          line_2_26                                 : out   std_logic;
          line_2_28                                 : out   std_logic;
          line_2_29                                 : out   std_logic;
          line_2_27                                 : out   std_logic;
          line_2_30                                 : out   std_logic;
          SHA256_Module_0_do_valid_o                : out   std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F       : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0      : in    std_logic;
          N_507                                     : out   std_logic;
          N_508                                     : out   std_logic;
          ren_pos                                   : out   std_logic;
          AHB_slave_dummy_0_read_en                 : in    std_logic;
          SHA256_Module_0_error_o                   : out   std_logic;
          SHA256_Module_0_di_req_o                  : out   std_logic;
          SHA256_Module_0_waiting_data              : out   std_logic;
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic;
          SHA256_Module_0_data_available            : out   std_logic;
          N_111_i_0                                 : in    std_logic;
          N_109_i_0                                 : in    std_logic;
          N_168_i_0                                 : in    std_logic;
          N_107_i_0                                 : in    std_logic;
          N_99_i_0                                  : in    std_logic;
          N_97_i_0                                  : in    std_logic;
          N_67_i_0                                  : in    std_logic;
          N_65_i_0                                  : in    std_logic;
          N_105_i_0                                 : in    std_logic;
          N_103_i_0                                 : in    std_logic;
          N_158_i_0                                 : in    std_logic;
          N_156_i_0                                 : in    std_logic;
          N_101_i_0                                 : in    std_logic;
          N_152_i_0                                 : in    std_logic;
          N_95_i_0                                  : in    std_logic;
          N_93_i_0                                  : in    std_logic;
          N_91_i_0                                  : in    std_logic;
          N_140_i_0                                 : in    std_logic;
          N_89_i_0                                  : in    std_logic;
          N_87_i_0                                  : in    std_logic;
          N_133_i_0                                 : in    std_logic;
          N_85_i_0                                  : in    std_logic;
          N_83_i_0                                  : in    std_logic;
          N_77_i_0                                  : in    std_logic;
          N_75_i_0                                  : in    std_logic;
          N_73_i_0                                  : in    std_logic;
          N_71_i_0                                  : in    std_logic;
          N_69_i_0                                  : in    std_logic;
          N_116_i_0                                 : in    std_logic;
          N_114_i_0                                 : in    std_logic;
          N_112_i_0                                 : in    std_logic;
          N_110_i_0                                 : in    std_logic;
          CertificationSystem_sb_0_GPIO_1_M2F       : in    std_logic;
          AHB_slave_dummy_0_write_en                : in    std_logic
        );

end SHA256_Module;

architecture DEF_ARCH of SHA256_Module is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SHA256_BLOCK
    port( SHA256_BLOCK_0_H0_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H1_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H2_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H3_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H4_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H5_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H6_o                       : out   std_logic_vector(31 downto 0);
          SHA256_BLOCK_0_H7_o                       : out   std_logic_vector(31 downto 0);
          waddr_in_net_0                            : in    std_logic_vector(4 downto 0) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0      : in    std_logic := 'U';
          SHA256_Module_0_di_req_o                  : out   std_logic;
          SHA256_BLOCK_0_do_valid_o                 : out   std_logic;
          SHA256_Module_0_waiting_data              : out   std_logic;
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic;
          SHA256_Module_0_error_o                   : out   std_logic;
          SHA256_BLOCK_0_start_o                    : out   std_logic;
          data_out_ready                            : out   std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F       : in    std_logic := 'U';
          SHA256_Module_0_data_available            : out   std_logic;
          N_111_i_0                                 : in    std_logic := 'U';
          N_109_i_0                                 : in    std_logic := 'U';
          N_168_i_0                                 : in    std_logic := 'U';
          N_107_i_0                                 : in    std_logic := 'U';
          N_99_i_0                                  : in    std_logic := 'U';
          N_97_i_0                                  : in    std_logic := 'U';
          N_67_i_0                                  : in    std_logic := 'U';
          N_65_i_0                                  : in    std_logic := 'U';
          CertificationSystem_sb_0_GPIO_9_M2F_i_0   : in    std_logic := 'U';
          N_105_i_0                                 : in    std_logic := 'U';
          N_103_i_0                                 : in    std_logic := 'U';
          N_158_i_0                                 : in    std_logic := 'U';
          N_156_i_0                                 : in    std_logic := 'U';
          N_101_i_0                                 : in    std_logic := 'U';
          N_152_i_0                                 : in    std_logic := 'U';
          N_95_i_0                                  : in    std_logic := 'U';
          N_93_i_0                                  : in    std_logic := 'U';
          N_91_i_0                                  : in    std_logic := 'U';
          N_140_i_0                                 : in    std_logic := 'U';
          N_89_i_0                                  : in    std_logic := 'U';
          N_87_i_0                                  : in    std_logic := 'U';
          N_133_i_0                                 : in    std_logic := 'U';
          N_85_i_0                                  : in    std_logic := 'U';
          N_83_i_0                                  : in    std_logic := 'U';
          N_77_i_0                                  : in    std_logic := 'U';
          N_75_i_0                                  : in    std_logic := 'U';
          N_73_i_0                                  : in    std_logic := 'U';
          N_71_i_0                                  : in    std_logic := 'U';
          N_69_i_0                                  : in    std_logic := 'U';
          N_116_i_0                                 : in    std_logic := 'U';
          N_114_i_0                                 : in    std_logic := 'U';
          N_112_i_0                                 : in    std_logic := 'U';
          N_110_i_0                                 : in    std_logic := 'U';
          CertificationSystem_sb_0_GPIO_1_M2F       : in    std_logic := 'U';
          AHB_slave_dummy_0_write_en                : in    std_logic := 'U'
        );
  end component;

  component reg9_1x32
    port( result_addr_net_0                    : in    std_logic_vector(3 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H0_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H1_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H2_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H3_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H4_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H5_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H6_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_BLOCK_0_H7_o                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          SHA256_Module_0_data_out_5           : out   std_logic;
          SHA256_Module_0_data_out_13          : out   std_logic;
          SHA256_Module_0_data_out_12          : out   std_logic;
          SHA256_Module_0_data_out_23          : out   std_logic;
          SHA256_Module_0_data_out_8           : out   std_logic;
          SHA256_Module_0_data_out_0           : out   std_logic;
          line_1_d0                            : out   std_logic;
          line_2_d0                            : out   std_logic;
          line_3_d0                            : out   std_logic;
          line_4_d0                            : out   std_logic;
          line_6_d0                            : out   std_logic;
          line_7_d0                            : out   std_logic;
          line_9                               : out   std_logic;
          line_10                              : out   std_logic;
          line_11                              : out   std_logic;
          line_14                              : out   std_logic;
          line_15                              : out   std_logic;
          line_16                              : out   std_logic;
          line_17                              : out   std_logic;
          line_18                              : out   std_logic;
          line_19                              : out   std_logic;
          line_20                              : out   std_logic;
          line_21                              : out   std_logic;
          line_22                              : out   std_logic;
          line_24                              : out   std_logic;
          line_25                              : out   std_logic;
          line_26                              : out   std_logic;
          line_27                              : out   std_logic;
          line_29                              : out   std_logic;
          line_30                              : out   std_logic;
          line_0_1                             : out   std_logic;
          line_0_2                             : out   std_logic;
          line_0_3                             : out   std_logic;
          line_0_4                             : out   std_logic;
          line_0_6                             : out   std_logic;
          line_0_7                             : out   std_logic;
          line_0_9                             : out   std_logic;
          line_0_10                            : out   std_logic;
          line_0_11                            : out   std_logic;
          line_0_14                            : out   std_logic;
          line_0_15                            : out   std_logic;
          line_0_16                            : out   std_logic;
          line_0_17                            : out   std_logic;
          line_0_18                            : out   std_logic;
          line_0_19                            : out   std_logic;
          line_0_20                            : out   std_logic;
          line_0_21                            : out   std_logic;
          line_0_22                            : out   std_logic;
          line_0_24                            : out   std_logic;
          line_0_25                            : out   std_logic;
          line_0_26                            : out   std_logic;
          line_0_27                            : out   std_logic;
          line_0_29                            : out   std_logic;
          line_0_30                            : out   std_logic;
          line_1_1                             : out   std_logic;
          line_1_2                             : out   std_logic;
          line_1_3                             : out   std_logic;
          line_1_4                             : out   std_logic;
          line_1_6                             : out   std_logic;
          line_1_7                             : out   std_logic;
          line_1_9                             : out   std_logic;
          line_1_10                            : out   std_logic;
          line_1_11                            : out   std_logic;
          line_1_14                            : out   std_logic;
          line_1_15                            : out   std_logic;
          line_1_16                            : out   std_logic;
          line_1_17                            : out   std_logic;
          line_1_18                            : out   std_logic;
          line_1_19                            : out   std_logic;
          line_1_20                            : out   std_logic;
          line_1_21                            : out   std_logic;
          line_1_22                            : out   std_logic;
          line_1_24                            : out   std_logic;
          line_1_25                            : out   std_logic;
          line_1_26                            : out   std_logic;
          line_1_27                            : out   std_logic;
          line_1_29                            : out   std_logic;
          line_1_30                            : out   std_logic;
          line_2_1                             : out   std_logic;
          line_2_2                             : out   std_logic;
          line_2_3                             : out   std_logic;
          line_2_4                             : out   std_logic;
          line_2_6                             : out   std_logic;
          line_2_7                             : out   std_logic;
          line_2_9                             : out   std_logic;
          line_2_10                            : out   std_logic;
          line_2_11                            : out   std_logic;
          line_2_14                            : out   std_logic;
          line_2_15                            : out   std_logic;
          line_2_16                            : out   std_logic;
          line_2_17                            : out   std_logic;
          line_2_18                            : out   std_logic;
          line_2_19                            : out   std_logic;
          line_2_20                            : out   std_logic;
          line_2_21                            : out   std_logic;
          line_2_22                            : out   std_logic;
          line_2_24                            : out   std_logic;
          line_2_25                            : out   std_logic;
          line_2_26                            : out   std_logic;
          line_2_27                            : out   std_logic;
          line_2_29                            : out   std_logic;
          line_2_30                            : out   std_logic;
          line_3_28                            : out   std_logic;
          line_3_31                            : out   std_logic;
          line_3_1                             : out   std_logic;
          line_3_2                             : out   std_logic;
          line_3_3                             : out   std_logic;
          line_3_4                             : out   std_logic;
          line_3_6                             : out   std_logic;
          line_3_7                             : out   std_logic;
          line_3_9                             : out   std_logic;
          line_3_10                            : out   std_logic;
          line_3_11                            : out   std_logic;
          line_3_14                            : out   std_logic;
          line_3_15                            : out   std_logic;
          line_3_16                            : out   std_logic;
          line_3_17                            : out   std_logic;
          line_3_18                            : out   std_logic;
          line_3_19                            : out   std_logic;
          line_3_20                            : out   std_logic;
          line_3_21                            : out   std_logic;
          line_3_22                            : out   std_logic;
          line_3_24                            : out   std_logic;
          line_3_25                            : out   std_logic;
          line_3_26                            : out   std_logic;
          line_3_27                            : out   std_logic;
          line_3_29                            : out   std_logic;
          line_3_30                            : out   std_logic;
          line_4_28                            : out   std_logic;
          line_4_31                            : out   std_logic;
          line_4_1                             : out   std_logic;
          line_4_2                             : out   std_logic;
          line_4_3                             : out   std_logic;
          line_4_4                             : out   std_logic;
          line_4_6                             : out   std_logic;
          line_4_7                             : out   std_logic;
          line_4_9                             : out   std_logic;
          line_4_10                            : out   std_logic;
          line_4_11                            : out   std_logic;
          line_4_14                            : out   std_logic;
          line_4_15                            : out   std_logic;
          line_4_16                            : out   std_logic;
          line_4_17                            : out   std_logic;
          line_4_18                            : out   std_logic;
          line_4_19                            : out   std_logic;
          line_4_20                            : out   std_logic;
          line_4_21                            : out   std_logic;
          line_4_22                            : out   std_logic;
          line_4_24                            : out   std_logic;
          line_4_25                            : out   std_logic;
          line_4_26                            : out   std_logic;
          line_4_27                            : out   std_logic;
          line_4_29                            : out   std_logic;
          line_4_30                            : out   std_logic;
          line_5_28                            : out   std_logic;
          line_5_31                            : out   std_logic;
          line_5_1                             : out   std_logic;
          line_5_2                             : out   std_logic;
          line_5_3                             : out   std_logic;
          line_5_4                             : out   std_logic;
          line_5_6                             : out   std_logic;
          line_5_7                             : out   std_logic;
          line_5_9                             : out   std_logic;
          line_5_10                            : out   std_logic;
          line_5_11                            : out   std_logic;
          line_5_14                            : out   std_logic;
          line_5_15                            : out   std_logic;
          line_5_16                            : out   std_logic;
          line_5_17                            : out   std_logic;
          line_5_18                            : out   std_logic;
          line_5_19                            : out   std_logic;
          line_5_20                            : out   std_logic;
          line_5_21                            : out   std_logic;
          line_5_22                            : out   std_logic;
          line_5_24                            : out   std_logic;
          line_5_25                            : out   std_logic;
          line_5_26                            : out   std_logic;
          line_5_27                            : out   std_logic;
          line_5_29                            : out   std_logic;
          line_5_30                            : out   std_logic;
          line_6_1                             : out   std_logic;
          line_6_2                             : out   std_logic;
          line_6_3                             : out   std_logic;
          line_6_4                             : out   std_logic;
          line_6_6                             : out   std_logic;
          line_6_7                             : out   std_logic;
          line_6_9                             : out   std_logic;
          line_6_10                            : out   std_logic;
          line_6_11                            : out   std_logic;
          line_6_14                            : out   std_logic;
          line_6_15                            : out   std_logic;
          line_6_16                            : out   std_logic;
          line_6_17                            : out   std_logic;
          line_6_18                            : out   std_logic;
          line_6_19                            : out   std_logic;
          line_6_20                            : out   std_logic;
          line_6_21                            : out   std_logic;
          line_6_22                            : out   std_logic;
          line_6_24                            : out   std_logic;
          line_6_25                            : out   std_logic;
          line_6_26                            : out   std_logic;
          line_6_27                            : out   std_logic;
          line_6_28                            : out   std_logic;
          line_6_29                            : out   std_logic;
          line_6_30                            : out   std_logic;
          line_6_31                            : out   std_logic;
          line_7_1                             : out   std_logic;
          line_7_2                             : out   std_logic;
          N_507                                : out   std_logic;
          N_508                                : out   std_logic;
          ren_pos                              : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          data_out_ready                       : in    std_logic := 'U';
          AHB_slave_dummy_0_read_en            : in    std_logic := 'U';
          start_wen                            : in    std_logic := 'U';
          SHA256_Module_0_error_o              : in    std_logic := 'U';
          SHA256_Module_0_di_req_o             : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o           : in    std_logic := 'U'
        );
  end component;

  component reg1_highonly
    port( CertificationSystem_sb_0_GPIO_9_M2F     : in    std_logic := 'U';
          CertificationSystem_sb_0_GPIO_9_M2F_i_0 : out   std_logic;
          start_wen                               : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0    : in    std_logic := 'U';
          SHA256_BLOCK_0_start_o                  : in    std_logic := 'U'
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \SHA256_Module_0_do_valid_o\, start_wen, 
        SHA256_BLOCK_0_do_valid_o, 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, 
        SHA256_BLOCK_0_start_o, \SHA256_BLOCK_0_H0_o[0]\, 
        \SHA256_BLOCK_0_H0_o[1]\, \SHA256_BLOCK_0_H0_o[2]\, 
        \SHA256_BLOCK_0_H0_o[3]\, \SHA256_BLOCK_0_H0_o[4]\, 
        \SHA256_BLOCK_0_H0_o[5]\, \SHA256_BLOCK_0_H0_o[6]\, 
        \SHA256_BLOCK_0_H0_o[7]\, \SHA256_BLOCK_0_H0_o[8]\, 
        \SHA256_BLOCK_0_H0_o[9]\, \SHA256_BLOCK_0_H0_o[10]\, 
        \SHA256_BLOCK_0_H0_o[11]\, \SHA256_BLOCK_0_H0_o[12]\, 
        \SHA256_BLOCK_0_H0_o[13]\, \SHA256_BLOCK_0_H0_o[14]\, 
        \SHA256_BLOCK_0_H0_o[15]\, \SHA256_BLOCK_0_H0_o[16]\, 
        \SHA256_BLOCK_0_H0_o[17]\, \SHA256_BLOCK_0_H0_o[18]\, 
        \SHA256_BLOCK_0_H0_o[19]\, \SHA256_BLOCK_0_H0_o[20]\, 
        \SHA256_BLOCK_0_H0_o[21]\, \SHA256_BLOCK_0_H0_o[22]\, 
        \SHA256_BLOCK_0_H0_o[23]\, \SHA256_BLOCK_0_H0_o[24]\, 
        \SHA256_BLOCK_0_H0_o[25]\, \SHA256_BLOCK_0_H0_o[26]\, 
        \SHA256_BLOCK_0_H0_o[27]\, \SHA256_BLOCK_0_H0_o[28]\, 
        \SHA256_BLOCK_0_H0_o[29]\, \SHA256_BLOCK_0_H0_o[30]\, 
        \SHA256_BLOCK_0_H0_o[31]\, \SHA256_BLOCK_0_H1_o[0]\, 
        \SHA256_BLOCK_0_H1_o[1]\, \SHA256_BLOCK_0_H1_o[2]\, 
        \SHA256_BLOCK_0_H1_o[3]\, \SHA256_BLOCK_0_H1_o[4]\, 
        \SHA256_BLOCK_0_H1_o[5]\, \SHA256_BLOCK_0_H1_o[6]\, 
        \SHA256_BLOCK_0_H1_o[7]\, \SHA256_BLOCK_0_H1_o[8]\, 
        \SHA256_BLOCK_0_H1_o[9]\, \SHA256_BLOCK_0_H1_o[10]\, 
        \SHA256_BLOCK_0_H1_o[11]\, \SHA256_BLOCK_0_H1_o[12]\, 
        \SHA256_BLOCK_0_H1_o[13]\, \SHA256_BLOCK_0_H1_o[14]\, 
        \SHA256_BLOCK_0_H1_o[15]\, \SHA256_BLOCK_0_H1_o[16]\, 
        \SHA256_BLOCK_0_H1_o[17]\, \SHA256_BLOCK_0_H1_o[18]\, 
        \SHA256_BLOCK_0_H1_o[19]\, \SHA256_BLOCK_0_H1_o[20]\, 
        \SHA256_BLOCK_0_H1_o[21]\, \SHA256_BLOCK_0_H1_o[22]\, 
        \SHA256_BLOCK_0_H1_o[23]\, \SHA256_BLOCK_0_H1_o[24]\, 
        \SHA256_BLOCK_0_H1_o[25]\, \SHA256_BLOCK_0_H1_o[26]\, 
        \SHA256_BLOCK_0_H1_o[27]\, \SHA256_BLOCK_0_H1_o[28]\, 
        \SHA256_BLOCK_0_H1_o[29]\, \SHA256_BLOCK_0_H1_o[30]\, 
        \SHA256_BLOCK_0_H1_o[31]\, \SHA256_BLOCK_0_H2_o[0]\, 
        \SHA256_BLOCK_0_H2_o[1]\, \SHA256_BLOCK_0_H2_o[2]\, 
        \SHA256_BLOCK_0_H2_o[3]\, \SHA256_BLOCK_0_H2_o[4]\, 
        \SHA256_BLOCK_0_H2_o[5]\, \SHA256_BLOCK_0_H2_o[6]\, 
        \SHA256_BLOCK_0_H2_o[7]\, \SHA256_BLOCK_0_H2_o[8]\, 
        \SHA256_BLOCK_0_H2_o[9]\, \SHA256_BLOCK_0_H2_o[10]\, 
        \SHA256_BLOCK_0_H2_o[11]\, \SHA256_BLOCK_0_H2_o[12]\, 
        \SHA256_BLOCK_0_H2_o[13]\, \SHA256_BLOCK_0_H2_o[14]\, 
        \SHA256_BLOCK_0_H2_o[15]\, \SHA256_BLOCK_0_H2_o[16]\, 
        \SHA256_BLOCK_0_H2_o[17]\, \SHA256_BLOCK_0_H2_o[18]\, 
        \SHA256_BLOCK_0_H2_o[19]\, \SHA256_BLOCK_0_H2_o[20]\, 
        \SHA256_BLOCK_0_H2_o[21]\, \SHA256_BLOCK_0_H2_o[22]\, 
        \SHA256_BLOCK_0_H2_o[23]\, \SHA256_BLOCK_0_H2_o[24]\, 
        \SHA256_BLOCK_0_H2_o[25]\, \SHA256_BLOCK_0_H2_o[26]\, 
        \SHA256_BLOCK_0_H2_o[27]\, \SHA256_BLOCK_0_H2_o[28]\, 
        \SHA256_BLOCK_0_H2_o[29]\, \SHA256_BLOCK_0_H2_o[30]\, 
        \SHA256_BLOCK_0_H2_o[31]\, \SHA256_BLOCK_0_H3_o[0]\, 
        \SHA256_BLOCK_0_H3_o[1]\, \SHA256_BLOCK_0_H3_o[2]\, 
        \SHA256_BLOCK_0_H3_o[3]\, \SHA256_BLOCK_0_H3_o[4]\, 
        \SHA256_BLOCK_0_H3_o[5]\, \SHA256_BLOCK_0_H3_o[6]\, 
        \SHA256_BLOCK_0_H3_o[7]\, \SHA256_BLOCK_0_H3_o[8]\, 
        \SHA256_BLOCK_0_H3_o[9]\, \SHA256_BLOCK_0_H3_o[10]\, 
        \SHA256_BLOCK_0_H3_o[11]\, \SHA256_BLOCK_0_H3_o[12]\, 
        \SHA256_BLOCK_0_H3_o[13]\, \SHA256_BLOCK_0_H3_o[14]\, 
        \SHA256_BLOCK_0_H3_o[15]\, \SHA256_BLOCK_0_H3_o[16]\, 
        \SHA256_BLOCK_0_H3_o[17]\, \SHA256_BLOCK_0_H3_o[18]\, 
        \SHA256_BLOCK_0_H3_o[19]\, \SHA256_BLOCK_0_H3_o[20]\, 
        \SHA256_BLOCK_0_H3_o[21]\, \SHA256_BLOCK_0_H3_o[22]\, 
        \SHA256_BLOCK_0_H3_o[23]\, \SHA256_BLOCK_0_H3_o[24]\, 
        \SHA256_BLOCK_0_H3_o[25]\, \SHA256_BLOCK_0_H3_o[26]\, 
        \SHA256_BLOCK_0_H3_o[27]\, \SHA256_BLOCK_0_H3_o[28]\, 
        \SHA256_BLOCK_0_H3_o[29]\, \SHA256_BLOCK_0_H3_o[30]\, 
        \SHA256_BLOCK_0_H3_o[31]\, \SHA256_BLOCK_0_H4_o[0]\, 
        \SHA256_BLOCK_0_H4_o[1]\, \SHA256_BLOCK_0_H4_o[2]\, 
        \SHA256_BLOCK_0_H4_o[3]\, \SHA256_BLOCK_0_H4_o[4]\, 
        \SHA256_BLOCK_0_H4_o[5]\, \SHA256_BLOCK_0_H4_o[6]\, 
        \SHA256_BLOCK_0_H4_o[7]\, \SHA256_BLOCK_0_H4_o[8]\, 
        \SHA256_BLOCK_0_H4_o[9]\, \SHA256_BLOCK_0_H4_o[10]\, 
        \SHA256_BLOCK_0_H4_o[11]\, \SHA256_BLOCK_0_H4_o[12]\, 
        \SHA256_BLOCK_0_H4_o[13]\, \SHA256_BLOCK_0_H4_o[14]\, 
        \SHA256_BLOCK_0_H4_o[15]\, \SHA256_BLOCK_0_H4_o[16]\, 
        \SHA256_BLOCK_0_H4_o[17]\, \SHA256_BLOCK_0_H4_o[18]\, 
        \SHA256_BLOCK_0_H4_o[19]\, \SHA256_BLOCK_0_H4_o[20]\, 
        \SHA256_BLOCK_0_H4_o[21]\, \SHA256_BLOCK_0_H4_o[22]\, 
        \SHA256_BLOCK_0_H4_o[23]\, \SHA256_BLOCK_0_H4_o[24]\, 
        \SHA256_BLOCK_0_H4_o[25]\, \SHA256_BLOCK_0_H4_o[26]\, 
        \SHA256_BLOCK_0_H4_o[27]\, \SHA256_BLOCK_0_H4_o[28]\, 
        \SHA256_BLOCK_0_H4_o[29]\, \SHA256_BLOCK_0_H4_o[30]\, 
        \SHA256_BLOCK_0_H4_o[31]\, \SHA256_BLOCK_0_H5_o[0]\, 
        \SHA256_BLOCK_0_H5_o[1]\, \SHA256_BLOCK_0_H5_o[2]\, 
        \SHA256_BLOCK_0_H5_o[3]\, \SHA256_BLOCK_0_H5_o[4]\, 
        \SHA256_BLOCK_0_H5_o[5]\, \SHA256_BLOCK_0_H5_o[6]\, 
        \SHA256_BLOCK_0_H5_o[7]\, \SHA256_BLOCK_0_H5_o[8]\, 
        \SHA256_BLOCK_0_H5_o[9]\, \SHA256_BLOCK_0_H5_o[10]\, 
        \SHA256_BLOCK_0_H5_o[11]\, \SHA256_BLOCK_0_H5_o[12]\, 
        \SHA256_BLOCK_0_H5_o[13]\, \SHA256_BLOCK_0_H5_o[14]\, 
        \SHA256_BLOCK_0_H5_o[15]\, \SHA256_BLOCK_0_H5_o[16]\, 
        \SHA256_BLOCK_0_H5_o[17]\, \SHA256_BLOCK_0_H5_o[18]\, 
        \SHA256_BLOCK_0_H5_o[19]\, \SHA256_BLOCK_0_H5_o[20]\, 
        \SHA256_BLOCK_0_H5_o[21]\, \SHA256_BLOCK_0_H5_o[22]\, 
        \SHA256_BLOCK_0_H5_o[23]\, \SHA256_BLOCK_0_H5_o[24]\, 
        \SHA256_BLOCK_0_H5_o[25]\, \SHA256_BLOCK_0_H5_o[26]\, 
        \SHA256_BLOCK_0_H5_o[27]\, \SHA256_BLOCK_0_H5_o[28]\, 
        \SHA256_BLOCK_0_H5_o[29]\, \SHA256_BLOCK_0_H5_o[30]\, 
        \SHA256_BLOCK_0_H5_o[31]\, \SHA256_BLOCK_0_H6_o[0]\, 
        \SHA256_BLOCK_0_H6_o[1]\, \SHA256_BLOCK_0_H6_o[2]\, 
        \SHA256_BLOCK_0_H6_o[3]\, \SHA256_BLOCK_0_H6_o[4]\, 
        \SHA256_BLOCK_0_H6_o[5]\, \SHA256_BLOCK_0_H6_o[6]\, 
        \SHA256_BLOCK_0_H6_o[7]\, \SHA256_BLOCK_0_H6_o[8]\, 
        \SHA256_BLOCK_0_H6_o[9]\, \SHA256_BLOCK_0_H6_o[10]\, 
        \SHA256_BLOCK_0_H6_o[11]\, \SHA256_BLOCK_0_H6_o[12]\, 
        \SHA256_BLOCK_0_H6_o[13]\, \SHA256_BLOCK_0_H6_o[14]\, 
        \SHA256_BLOCK_0_H6_o[15]\, \SHA256_BLOCK_0_H6_o[16]\, 
        \SHA256_BLOCK_0_H6_o[17]\, \SHA256_BLOCK_0_H6_o[18]\, 
        \SHA256_BLOCK_0_H6_o[19]\, \SHA256_BLOCK_0_H6_o[20]\, 
        \SHA256_BLOCK_0_H6_o[21]\, \SHA256_BLOCK_0_H6_o[22]\, 
        \SHA256_BLOCK_0_H6_o[23]\, \SHA256_BLOCK_0_H6_o[24]\, 
        \SHA256_BLOCK_0_H6_o[25]\, \SHA256_BLOCK_0_H6_o[26]\, 
        \SHA256_BLOCK_0_H6_o[27]\, \SHA256_BLOCK_0_H6_o[28]\, 
        \SHA256_BLOCK_0_H6_o[29]\, \SHA256_BLOCK_0_H6_o[30]\, 
        \SHA256_BLOCK_0_H6_o[31]\, \SHA256_BLOCK_0_H7_o[0]\, 
        \SHA256_BLOCK_0_H7_o[1]\, \SHA256_BLOCK_0_H7_o[2]\, 
        \SHA256_BLOCK_0_H7_o[3]\, \SHA256_BLOCK_0_H7_o[4]\, 
        \SHA256_BLOCK_0_H7_o[5]\, \SHA256_BLOCK_0_H7_o[6]\, 
        \SHA256_BLOCK_0_H7_o[7]\, \SHA256_BLOCK_0_H7_o[8]\, 
        \SHA256_BLOCK_0_H7_o[9]\, \SHA256_BLOCK_0_H7_o[10]\, 
        \SHA256_BLOCK_0_H7_o[11]\, \SHA256_BLOCK_0_H7_o[12]\, 
        \SHA256_BLOCK_0_H7_o[13]\, \SHA256_BLOCK_0_H7_o[14]\, 
        \SHA256_BLOCK_0_H7_o[15]\, \SHA256_BLOCK_0_H7_o[16]\, 
        \SHA256_BLOCK_0_H7_o[17]\, \SHA256_BLOCK_0_H7_o[18]\, 
        \SHA256_BLOCK_0_H7_o[19]\, \SHA256_BLOCK_0_H7_o[20]\, 
        \SHA256_BLOCK_0_H7_o[21]\, \SHA256_BLOCK_0_H7_o[22]\, 
        \SHA256_BLOCK_0_H7_o[23]\, \SHA256_BLOCK_0_H7_o[24]\, 
        \SHA256_BLOCK_0_H7_o[25]\, \SHA256_BLOCK_0_H7_o[26]\, 
        \SHA256_BLOCK_0_H7_o[27]\, \SHA256_BLOCK_0_H7_o[28]\, 
        \SHA256_BLOCK_0_H7_o[29]\, \SHA256_BLOCK_0_H7_o[30]\, 
        \SHA256_BLOCK_0_H7_o[31]\, data_out_ready, 
        \SHA256_Module_0_error_o\, \SHA256_Module_0_di_req_o\, 
        GND_net_1, VCC_net_1 : std_logic;

    for all : SHA256_BLOCK
	Use entity work.SHA256_BLOCK(DEF_ARCH);
    for all : reg9_1x32
	Use entity work.reg9_1x32(DEF_ARCH);
    for all : reg1_highonly
	Use entity work.reg1_highonly(DEF_ARCH);
begin 

    SHA256_Module_0_do_valid_o <= \SHA256_Module_0_do_valid_o\;
    SHA256_Module_0_error_o <= \SHA256_Module_0_error_o\;
    SHA256_Module_0_di_req_o <= \SHA256_Module_0_di_req_o\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    SHA256_BLOCK_0 : SHA256_BLOCK
      port map(SHA256_BLOCK_0_H0_o(31) => 
        \SHA256_BLOCK_0_H0_o[31]\, SHA256_BLOCK_0_H0_o(30) => 
        \SHA256_BLOCK_0_H0_o[30]\, SHA256_BLOCK_0_H0_o(29) => 
        \SHA256_BLOCK_0_H0_o[29]\, SHA256_BLOCK_0_H0_o(28) => 
        \SHA256_BLOCK_0_H0_o[28]\, SHA256_BLOCK_0_H0_o(27) => 
        \SHA256_BLOCK_0_H0_o[27]\, SHA256_BLOCK_0_H0_o(26) => 
        \SHA256_BLOCK_0_H0_o[26]\, SHA256_BLOCK_0_H0_o(25) => 
        \SHA256_BLOCK_0_H0_o[25]\, SHA256_BLOCK_0_H0_o(24) => 
        \SHA256_BLOCK_0_H0_o[24]\, SHA256_BLOCK_0_H0_o(23) => 
        \SHA256_BLOCK_0_H0_o[23]\, SHA256_BLOCK_0_H0_o(22) => 
        \SHA256_BLOCK_0_H0_o[22]\, SHA256_BLOCK_0_H0_o(21) => 
        \SHA256_BLOCK_0_H0_o[21]\, SHA256_BLOCK_0_H0_o(20) => 
        \SHA256_BLOCK_0_H0_o[20]\, SHA256_BLOCK_0_H0_o(19) => 
        \SHA256_BLOCK_0_H0_o[19]\, SHA256_BLOCK_0_H0_o(18) => 
        \SHA256_BLOCK_0_H0_o[18]\, SHA256_BLOCK_0_H0_o(17) => 
        \SHA256_BLOCK_0_H0_o[17]\, SHA256_BLOCK_0_H0_o(16) => 
        \SHA256_BLOCK_0_H0_o[16]\, SHA256_BLOCK_0_H0_o(15) => 
        \SHA256_BLOCK_0_H0_o[15]\, SHA256_BLOCK_0_H0_o(14) => 
        \SHA256_BLOCK_0_H0_o[14]\, SHA256_BLOCK_0_H0_o(13) => 
        \SHA256_BLOCK_0_H0_o[13]\, SHA256_BLOCK_0_H0_o(12) => 
        \SHA256_BLOCK_0_H0_o[12]\, SHA256_BLOCK_0_H0_o(11) => 
        \SHA256_BLOCK_0_H0_o[11]\, SHA256_BLOCK_0_H0_o(10) => 
        \SHA256_BLOCK_0_H0_o[10]\, SHA256_BLOCK_0_H0_o(9) => 
        \SHA256_BLOCK_0_H0_o[9]\, SHA256_BLOCK_0_H0_o(8) => 
        \SHA256_BLOCK_0_H0_o[8]\, SHA256_BLOCK_0_H0_o(7) => 
        \SHA256_BLOCK_0_H0_o[7]\, SHA256_BLOCK_0_H0_o(6) => 
        \SHA256_BLOCK_0_H0_o[6]\, SHA256_BLOCK_0_H0_o(5) => 
        \SHA256_BLOCK_0_H0_o[5]\, SHA256_BLOCK_0_H0_o(4) => 
        \SHA256_BLOCK_0_H0_o[4]\, SHA256_BLOCK_0_H0_o(3) => 
        \SHA256_BLOCK_0_H0_o[3]\, SHA256_BLOCK_0_H0_o(2) => 
        \SHA256_BLOCK_0_H0_o[2]\, SHA256_BLOCK_0_H0_o(1) => 
        \SHA256_BLOCK_0_H0_o[1]\, SHA256_BLOCK_0_H0_o(0) => 
        \SHA256_BLOCK_0_H0_o[0]\, SHA256_BLOCK_0_H1_o(31) => 
        \SHA256_BLOCK_0_H1_o[31]\, SHA256_BLOCK_0_H1_o(30) => 
        \SHA256_BLOCK_0_H1_o[30]\, SHA256_BLOCK_0_H1_o(29) => 
        \SHA256_BLOCK_0_H1_o[29]\, SHA256_BLOCK_0_H1_o(28) => 
        \SHA256_BLOCK_0_H1_o[28]\, SHA256_BLOCK_0_H1_o(27) => 
        \SHA256_BLOCK_0_H1_o[27]\, SHA256_BLOCK_0_H1_o(26) => 
        \SHA256_BLOCK_0_H1_o[26]\, SHA256_BLOCK_0_H1_o(25) => 
        \SHA256_BLOCK_0_H1_o[25]\, SHA256_BLOCK_0_H1_o(24) => 
        \SHA256_BLOCK_0_H1_o[24]\, SHA256_BLOCK_0_H1_o(23) => 
        \SHA256_BLOCK_0_H1_o[23]\, SHA256_BLOCK_0_H1_o(22) => 
        \SHA256_BLOCK_0_H1_o[22]\, SHA256_BLOCK_0_H1_o(21) => 
        \SHA256_BLOCK_0_H1_o[21]\, SHA256_BLOCK_0_H1_o(20) => 
        \SHA256_BLOCK_0_H1_o[20]\, SHA256_BLOCK_0_H1_o(19) => 
        \SHA256_BLOCK_0_H1_o[19]\, SHA256_BLOCK_0_H1_o(18) => 
        \SHA256_BLOCK_0_H1_o[18]\, SHA256_BLOCK_0_H1_o(17) => 
        \SHA256_BLOCK_0_H1_o[17]\, SHA256_BLOCK_0_H1_o(16) => 
        \SHA256_BLOCK_0_H1_o[16]\, SHA256_BLOCK_0_H1_o(15) => 
        \SHA256_BLOCK_0_H1_o[15]\, SHA256_BLOCK_0_H1_o(14) => 
        \SHA256_BLOCK_0_H1_o[14]\, SHA256_BLOCK_0_H1_o(13) => 
        \SHA256_BLOCK_0_H1_o[13]\, SHA256_BLOCK_0_H1_o(12) => 
        \SHA256_BLOCK_0_H1_o[12]\, SHA256_BLOCK_0_H1_o(11) => 
        \SHA256_BLOCK_0_H1_o[11]\, SHA256_BLOCK_0_H1_o(10) => 
        \SHA256_BLOCK_0_H1_o[10]\, SHA256_BLOCK_0_H1_o(9) => 
        \SHA256_BLOCK_0_H1_o[9]\, SHA256_BLOCK_0_H1_o(8) => 
        \SHA256_BLOCK_0_H1_o[8]\, SHA256_BLOCK_0_H1_o(7) => 
        \SHA256_BLOCK_0_H1_o[7]\, SHA256_BLOCK_0_H1_o(6) => 
        \SHA256_BLOCK_0_H1_o[6]\, SHA256_BLOCK_0_H1_o(5) => 
        \SHA256_BLOCK_0_H1_o[5]\, SHA256_BLOCK_0_H1_o(4) => 
        \SHA256_BLOCK_0_H1_o[4]\, SHA256_BLOCK_0_H1_o(3) => 
        \SHA256_BLOCK_0_H1_o[3]\, SHA256_BLOCK_0_H1_o(2) => 
        \SHA256_BLOCK_0_H1_o[2]\, SHA256_BLOCK_0_H1_o(1) => 
        \SHA256_BLOCK_0_H1_o[1]\, SHA256_BLOCK_0_H1_o(0) => 
        \SHA256_BLOCK_0_H1_o[0]\, SHA256_BLOCK_0_H2_o(31) => 
        \SHA256_BLOCK_0_H2_o[31]\, SHA256_BLOCK_0_H2_o(30) => 
        \SHA256_BLOCK_0_H2_o[30]\, SHA256_BLOCK_0_H2_o(29) => 
        \SHA256_BLOCK_0_H2_o[29]\, SHA256_BLOCK_0_H2_o(28) => 
        \SHA256_BLOCK_0_H2_o[28]\, SHA256_BLOCK_0_H2_o(27) => 
        \SHA256_BLOCK_0_H2_o[27]\, SHA256_BLOCK_0_H2_o(26) => 
        \SHA256_BLOCK_0_H2_o[26]\, SHA256_BLOCK_0_H2_o(25) => 
        \SHA256_BLOCK_0_H2_o[25]\, SHA256_BLOCK_0_H2_o(24) => 
        \SHA256_BLOCK_0_H2_o[24]\, SHA256_BLOCK_0_H2_o(23) => 
        \SHA256_BLOCK_0_H2_o[23]\, SHA256_BLOCK_0_H2_o(22) => 
        \SHA256_BLOCK_0_H2_o[22]\, SHA256_BLOCK_0_H2_o(21) => 
        \SHA256_BLOCK_0_H2_o[21]\, SHA256_BLOCK_0_H2_o(20) => 
        \SHA256_BLOCK_0_H2_o[20]\, SHA256_BLOCK_0_H2_o(19) => 
        \SHA256_BLOCK_0_H2_o[19]\, SHA256_BLOCK_0_H2_o(18) => 
        \SHA256_BLOCK_0_H2_o[18]\, SHA256_BLOCK_0_H2_o(17) => 
        \SHA256_BLOCK_0_H2_o[17]\, SHA256_BLOCK_0_H2_o(16) => 
        \SHA256_BLOCK_0_H2_o[16]\, SHA256_BLOCK_0_H2_o(15) => 
        \SHA256_BLOCK_0_H2_o[15]\, SHA256_BLOCK_0_H2_o(14) => 
        \SHA256_BLOCK_0_H2_o[14]\, SHA256_BLOCK_0_H2_o(13) => 
        \SHA256_BLOCK_0_H2_o[13]\, SHA256_BLOCK_0_H2_o(12) => 
        \SHA256_BLOCK_0_H2_o[12]\, SHA256_BLOCK_0_H2_o(11) => 
        \SHA256_BLOCK_0_H2_o[11]\, SHA256_BLOCK_0_H2_o(10) => 
        \SHA256_BLOCK_0_H2_o[10]\, SHA256_BLOCK_0_H2_o(9) => 
        \SHA256_BLOCK_0_H2_o[9]\, SHA256_BLOCK_0_H2_o(8) => 
        \SHA256_BLOCK_0_H2_o[8]\, SHA256_BLOCK_0_H2_o(7) => 
        \SHA256_BLOCK_0_H2_o[7]\, SHA256_BLOCK_0_H2_o(6) => 
        \SHA256_BLOCK_0_H2_o[6]\, SHA256_BLOCK_0_H2_o(5) => 
        \SHA256_BLOCK_0_H2_o[5]\, SHA256_BLOCK_0_H2_o(4) => 
        \SHA256_BLOCK_0_H2_o[4]\, SHA256_BLOCK_0_H2_o(3) => 
        \SHA256_BLOCK_0_H2_o[3]\, SHA256_BLOCK_0_H2_o(2) => 
        \SHA256_BLOCK_0_H2_o[2]\, SHA256_BLOCK_0_H2_o(1) => 
        \SHA256_BLOCK_0_H2_o[1]\, SHA256_BLOCK_0_H2_o(0) => 
        \SHA256_BLOCK_0_H2_o[0]\, SHA256_BLOCK_0_H3_o(31) => 
        \SHA256_BLOCK_0_H3_o[31]\, SHA256_BLOCK_0_H3_o(30) => 
        \SHA256_BLOCK_0_H3_o[30]\, SHA256_BLOCK_0_H3_o(29) => 
        \SHA256_BLOCK_0_H3_o[29]\, SHA256_BLOCK_0_H3_o(28) => 
        \SHA256_BLOCK_0_H3_o[28]\, SHA256_BLOCK_0_H3_o(27) => 
        \SHA256_BLOCK_0_H3_o[27]\, SHA256_BLOCK_0_H3_o(26) => 
        \SHA256_BLOCK_0_H3_o[26]\, SHA256_BLOCK_0_H3_o(25) => 
        \SHA256_BLOCK_0_H3_o[25]\, SHA256_BLOCK_0_H3_o(24) => 
        \SHA256_BLOCK_0_H3_o[24]\, SHA256_BLOCK_0_H3_o(23) => 
        \SHA256_BLOCK_0_H3_o[23]\, SHA256_BLOCK_0_H3_o(22) => 
        \SHA256_BLOCK_0_H3_o[22]\, SHA256_BLOCK_0_H3_o(21) => 
        \SHA256_BLOCK_0_H3_o[21]\, SHA256_BLOCK_0_H3_o(20) => 
        \SHA256_BLOCK_0_H3_o[20]\, SHA256_BLOCK_0_H3_o(19) => 
        \SHA256_BLOCK_0_H3_o[19]\, SHA256_BLOCK_0_H3_o(18) => 
        \SHA256_BLOCK_0_H3_o[18]\, SHA256_BLOCK_0_H3_o(17) => 
        \SHA256_BLOCK_0_H3_o[17]\, SHA256_BLOCK_0_H3_o(16) => 
        \SHA256_BLOCK_0_H3_o[16]\, SHA256_BLOCK_0_H3_o(15) => 
        \SHA256_BLOCK_0_H3_o[15]\, SHA256_BLOCK_0_H3_o(14) => 
        \SHA256_BLOCK_0_H3_o[14]\, SHA256_BLOCK_0_H3_o(13) => 
        \SHA256_BLOCK_0_H3_o[13]\, SHA256_BLOCK_0_H3_o(12) => 
        \SHA256_BLOCK_0_H3_o[12]\, SHA256_BLOCK_0_H3_o(11) => 
        \SHA256_BLOCK_0_H3_o[11]\, SHA256_BLOCK_0_H3_o(10) => 
        \SHA256_BLOCK_0_H3_o[10]\, SHA256_BLOCK_0_H3_o(9) => 
        \SHA256_BLOCK_0_H3_o[9]\, SHA256_BLOCK_0_H3_o(8) => 
        \SHA256_BLOCK_0_H3_o[8]\, SHA256_BLOCK_0_H3_o(7) => 
        \SHA256_BLOCK_0_H3_o[7]\, SHA256_BLOCK_0_H3_o(6) => 
        \SHA256_BLOCK_0_H3_o[6]\, SHA256_BLOCK_0_H3_o(5) => 
        \SHA256_BLOCK_0_H3_o[5]\, SHA256_BLOCK_0_H3_o(4) => 
        \SHA256_BLOCK_0_H3_o[4]\, SHA256_BLOCK_0_H3_o(3) => 
        \SHA256_BLOCK_0_H3_o[3]\, SHA256_BLOCK_0_H3_o(2) => 
        \SHA256_BLOCK_0_H3_o[2]\, SHA256_BLOCK_0_H3_o(1) => 
        \SHA256_BLOCK_0_H3_o[1]\, SHA256_BLOCK_0_H3_o(0) => 
        \SHA256_BLOCK_0_H3_o[0]\, SHA256_BLOCK_0_H4_o(31) => 
        \SHA256_BLOCK_0_H4_o[31]\, SHA256_BLOCK_0_H4_o(30) => 
        \SHA256_BLOCK_0_H4_o[30]\, SHA256_BLOCK_0_H4_o(29) => 
        \SHA256_BLOCK_0_H4_o[29]\, SHA256_BLOCK_0_H4_o(28) => 
        \SHA256_BLOCK_0_H4_o[28]\, SHA256_BLOCK_0_H4_o(27) => 
        \SHA256_BLOCK_0_H4_o[27]\, SHA256_BLOCK_0_H4_o(26) => 
        \SHA256_BLOCK_0_H4_o[26]\, SHA256_BLOCK_0_H4_o(25) => 
        \SHA256_BLOCK_0_H4_o[25]\, SHA256_BLOCK_0_H4_o(24) => 
        \SHA256_BLOCK_0_H4_o[24]\, SHA256_BLOCK_0_H4_o(23) => 
        \SHA256_BLOCK_0_H4_o[23]\, SHA256_BLOCK_0_H4_o(22) => 
        \SHA256_BLOCK_0_H4_o[22]\, SHA256_BLOCK_0_H4_o(21) => 
        \SHA256_BLOCK_0_H4_o[21]\, SHA256_BLOCK_0_H4_o(20) => 
        \SHA256_BLOCK_0_H4_o[20]\, SHA256_BLOCK_0_H4_o(19) => 
        \SHA256_BLOCK_0_H4_o[19]\, SHA256_BLOCK_0_H4_o(18) => 
        \SHA256_BLOCK_0_H4_o[18]\, SHA256_BLOCK_0_H4_o(17) => 
        \SHA256_BLOCK_0_H4_o[17]\, SHA256_BLOCK_0_H4_o(16) => 
        \SHA256_BLOCK_0_H4_o[16]\, SHA256_BLOCK_0_H4_o(15) => 
        \SHA256_BLOCK_0_H4_o[15]\, SHA256_BLOCK_0_H4_o(14) => 
        \SHA256_BLOCK_0_H4_o[14]\, SHA256_BLOCK_0_H4_o(13) => 
        \SHA256_BLOCK_0_H4_o[13]\, SHA256_BLOCK_0_H4_o(12) => 
        \SHA256_BLOCK_0_H4_o[12]\, SHA256_BLOCK_0_H4_o(11) => 
        \SHA256_BLOCK_0_H4_o[11]\, SHA256_BLOCK_0_H4_o(10) => 
        \SHA256_BLOCK_0_H4_o[10]\, SHA256_BLOCK_0_H4_o(9) => 
        \SHA256_BLOCK_0_H4_o[9]\, SHA256_BLOCK_0_H4_o(8) => 
        \SHA256_BLOCK_0_H4_o[8]\, SHA256_BLOCK_0_H4_o(7) => 
        \SHA256_BLOCK_0_H4_o[7]\, SHA256_BLOCK_0_H4_o(6) => 
        \SHA256_BLOCK_0_H4_o[6]\, SHA256_BLOCK_0_H4_o(5) => 
        \SHA256_BLOCK_0_H4_o[5]\, SHA256_BLOCK_0_H4_o(4) => 
        \SHA256_BLOCK_0_H4_o[4]\, SHA256_BLOCK_0_H4_o(3) => 
        \SHA256_BLOCK_0_H4_o[3]\, SHA256_BLOCK_0_H4_o(2) => 
        \SHA256_BLOCK_0_H4_o[2]\, SHA256_BLOCK_0_H4_o(1) => 
        \SHA256_BLOCK_0_H4_o[1]\, SHA256_BLOCK_0_H4_o(0) => 
        \SHA256_BLOCK_0_H4_o[0]\, SHA256_BLOCK_0_H5_o(31) => 
        \SHA256_BLOCK_0_H5_o[31]\, SHA256_BLOCK_0_H5_o(30) => 
        \SHA256_BLOCK_0_H5_o[30]\, SHA256_BLOCK_0_H5_o(29) => 
        \SHA256_BLOCK_0_H5_o[29]\, SHA256_BLOCK_0_H5_o(28) => 
        \SHA256_BLOCK_0_H5_o[28]\, SHA256_BLOCK_0_H5_o(27) => 
        \SHA256_BLOCK_0_H5_o[27]\, SHA256_BLOCK_0_H5_o(26) => 
        \SHA256_BLOCK_0_H5_o[26]\, SHA256_BLOCK_0_H5_o(25) => 
        \SHA256_BLOCK_0_H5_o[25]\, SHA256_BLOCK_0_H5_o(24) => 
        \SHA256_BLOCK_0_H5_o[24]\, SHA256_BLOCK_0_H5_o(23) => 
        \SHA256_BLOCK_0_H5_o[23]\, SHA256_BLOCK_0_H5_o(22) => 
        \SHA256_BLOCK_0_H5_o[22]\, SHA256_BLOCK_0_H5_o(21) => 
        \SHA256_BLOCK_0_H5_o[21]\, SHA256_BLOCK_0_H5_o(20) => 
        \SHA256_BLOCK_0_H5_o[20]\, SHA256_BLOCK_0_H5_o(19) => 
        \SHA256_BLOCK_0_H5_o[19]\, SHA256_BLOCK_0_H5_o(18) => 
        \SHA256_BLOCK_0_H5_o[18]\, SHA256_BLOCK_0_H5_o(17) => 
        \SHA256_BLOCK_0_H5_o[17]\, SHA256_BLOCK_0_H5_o(16) => 
        \SHA256_BLOCK_0_H5_o[16]\, SHA256_BLOCK_0_H5_o(15) => 
        \SHA256_BLOCK_0_H5_o[15]\, SHA256_BLOCK_0_H5_o(14) => 
        \SHA256_BLOCK_0_H5_o[14]\, SHA256_BLOCK_0_H5_o(13) => 
        \SHA256_BLOCK_0_H5_o[13]\, SHA256_BLOCK_0_H5_o(12) => 
        \SHA256_BLOCK_0_H5_o[12]\, SHA256_BLOCK_0_H5_o(11) => 
        \SHA256_BLOCK_0_H5_o[11]\, SHA256_BLOCK_0_H5_o(10) => 
        \SHA256_BLOCK_0_H5_o[10]\, SHA256_BLOCK_0_H5_o(9) => 
        \SHA256_BLOCK_0_H5_o[9]\, SHA256_BLOCK_0_H5_o(8) => 
        \SHA256_BLOCK_0_H5_o[8]\, SHA256_BLOCK_0_H5_o(7) => 
        \SHA256_BLOCK_0_H5_o[7]\, SHA256_BLOCK_0_H5_o(6) => 
        \SHA256_BLOCK_0_H5_o[6]\, SHA256_BLOCK_0_H5_o(5) => 
        \SHA256_BLOCK_0_H5_o[5]\, SHA256_BLOCK_0_H5_o(4) => 
        \SHA256_BLOCK_0_H5_o[4]\, SHA256_BLOCK_0_H5_o(3) => 
        \SHA256_BLOCK_0_H5_o[3]\, SHA256_BLOCK_0_H5_o(2) => 
        \SHA256_BLOCK_0_H5_o[2]\, SHA256_BLOCK_0_H5_o(1) => 
        \SHA256_BLOCK_0_H5_o[1]\, SHA256_BLOCK_0_H5_o(0) => 
        \SHA256_BLOCK_0_H5_o[0]\, SHA256_BLOCK_0_H6_o(31) => 
        \SHA256_BLOCK_0_H6_o[31]\, SHA256_BLOCK_0_H6_o(30) => 
        \SHA256_BLOCK_0_H6_o[30]\, SHA256_BLOCK_0_H6_o(29) => 
        \SHA256_BLOCK_0_H6_o[29]\, SHA256_BLOCK_0_H6_o(28) => 
        \SHA256_BLOCK_0_H6_o[28]\, SHA256_BLOCK_0_H6_o(27) => 
        \SHA256_BLOCK_0_H6_o[27]\, SHA256_BLOCK_0_H6_o(26) => 
        \SHA256_BLOCK_0_H6_o[26]\, SHA256_BLOCK_0_H6_o(25) => 
        \SHA256_BLOCK_0_H6_o[25]\, SHA256_BLOCK_0_H6_o(24) => 
        \SHA256_BLOCK_0_H6_o[24]\, SHA256_BLOCK_0_H6_o(23) => 
        \SHA256_BLOCK_0_H6_o[23]\, SHA256_BLOCK_0_H6_o(22) => 
        \SHA256_BLOCK_0_H6_o[22]\, SHA256_BLOCK_0_H6_o(21) => 
        \SHA256_BLOCK_0_H6_o[21]\, SHA256_BLOCK_0_H6_o(20) => 
        \SHA256_BLOCK_0_H6_o[20]\, SHA256_BLOCK_0_H6_o(19) => 
        \SHA256_BLOCK_0_H6_o[19]\, SHA256_BLOCK_0_H6_o(18) => 
        \SHA256_BLOCK_0_H6_o[18]\, SHA256_BLOCK_0_H6_o(17) => 
        \SHA256_BLOCK_0_H6_o[17]\, SHA256_BLOCK_0_H6_o(16) => 
        \SHA256_BLOCK_0_H6_o[16]\, SHA256_BLOCK_0_H6_o(15) => 
        \SHA256_BLOCK_0_H6_o[15]\, SHA256_BLOCK_0_H6_o(14) => 
        \SHA256_BLOCK_0_H6_o[14]\, SHA256_BLOCK_0_H6_o(13) => 
        \SHA256_BLOCK_0_H6_o[13]\, SHA256_BLOCK_0_H6_o(12) => 
        \SHA256_BLOCK_0_H6_o[12]\, SHA256_BLOCK_0_H6_o(11) => 
        \SHA256_BLOCK_0_H6_o[11]\, SHA256_BLOCK_0_H6_o(10) => 
        \SHA256_BLOCK_0_H6_o[10]\, SHA256_BLOCK_0_H6_o(9) => 
        \SHA256_BLOCK_0_H6_o[9]\, SHA256_BLOCK_0_H6_o(8) => 
        \SHA256_BLOCK_0_H6_o[8]\, SHA256_BLOCK_0_H6_o(7) => 
        \SHA256_BLOCK_0_H6_o[7]\, SHA256_BLOCK_0_H6_o(6) => 
        \SHA256_BLOCK_0_H6_o[6]\, SHA256_BLOCK_0_H6_o(5) => 
        \SHA256_BLOCK_0_H6_o[5]\, SHA256_BLOCK_0_H6_o(4) => 
        \SHA256_BLOCK_0_H6_o[4]\, SHA256_BLOCK_0_H6_o(3) => 
        \SHA256_BLOCK_0_H6_o[3]\, SHA256_BLOCK_0_H6_o(2) => 
        \SHA256_BLOCK_0_H6_o[2]\, SHA256_BLOCK_0_H6_o(1) => 
        \SHA256_BLOCK_0_H6_o[1]\, SHA256_BLOCK_0_H6_o(0) => 
        \SHA256_BLOCK_0_H6_o[0]\, SHA256_BLOCK_0_H7_o(31) => 
        \SHA256_BLOCK_0_H7_o[31]\, SHA256_BLOCK_0_H7_o(30) => 
        \SHA256_BLOCK_0_H7_o[30]\, SHA256_BLOCK_0_H7_o(29) => 
        \SHA256_BLOCK_0_H7_o[29]\, SHA256_BLOCK_0_H7_o(28) => 
        \SHA256_BLOCK_0_H7_o[28]\, SHA256_BLOCK_0_H7_o(27) => 
        \SHA256_BLOCK_0_H7_o[27]\, SHA256_BLOCK_0_H7_o(26) => 
        \SHA256_BLOCK_0_H7_o[26]\, SHA256_BLOCK_0_H7_o(25) => 
        \SHA256_BLOCK_0_H7_o[25]\, SHA256_BLOCK_0_H7_o(24) => 
        \SHA256_BLOCK_0_H7_o[24]\, SHA256_BLOCK_0_H7_o(23) => 
        \SHA256_BLOCK_0_H7_o[23]\, SHA256_BLOCK_0_H7_o(22) => 
        \SHA256_BLOCK_0_H7_o[22]\, SHA256_BLOCK_0_H7_o(21) => 
        \SHA256_BLOCK_0_H7_o[21]\, SHA256_BLOCK_0_H7_o(20) => 
        \SHA256_BLOCK_0_H7_o[20]\, SHA256_BLOCK_0_H7_o(19) => 
        \SHA256_BLOCK_0_H7_o[19]\, SHA256_BLOCK_0_H7_o(18) => 
        \SHA256_BLOCK_0_H7_o[18]\, SHA256_BLOCK_0_H7_o(17) => 
        \SHA256_BLOCK_0_H7_o[17]\, SHA256_BLOCK_0_H7_o(16) => 
        \SHA256_BLOCK_0_H7_o[16]\, SHA256_BLOCK_0_H7_o(15) => 
        \SHA256_BLOCK_0_H7_o[15]\, SHA256_BLOCK_0_H7_o(14) => 
        \SHA256_BLOCK_0_H7_o[14]\, SHA256_BLOCK_0_H7_o(13) => 
        \SHA256_BLOCK_0_H7_o[13]\, SHA256_BLOCK_0_H7_o(12) => 
        \SHA256_BLOCK_0_H7_o[12]\, SHA256_BLOCK_0_H7_o(11) => 
        \SHA256_BLOCK_0_H7_o[11]\, SHA256_BLOCK_0_H7_o(10) => 
        \SHA256_BLOCK_0_H7_o[10]\, SHA256_BLOCK_0_H7_o(9) => 
        \SHA256_BLOCK_0_H7_o[9]\, SHA256_BLOCK_0_H7_o(8) => 
        \SHA256_BLOCK_0_H7_o[8]\, SHA256_BLOCK_0_H7_o(7) => 
        \SHA256_BLOCK_0_H7_o[7]\, SHA256_BLOCK_0_H7_o(6) => 
        \SHA256_BLOCK_0_H7_o[6]\, SHA256_BLOCK_0_H7_o(5) => 
        \SHA256_BLOCK_0_H7_o[5]\, SHA256_BLOCK_0_H7_o(4) => 
        \SHA256_BLOCK_0_H7_o[4]\, SHA256_BLOCK_0_H7_o(3) => 
        \SHA256_BLOCK_0_H7_o[3]\, SHA256_BLOCK_0_H7_o(2) => 
        \SHA256_BLOCK_0_H7_o[2]\, SHA256_BLOCK_0_H7_o(1) => 
        \SHA256_BLOCK_0_H7_o[1]\, SHA256_BLOCK_0_H7_o(0) => 
        \SHA256_BLOCK_0_H7_o[0]\, waddr_in_net_0(4) => 
        waddr_in_net_0(4), waddr_in_net_0(3) => waddr_in_net_0(3), 
        waddr_in_net_0(2) => waddr_in_net_0(2), waddr_in_net_0(1)
         => waddr_in_net_0(1), waddr_in_net_0(0) => 
        waddr_in_net_0(0), CertificationSystem_sb_0_FAB_CCC_GL0
         => CertificationSystem_sb_0_FAB_CCC_GL0, 
        SHA256_Module_0_di_req_o => \SHA256_Module_0_di_req_o\, 
        SHA256_BLOCK_0_do_valid_o => SHA256_BLOCK_0_do_valid_o, 
        SHA256_Module_0_waiting_data => 
        SHA256_Module_0_waiting_data, 
        SHA256_Module_0_data_available_lastbank_8 => 
        SHA256_Module_0_data_available_lastbank_8, 
        SHA256_Module_0_error_o => \SHA256_Module_0_error_o\, 
        SHA256_BLOCK_0_start_o => SHA256_BLOCK_0_start_o, 
        data_out_ready => data_out_ready, 
        CertificationSystem_sb_0_GPIO_9_M2F => 
        CertificationSystem_sb_0_GPIO_9_M2F, 
        SHA256_Module_0_data_available => 
        SHA256_Module_0_data_available, N_111_i_0 => N_111_i_0, 
        N_109_i_0 => N_109_i_0, N_168_i_0 => N_168_i_0, N_107_i_0
         => N_107_i_0, N_99_i_0 => N_99_i_0, N_97_i_0 => N_97_i_0, 
        N_67_i_0 => N_67_i_0, N_65_i_0 => N_65_i_0, 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0 => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, N_105_i_0 => 
        N_105_i_0, N_103_i_0 => N_103_i_0, N_158_i_0 => N_158_i_0, 
        N_156_i_0 => N_156_i_0, N_101_i_0 => N_101_i_0, N_152_i_0
         => N_152_i_0, N_95_i_0 => N_95_i_0, N_93_i_0 => N_93_i_0, 
        N_91_i_0 => N_91_i_0, N_140_i_0 => N_140_i_0, N_89_i_0
         => N_89_i_0, N_87_i_0 => N_87_i_0, N_133_i_0 => 
        N_133_i_0, N_85_i_0 => N_85_i_0, N_83_i_0 => N_83_i_0, 
        N_77_i_0 => N_77_i_0, N_75_i_0 => N_75_i_0, N_73_i_0 => 
        N_73_i_0, N_71_i_0 => N_71_i_0, N_69_i_0 => N_69_i_0, 
        N_116_i_0 => N_116_i_0, N_114_i_0 => N_114_i_0, N_112_i_0
         => N_112_i_0, N_110_i_0 => N_110_i_0, 
        CertificationSystem_sb_0_GPIO_1_M2F => 
        CertificationSystem_sb_0_GPIO_1_M2F, 
        AHB_slave_dummy_0_write_en => AHB_slave_dummy_0_write_en);
    
    reg9_1x32_0 : reg9_1x32
      port map(result_addr_net_0(3) => result_addr_net_0(3), 
        result_addr_net_0(2) => result_addr_net_0(2), 
        result_addr_net_0(1) => result_addr_net_0(1), 
        result_addr_net_0(0) => result_addr_net_0(0), 
        SHA256_BLOCK_0_H0_o(31) => \SHA256_BLOCK_0_H0_o[31]\, 
        SHA256_BLOCK_0_H0_o(30) => \SHA256_BLOCK_0_H0_o[30]\, 
        SHA256_BLOCK_0_H0_o(29) => \SHA256_BLOCK_0_H0_o[29]\, 
        SHA256_BLOCK_0_H0_o(28) => \SHA256_BLOCK_0_H0_o[28]\, 
        SHA256_BLOCK_0_H0_o(27) => \SHA256_BLOCK_0_H0_o[27]\, 
        SHA256_BLOCK_0_H0_o(26) => \SHA256_BLOCK_0_H0_o[26]\, 
        SHA256_BLOCK_0_H0_o(25) => \SHA256_BLOCK_0_H0_o[25]\, 
        SHA256_BLOCK_0_H0_o(24) => \SHA256_BLOCK_0_H0_o[24]\, 
        SHA256_BLOCK_0_H0_o(23) => \SHA256_BLOCK_0_H0_o[23]\, 
        SHA256_BLOCK_0_H0_o(22) => \SHA256_BLOCK_0_H0_o[22]\, 
        SHA256_BLOCK_0_H0_o(21) => \SHA256_BLOCK_0_H0_o[21]\, 
        SHA256_BLOCK_0_H0_o(20) => \SHA256_BLOCK_0_H0_o[20]\, 
        SHA256_BLOCK_0_H0_o(19) => \SHA256_BLOCK_0_H0_o[19]\, 
        SHA256_BLOCK_0_H0_o(18) => \SHA256_BLOCK_0_H0_o[18]\, 
        SHA256_BLOCK_0_H0_o(17) => \SHA256_BLOCK_0_H0_o[17]\, 
        SHA256_BLOCK_0_H0_o(16) => \SHA256_BLOCK_0_H0_o[16]\, 
        SHA256_BLOCK_0_H0_o(15) => \SHA256_BLOCK_0_H0_o[15]\, 
        SHA256_BLOCK_0_H0_o(14) => \SHA256_BLOCK_0_H0_o[14]\, 
        SHA256_BLOCK_0_H0_o(13) => \SHA256_BLOCK_0_H0_o[13]\, 
        SHA256_BLOCK_0_H0_o(12) => \SHA256_BLOCK_0_H0_o[12]\, 
        SHA256_BLOCK_0_H0_o(11) => \SHA256_BLOCK_0_H0_o[11]\, 
        SHA256_BLOCK_0_H0_o(10) => \SHA256_BLOCK_0_H0_o[10]\, 
        SHA256_BLOCK_0_H0_o(9) => \SHA256_BLOCK_0_H0_o[9]\, 
        SHA256_BLOCK_0_H0_o(8) => \SHA256_BLOCK_0_H0_o[8]\, 
        SHA256_BLOCK_0_H0_o(7) => \SHA256_BLOCK_0_H0_o[7]\, 
        SHA256_BLOCK_0_H0_o(6) => \SHA256_BLOCK_0_H0_o[6]\, 
        SHA256_BLOCK_0_H0_o(5) => \SHA256_BLOCK_0_H0_o[5]\, 
        SHA256_BLOCK_0_H0_o(4) => \SHA256_BLOCK_0_H0_o[4]\, 
        SHA256_BLOCK_0_H0_o(3) => \SHA256_BLOCK_0_H0_o[3]\, 
        SHA256_BLOCK_0_H0_o(2) => \SHA256_BLOCK_0_H0_o[2]\, 
        SHA256_BLOCK_0_H0_o(1) => \SHA256_BLOCK_0_H0_o[1]\, 
        SHA256_BLOCK_0_H0_o(0) => \SHA256_BLOCK_0_H0_o[0]\, 
        SHA256_BLOCK_0_H1_o(31) => \SHA256_BLOCK_0_H1_o[31]\, 
        SHA256_BLOCK_0_H1_o(30) => \SHA256_BLOCK_0_H1_o[30]\, 
        SHA256_BLOCK_0_H1_o(29) => \SHA256_BLOCK_0_H1_o[29]\, 
        SHA256_BLOCK_0_H1_o(28) => \SHA256_BLOCK_0_H1_o[28]\, 
        SHA256_BLOCK_0_H1_o(27) => \SHA256_BLOCK_0_H1_o[27]\, 
        SHA256_BLOCK_0_H1_o(26) => \SHA256_BLOCK_0_H1_o[26]\, 
        SHA256_BLOCK_0_H1_o(25) => \SHA256_BLOCK_0_H1_o[25]\, 
        SHA256_BLOCK_0_H1_o(24) => \SHA256_BLOCK_0_H1_o[24]\, 
        SHA256_BLOCK_0_H1_o(23) => \SHA256_BLOCK_0_H1_o[23]\, 
        SHA256_BLOCK_0_H1_o(22) => \SHA256_BLOCK_0_H1_o[22]\, 
        SHA256_BLOCK_0_H1_o(21) => \SHA256_BLOCK_0_H1_o[21]\, 
        SHA256_BLOCK_0_H1_o(20) => \SHA256_BLOCK_0_H1_o[20]\, 
        SHA256_BLOCK_0_H1_o(19) => \SHA256_BLOCK_0_H1_o[19]\, 
        SHA256_BLOCK_0_H1_o(18) => \SHA256_BLOCK_0_H1_o[18]\, 
        SHA256_BLOCK_0_H1_o(17) => \SHA256_BLOCK_0_H1_o[17]\, 
        SHA256_BLOCK_0_H1_o(16) => \SHA256_BLOCK_0_H1_o[16]\, 
        SHA256_BLOCK_0_H1_o(15) => \SHA256_BLOCK_0_H1_o[15]\, 
        SHA256_BLOCK_0_H1_o(14) => \SHA256_BLOCK_0_H1_o[14]\, 
        SHA256_BLOCK_0_H1_o(13) => \SHA256_BLOCK_0_H1_o[13]\, 
        SHA256_BLOCK_0_H1_o(12) => \SHA256_BLOCK_0_H1_o[12]\, 
        SHA256_BLOCK_0_H1_o(11) => \SHA256_BLOCK_0_H1_o[11]\, 
        SHA256_BLOCK_0_H1_o(10) => \SHA256_BLOCK_0_H1_o[10]\, 
        SHA256_BLOCK_0_H1_o(9) => \SHA256_BLOCK_0_H1_o[9]\, 
        SHA256_BLOCK_0_H1_o(8) => \SHA256_BLOCK_0_H1_o[8]\, 
        SHA256_BLOCK_0_H1_o(7) => \SHA256_BLOCK_0_H1_o[7]\, 
        SHA256_BLOCK_0_H1_o(6) => \SHA256_BLOCK_0_H1_o[6]\, 
        SHA256_BLOCK_0_H1_o(5) => \SHA256_BLOCK_0_H1_o[5]\, 
        SHA256_BLOCK_0_H1_o(4) => \SHA256_BLOCK_0_H1_o[4]\, 
        SHA256_BLOCK_0_H1_o(3) => \SHA256_BLOCK_0_H1_o[3]\, 
        SHA256_BLOCK_0_H1_o(2) => \SHA256_BLOCK_0_H1_o[2]\, 
        SHA256_BLOCK_0_H1_o(1) => \SHA256_BLOCK_0_H1_o[1]\, 
        SHA256_BLOCK_0_H1_o(0) => \SHA256_BLOCK_0_H1_o[0]\, 
        SHA256_BLOCK_0_H2_o(31) => \SHA256_BLOCK_0_H2_o[31]\, 
        SHA256_BLOCK_0_H2_o(30) => \SHA256_BLOCK_0_H2_o[30]\, 
        SHA256_BLOCK_0_H2_o(29) => \SHA256_BLOCK_0_H2_o[29]\, 
        SHA256_BLOCK_0_H2_o(28) => \SHA256_BLOCK_0_H2_o[28]\, 
        SHA256_BLOCK_0_H2_o(27) => \SHA256_BLOCK_0_H2_o[27]\, 
        SHA256_BLOCK_0_H2_o(26) => \SHA256_BLOCK_0_H2_o[26]\, 
        SHA256_BLOCK_0_H2_o(25) => \SHA256_BLOCK_0_H2_o[25]\, 
        SHA256_BLOCK_0_H2_o(24) => \SHA256_BLOCK_0_H2_o[24]\, 
        SHA256_BLOCK_0_H2_o(23) => \SHA256_BLOCK_0_H2_o[23]\, 
        SHA256_BLOCK_0_H2_o(22) => \SHA256_BLOCK_0_H2_o[22]\, 
        SHA256_BLOCK_0_H2_o(21) => \SHA256_BLOCK_0_H2_o[21]\, 
        SHA256_BLOCK_0_H2_o(20) => \SHA256_BLOCK_0_H2_o[20]\, 
        SHA256_BLOCK_0_H2_o(19) => \SHA256_BLOCK_0_H2_o[19]\, 
        SHA256_BLOCK_0_H2_o(18) => \SHA256_BLOCK_0_H2_o[18]\, 
        SHA256_BLOCK_0_H2_o(17) => \SHA256_BLOCK_0_H2_o[17]\, 
        SHA256_BLOCK_0_H2_o(16) => \SHA256_BLOCK_0_H2_o[16]\, 
        SHA256_BLOCK_0_H2_o(15) => \SHA256_BLOCK_0_H2_o[15]\, 
        SHA256_BLOCK_0_H2_o(14) => \SHA256_BLOCK_0_H2_o[14]\, 
        SHA256_BLOCK_0_H2_o(13) => \SHA256_BLOCK_0_H2_o[13]\, 
        SHA256_BLOCK_0_H2_o(12) => \SHA256_BLOCK_0_H2_o[12]\, 
        SHA256_BLOCK_0_H2_o(11) => \SHA256_BLOCK_0_H2_o[11]\, 
        SHA256_BLOCK_0_H2_o(10) => \SHA256_BLOCK_0_H2_o[10]\, 
        SHA256_BLOCK_0_H2_o(9) => \SHA256_BLOCK_0_H2_o[9]\, 
        SHA256_BLOCK_0_H2_o(8) => \SHA256_BLOCK_0_H2_o[8]\, 
        SHA256_BLOCK_0_H2_o(7) => \SHA256_BLOCK_0_H2_o[7]\, 
        SHA256_BLOCK_0_H2_o(6) => \SHA256_BLOCK_0_H2_o[6]\, 
        SHA256_BLOCK_0_H2_o(5) => \SHA256_BLOCK_0_H2_o[5]\, 
        SHA256_BLOCK_0_H2_o(4) => \SHA256_BLOCK_0_H2_o[4]\, 
        SHA256_BLOCK_0_H2_o(3) => \SHA256_BLOCK_0_H2_o[3]\, 
        SHA256_BLOCK_0_H2_o(2) => \SHA256_BLOCK_0_H2_o[2]\, 
        SHA256_BLOCK_0_H2_o(1) => \SHA256_BLOCK_0_H2_o[1]\, 
        SHA256_BLOCK_0_H2_o(0) => \SHA256_BLOCK_0_H2_o[0]\, 
        SHA256_BLOCK_0_H3_o(31) => \SHA256_BLOCK_0_H3_o[31]\, 
        SHA256_BLOCK_0_H3_o(30) => \SHA256_BLOCK_0_H3_o[30]\, 
        SHA256_BLOCK_0_H3_o(29) => \SHA256_BLOCK_0_H3_o[29]\, 
        SHA256_BLOCK_0_H3_o(28) => \SHA256_BLOCK_0_H3_o[28]\, 
        SHA256_BLOCK_0_H3_o(27) => \SHA256_BLOCK_0_H3_o[27]\, 
        SHA256_BLOCK_0_H3_o(26) => \SHA256_BLOCK_0_H3_o[26]\, 
        SHA256_BLOCK_0_H3_o(25) => \SHA256_BLOCK_0_H3_o[25]\, 
        SHA256_BLOCK_0_H3_o(24) => \SHA256_BLOCK_0_H3_o[24]\, 
        SHA256_BLOCK_0_H3_o(23) => \SHA256_BLOCK_0_H3_o[23]\, 
        SHA256_BLOCK_0_H3_o(22) => \SHA256_BLOCK_0_H3_o[22]\, 
        SHA256_BLOCK_0_H3_o(21) => \SHA256_BLOCK_0_H3_o[21]\, 
        SHA256_BLOCK_0_H3_o(20) => \SHA256_BLOCK_0_H3_o[20]\, 
        SHA256_BLOCK_0_H3_o(19) => \SHA256_BLOCK_0_H3_o[19]\, 
        SHA256_BLOCK_0_H3_o(18) => \SHA256_BLOCK_0_H3_o[18]\, 
        SHA256_BLOCK_0_H3_o(17) => \SHA256_BLOCK_0_H3_o[17]\, 
        SHA256_BLOCK_0_H3_o(16) => \SHA256_BLOCK_0_H3_o[16]\, 
        SHA256_BLOCK_0_H3_o(15) => \SHA256_BLOCK_0_H3_o[15]\, 
        SHA256_BLOCK_0_H3_o(14) => \SHA256_BLOCK_0_H3_o[14]\, 
        SHA256_BLOCK_0_H3_o(13) => \SHA256_BLOCK_0_H3_o[13]\, 
        SHA256_BLOCK_0_H3_o(12) => \SHA256_BLOCK_0_H3_o[12]\, 
        SHA256_BLOCK_0_H3_o(11) => \SHA256_BLOCK_0_H3_o[11]\, 
        SHA256_BLOCK_0_H3_o(10) => \SHA256_BLOCK_0_H3_o[10]\, 
        SHA256_BLOCK_0_H3_o(9) => \SHA256_BLOCK_0_H3_o[9]\, 
        SHA256_BLOCK_0_H3_o(8) => \SHA256_BLOCK_0_H3_o[8]\, 
        SHA256_BLOCK_0_H3_o(7) => \SHA256_BLOCK_0_H3_o[7]\, 
        SHA256_BLOCK_0_H3_o(6) => \SHA256_BLOCK_0_H3_o[6]\, 
        SHA256_BLOCK_0_H3_o(5) => \SHA256_BLOCK_0_H3_o[5]\, 
        SHA256_BLOCK_0_H3_o(4) => \SHA256_BLOCK_0_H3_o[4]\, 
        SHA256_BLOCK_0_H3_o(3) => \SHA256_BLOCK_0_H3_o[3]\, 
        SHA256_BLOCK_0_H3_o(2) => \SHA256_BLOCK_0_H3_o[2]\, 
        SHA256_BLOCK_0_H3_o(1) => \SHA256_BLOCK_0_H3_o[1]\, 
        SHA256_BLOCK_0_H3_o(0) => \SHA256_BLOCK_0_H3_o[0]\, 
        SHA256_BLOCK_0_H4_o(31) => \SHA256_BLOCK_0_H4_o[31]\, 
        SHA256_BLOCK_0_H4_o(30) => \SHA256_BLOCK_0_H4_o[30]\, 
        SHA256_BLOCK_0_H4_o(29) => \SHA256_BLOCK_0_H4_o[29]\, 
        SHA256_BLOCK_0_H4_o(28) => \SHA256_BLOCK_0_H4_o[28]\, 
        SHA256_BLOCK_0_H4_o(27) => \SHA256_BLOCK_0_H4_o[27]\, 
        SHA256_BLOCK_0_H4_o(26) => \SHA256_BLOCK_0_H4_o[26]\, 
        SHA256_BLOCK_0_H4_o(25) => \SHA256_BLOCK_0_H4_o[25]\, 
        SHA256_BLOCK_0_H4_o(24) => \SHA256_BLOCK_0_H4_o[24]\, 
        SHA256_BLOCK_0_H4_o(23) => \SHA256_BLOCK_0_H4_o[23]\, 
        SHA256_BLOCK_0_H4_o(22) => \SHA256_BLOCK_0_H4_o[22]\, 
        SHA256_BLOCK_0_H4_o(21) => \SHA256_BLOCK_0_H4_o[21]\, 
        SHA256_BLOCK_0_H4_o(20) => \SHA256_BLOCK_0_H4_o[20]\, 
        SHA256_BLOCK_0_H4_o(19) => \SHA256_BLOCK_0_H4_o[19]\, 
        SHA256_BLOCK_0_H4_o(18) => \SHA256_BLOCK_0_H4_o[18]\, 
        SHA256_BLOCK_0_H4_o(17) => \SHA256_BLOCK_0_H4_o[17]\, 
        SHA256_BLOCK_0_H4_o(16) => \SHA256_BLOCK_0_H4_o[16]\, 
        SHA256_BLOCK_0_H4_o(15) => \SHA256_BLOCK_0_H4_o[15]\, 
        SHA256_BLOCK_0_H4_o(14) => \SHA256_BLOCK_0_H4_o[14]\, 
        SHA256_BLOCK_0_H4_o(13) => \SHA256_BLOCK_0_H4_o[13]\, 
        SHA256_BLOCK_0_H4_o(12) => \SHA256_BLOCK_0_H4_o[12]\, 
        SHA256_BLOCK_0_H4_o(11) => \SHA256_BLOCK_0_H4_o[11]\, 
        SHA256_BLOCK_0_H4_o(10) => \SHA256_BLOCK_0_H4_o[10]\, 
        SHA256_BLOCK_0_H4_o(9) => \SHA256_BLOCK_0_H4_o[9]\, 
        SHA256_BLOCK_0_H4_o(8) => \SHA256_BLOCK_0_H4_o[8]\, 
        SHA256_BLOCK_0_H4_o(7) => \SHA256_BLOCK_0_H4_o[7]\, 
        SHA256_BLOCK_0_H4_o(6) => \SHA256_BLOCK_0_H4_o[6]\, 
        SHA256_BLOCK_0_H4_o(5) => \SHA256_BLOCK_0_H4_o[5]\, 
        SHA256_BLOCK_0_H4_o(4) => \SHA256_BLOCK_0_H4_o[4]\, 
        SHA256_BLOCK_0_H4_o(3) => \SHA256_BLOCK_0_H4_o[3]\, 
        SHA256_BLOCK_0_H4_o(2) => \SHA256_BLOCK_0_H4_o[2]\, 
        SHA256_BLOCK_0_H4_o(1) => \SHA256_BLOCK_0_H4_o[1]\, 
        SHA256_BLOCK_0_H4_o(0) => \SHA256_BLOCK_0_H4_o[0]\, 
        SHA256_BLOCK_0_H5_o(31) => \SHA256_BLOCK_0_H5_o[31]\, 
        SHA256_BLOCK_0_H5_o(30) => \SHA256_BLOCK_0_H5_o[30]\, 
        SHA256_BLOCK_0_H5_o(29) => \SHA256_BLOCK_0_H5_o[29]\, 
        SHA256_BLOCK_0_H5_o(28) => \SHA256_BLOCK_0_H5_o[28]\, 
        SHA256_BLOCK_0_H5_o(27) => \SHA256_BLOCK_0_H5_o[27]\, 
        SHA256_BLOCK_0_H5_o(26) => \SHA256_BLOCK_0_H5_o[26]\, 
        SHA256_BLOCK_0_H5_o(25) => \SHA256_BLOCK_0_H5_o[25]\, 
        SHA256_BLOCK_0_H5_o(24) => \SHA256_BLOCK_0_H5_o[24]\, 
        SHA256_BLOCK_0_H5_o(23) => \SHA256_BLOCK_0_H5_o[23]\, 
        SHA256_BLOCK_0_H5_o(22) => \SHA256_BLOCK_0_H5_o[22]\, 
        SHA256_BLOCK_0_H5_o(21) => \SHA256_BLOCK_0_H5_o[21]\, 
        SHA256_BLOCK_0_H5_o(20) => \SHA256_BLOCK_0_H5_o[20]\, 
        SHA256_BLOCK_0_H5_o(19) => \SHA256_BLOCK_0_H5_o[19]\, 
        SHA256_BLOCK_0_H5_o(18) => \SHA256_BLOCK_0_H5_o[18]\, 
        SHA256_BLOCK_0_H5_o(17) => \SHA256_BLOCK_0_H5_o[17]\, 
        SHA256_BLOCK_0_H5_o(16) => \SHA256_BLOCK_0_H5_o[16]\, 
        SHA256_BLOCK_0_H5_o(15) => \SHA256_BLOCK_0_H5_o[15]\, 
        SHA256_BLOCK_0_H5_o(14) => \SHA256_BLOCK_0_H5_o[14]\, 
        SHA256_BLOCK_0_H5_o(13) => \SHA256_BLOCK_0_H5_o[13]\, 
        SHA256_BLOCK_0_H5_o(12) => \SHA256_BLOCK_0_H5_o[12]\, 
        SHA256_BLOCK_0_H5_o(11) => \SHA256_BLOCK_0_H5_o[11]\, 
        SHA256_BLOCK_0_H5_o(10) => \SHA256_BLOCK_0_H5_o[10]\, 
        SHA256_BLOCK_0_H5_o(9) => \SHA256_BLOCK_0_H5_o[9]\, 
        SHA256_BLOCK_0_H5_o(8) => \SHA256_BLOCK_0_H5_o[8]\, 
        SHA256_BLOCK_0_H5_o(7) => \SHA256_BLOCK_0_H5_o[7]\, 
        SHA256_BLOCK_0_H5_o(6) => \SHA256_BLOCK_0_H5_o[6]\, 
        SHA256_BLOCK_0_H5_o(5) => \SHA256_BLOCK_0_H5_o[5]\, 
        SHA256_BLOCK_0_H5_o(4) => \SHA256_BLOCK_0_H5_o[4]\, 
        SHA256_BLOCK_0_H5_o(3) => \SHA256_BLOCK_0_H5_o[3]\, 
        SHA256_BLOCK_0_H5_o(2) => \SHA256_BLOCK_0_H5_o[2]\, 
        SHA256_BLOCK_0_H5_o(1) => \SHA256_BLOCK_0_H5_o[1]\, 
        SHA256_BLOCK_0_H5_o(0) => \SHA256_BLOCK_0_H5_o[0]\, 
        SHA256_BLOCK_0_H6_o(31) => \SHA256_BLOCK_0_H6_o[31]\, 
        SHA256_BLOCK_0_H6_o(30) => \SHA256_BLOCK_0_H6_o[30]\, 
        SHA256_BLOCK_0_H6_o(29) => \SHA256_BLOCK_0_H6_o[29]\, 
        SHA256_BLOCK_0_H6_o(28) => \SHA256_BLOCK_0_H6_o[28]\, 
        SHA256_BLOCK_0_H6_o(27) => \SHA256_BLOCK_0_H6_o[27]\, 
        SHA256_BLOCK_0_H6_o(26) => \SHA256_BLOCK_0_H6_o[26]\, 
        SHA256_BLOCK_0_H6_o(25) => \SHA256_BLOCK_0_H6_o[25]\, 
        SHA256_BLOCK_0_H6_o(24) => \SHA256_BLOCK_0_H6_o[24]\, 
        SHA256_BLOCK_0_H6_o(23) => \SHA256_BLOCK_0_H6_o[23]\, 
        SHA256_BLOCK_0_H6_o(22) => \SHA256_BLOCK_0_H6_o[22]\, 
        SHA256_BLOCK_0_H6_o(21) => \SHA256_BLOCK_0_H6_o[21]\, 
        SHA256_BLOCK_0_H6_o(20) => \SHA256_BLOCK_0_H6_o[20]\, 
        SHA256_BLOCK_0_H6_o(19) => \SHA256_BLOCK_0_H6_o[19]\, 
        SHA256_BLOCK_0_H6_o(18) => \SHA256_BLOCK_0_H6_o[18]\, 
        SHA256_BLOCK_0_H6_o(17) => \SHA256_BLOCK_0_H6_o[17]\, 
        SHA256_BLOCK_0_H6_o(16) => \SHA256_BLOCK_0_H6_o[16]\, 
        SHA256_BLOCK_0_H6_o(15) => \SHA256_BLOCK_0_H6_o[15]\, 
        SHA256_BLOCK_0_H6_o(14) => \SHA256_BLOCK_0_H6_o[14]\, 
        SHA256_BLOCK_0_H6_o(13) => \SHA256_BLOCK_0_H6_o[13]\, 
        SHA256_BLOCK_0_H6_o(12) => \SHA256_BLOCK_0_H6_o[12]\, 
        SHA256_BLOCK_0_H6_o(11) => \SHA256_BLOCK_0_H6_o[11]\, 
        SHA256_BLOCK_0_H6_o(10) => \SHA256_BLOCK_0_H6_o[10]\, 
        SHA256_BLOCK_0_H6_o(9) => \SHA256_BLOCK_0_H6_o[9]\, 
        SHA256_BLOCK_0_H6_o(8) => \SHA256_BLOCK_0_H6_o[8]\, 
        SHA256_BLOCK_0_H6_o(7) => \SHA256_BLOCK_0_H6_o[7]\, 
        SHA256_BLOCK_0_H6_o(6) => \SHA256_BLOCK_0_H6_o[6]\, 
        SHA256_BLOCK_0_H6_o(5) => \SHA256_BLOCK_0_H6_o[5]\, 
        SHA256_BLOCK_0_H6_o(4) => \SHA256_BLOCK_0_H6_o[4]\, 
        SHA256_BLOCK_0_H6_o(3) => \SHA256_BLOCK_0_H6_o[3]\, 
        SHA256_BLOCK_0_H6_o(2) => \SHA256_BLOCK_0_H6_o[2]\, 
        SHA256_BLOCK_0_H6_o(1) => \SHA256_BLOCK_0_H6_o[1]\, 
        SHA256_BLOCK_0_H6_o(0) => \SHA256_BLOCK_0_H6_o[0]\, 
        SHA256_BLOCK_0_H7_o(31) => \SHA256_BLOCK_0_H7_o[31]\, 
        SHA256_BLOCK_0_H7_o(30) => \SHA256_BLOCK_0_H7_o[30]\, 
        SHA256_BLOCK_0_H7_o(29) => \SHA256_BLOCK_0_H7_o[29]\, 
        SHA256_BLOCK_0_H7_o(28) => \SHA256_BLOCK_0_H7_o[28]\, 
        SHA256_BLOCK_0_H7_o(27) => \SHA256_BLOCK_0_H7_o[27]\, 
        SHA256_BLOCK_0_H7_o(26) => \SHA256_BLOCK_0_H7_o[26]\, 
        SHA256_BLOCK_0_H7_o(25) => \SHA256_BLOCK_0_H7_o[25]\, 
        SHA256_BLOCK_0_H7_o(24) => \SHA256_BLOCK_0_H7_o[24]\, 
        SHA256_BLOCK_0_H7_o(23) => \SHA256_BLOCK_0_H7_o[23]\, 
        SHA256_BLOCK_0_H7_o(22) => \SHA256_BLOCK_0_H7_o[22]\, 
        SHA256_BLOCK_0_H7_o(21) => \SHA256_BLOCK_0_H7_o[21]\, 
        SHA256_BLOCK_0_H7_o(20) => \SHA256_BLOCK_0_H7_o[20]\, 
        SHA256_BLOCK_0_H7_o(19) => \SHA256_BLOCK_0_H7_o[19]\, 
        SHA256_BLOCK_0_H7_o(18) => \SHA256_BLOCK_0_H7_o[18]\, 
        SHA256_BLOCK_0_H7_o(17) => \SHA256_BLOCK_0_H7_o[17]\, 
        SHA256_BLOCK_0_H7_o(16) => \SHA256_BLOCK_0_H7_o[16]\, 
        SHA256_BLOCK_0_H7_o(15) => \SHA256_BLOCK_0_H7_o[15]\, 
        SHA256_BLOCK_0_H7_o(14) => \SHA256_BLOCK_0_H7_o[14]\, 
        SHA256_BLOCK_0_H7_o(13) => \SHA256_BLOCK_0_H7_o[13]\, 
        SHA256_BLOCK_0_H7_o(12) => \SHA256_BLOCK_0_H7_o[12]\, 
        SHA256_BLOCK_0_H7_o(11) => \SHA256_BLOCK_0_H7_o[11]\, 
        SHA256_BLOCK_0_H7_o(10) => \SHA256_BLOCK_0_H7_o[10]\, 
        SHA256_BLOCK_0_H7_o(9) => \SHA256_BLOCK_0_H7_o[9]\, 
        SHA256_BLOCK_0_H7_o(8) => \SHA256_BLOCK_0_H7_o[8]\, 
        SHA256_BLOCK_0_H7_o(7) => \SHA256_BLOCK_0_H7_o[7]\, 
        SHA256_BLOCK_0_H7_o(6) => \SHA256_BLOCK_0_H7_o[6]\, 
        SHA256_BLOCK_0_H7_o(5) => \SHA256_BLOCK_0_H7_o[5]\, 
        SHA256_BLOCK_0_H7_o(4) => \SHA256_BLOCK_0_H7_o[4]\, 
        SHA256_BLOCK_0_H7_o(3) => \SHA256_BLOCK_0_H7_o[3]\, 
        SHA256_BLOCK_0_H7_o(2) => \SHA256_BLOCK_0_H7_o[2]\, 
        SHA256_BLOCK_0_H7_o(1) => \SHA256_BLOCK_0_H7_o[1]\, 
        SHA256_BLOCK_0_H7_o(0) => \SHA256_BLOCK_0_H7_o[0]\, 
        SHA256_Module_0_data_out_5 => SHA256_Module_0_data_out_5, 
        SHA256_Module_0_data_out_13 => 
        SHA256_Module_0_data_out_13, SHA256_Module_0_data_out_12
         => SHA256_Module_0_data_out_12, 
        SHA256_Module_0_data_out_23 => 
        SHA256_Module_0_data_out_23, SHA256_Module_0_data_out_8
         => SHA256_Module_0_data_out_8, 
        SHA256_Module_0_data_out_0 => SHA256_Module_0_data_out_0, 
        line_1_d0 => line_0_d0, line_2_d0 => line_1_d0, line_3_d0
         => line_2_d0, line_4_d0 => line_3_d0, line_6_d0 => 
        line_5_d0, line_7_d0 => line_6_d0, line_9 => line_8, 
        line_10 => line_9, line_11 => line_10, line_14 => line_13, 
        line_15 => line_14, line_16 => line_15, line_17 => 
        line_16, line_18 => line_17, line_19 => line_18, line_20
         => line_19, line_21 => line_20, line_22 => line_21, 
        line_24 => line_23, line_25 => line_24, line_26 => 
        line_25, line_27 => line_26, line_29 => line_28, line_30
         => line_29, line_0_1 => line_0_0, line_0_2 => line_0_1, 
        line_0_3 => line_0_2, line_0_4 => line_0_3, line_0_6 => 
        line_0_5, line_0_7 => line_0_6, line_0_9 => line_0_8, 
        line_0_10 => line_0_9, line_0_11 => line_0_10, line_0_14
         => line_0_13, line_0_15 => line_0_14, line_0_16 => 
        line_0_15, line_0_17 => line_0_16, line_0_18 => line_0_17, 
        line_0_19 => line_0_18, line_0_20 => line_0_19, line_0_21
         => line_0_20, line_0_22 => line_0_21, line_0_24 => 
        line_0_23, line_0_25 => line_0_24, line_0_26 => line_0_25, 
        line_0_27 => line_0_26, line_0_29 => line_0_28, line_0_30
         => line_0_29, line_1_1 => line_1_0, line_1_2 => line_1_1, 
        line_1_3 => line_1_2, line_1_4 => line_1_3, line_1_6 => 
        line_1_5, line_1_7 => line_1_6, line_1_9 => line_1_8, 
        line_1_10 => line_1_9, line_1_11 => line_1_10, line_1_14
         => line_1_13, line_1_15 => line_1_14, line_1_16 => 
        line_1_15, line_1_17 => line_1_16, line_1_18 => line_1_17, 
        line_1_19 => line_1_18, line_1_20 => line_1_19, line_1_21
         => line_1_20, line_1_22 => line_1_21, line_1_24 => 
        line_1_23, line_1_25 => line_1_24, line_1_26 => line_1_25, 
        line_1_27 => line_1_26, line_1_29 => line_1_28, line_1_30
         => line_1_29, line_2_1 => line_2_0, line_2_2 => line_2_1, 
        line_2_3 => line_2_2, line_2_4 => line_2_3, line_2_6 => 
        line_2_5, line_2_7 => line_2_6, line_2_9 => line_2_8, 
        line_2_10 => line_2_9, line_2_11 => line_2_10, line_2_14
         => line_2_13, line_2_15 => line_2_14, line_2_16 => 
        line_2_15, line_2_17 => line_2_16, line_2_18 => line_2_17, 
        line_2_19 => line_2_18, line_2_20 => line_2_19, line_2_21
         => line_2_20, line_2_22 => line_2_21, line_2_24 => 
        line_2_23, line_2_25 => line_2_24, line_2_26 => line_2_25, 
        line_2_27 => line_2_26, line_2_29 => line_2_28, line_2_30
         => line_2_29, line_3_28 => line_27, line_3_31 => line_30, 
        line_3_1 => line_3_0, line_3_2 => line_3_1, line_3_3 => 
        line_3_2, line_3_4 => line_3_3, line_3_6 => line_3_5, 
        line_3_7 => line_3_6, line_3_9 => line_3_8, line_3_10 => 
        line_3_9, line_3_11 => line_3_10, line_3_14 => line_3_13, 
        line_3_15 => line_3_14, line_3_16 => line_3_15, line_3_17
         => line_3_16, line_3_18 => line_3_17, line_3_19 => 
        line_3_18, line_3_20 => line_3_19, line_3_21 => line_3_20, 
        line_3_22 => line_3_21, line_3_24 => line_3_23, line_3_25
         => line_3_24, line_3_26 => line_3_25, line_3_27 => 
        line_3_26, line_3_29 => line_3_28, line_3_30 => line_3_29, 
        line_4_28 => line_0_27, line_4_31 => line_0_30, line_4_1
         => line_4_0, line_4_2 => line_4_1, line_4_3 => line_4_2, 
        line_4_4 => line_4_3, line_4_6 => line_4_5, line_4_7 => 
        line_4_6, line_4_9 => line_4_8, line_4_10 => line_4_9, 
        line_4_11 => line_4_10, line_4_14 => line_4_13, line_4_15
         => line_4_14, line_4_16 => line_4_15, line_4_17 => 
        line_4_16, line_4_18 => line_4_17, line_4_19 => line_4_18, 
        line_4_20 => line_4_19, line_4_21 => line_4_20, line_4_22
         => line_4_21, line_4_24 => line_4_23, line_4_25 => 
        line_4_24, line_4_26 => line_4_25, line_4_27 => line_4_26, 
        line_4_29 => line_4_28, line_4_30 => line_4_29, line_5_28
         => line_1_27, line_5_31 => line_1_30, line_5_1 => 
        line_5_0, line_5_2 => line_5_1, line_5_3 => line_5_2, 
        line_5_4 => line_5_3, line_5_6 => line_5_5, line_5_7 => 
        line_5_6, line_5_9 => line_5_8, line_5_10 => line_5_9, 
        line_5_11 => line_5_10, line_5_14 => line_5_13, line_5_15
         => line_5_14, line_5_16 => line_5_15, line_5_17 => 
        line_5_16, line_5_18 => line_5_17, line_5_19 => line_5_18, 
        line_5_20 => line_5_19, line_5_21 => line_5_20, line_5_22
         => line_5_21, line_5_24 => line_5_23, line_5_25 => 
        line_5_24, line_5_26 => line_5_25, line_5_27 => line_5_26, 
        line_5_29 => line_5_28, line_5_30 => line_5_29, line_6_1
         => line_6_0, line_6_2 => line_6_1, line_6_3 => line_6_2, 
        line_6_4 => line_6_3, line_6_6 => line_6_5, line_6_7 => 
        line_6_6, line_6_9 => line_6_8, line_6_10 => line_6_9, 
        line_6_11 => line_6_10, line_6_14 => line_6_13, line_6_15
         => line_6_14, line_6_16 => line_6_15, line_6_17 => 
        line_6_16, line_6_18 => line_6_17, line_6_19 => line_6_18, 
        line_6_20 => line_6_19, line_6_21 => line_6_20, line_6_22
         => line_6_21, line_6_24 => line_6_23, line_6_25 => 
        line_6_24, line_6_26 => line_6_25, line_6_27 => line_6_26, 
        line_6_28 => line_2_27, line_6_29 => line_6_28, line_6_30
         => line_6_29, line_6_31 => line_2_30, line_7_1 => 
        line_7(1), line_7_2 => line_7(2), N_507 => N_507, N_508
         => N_508, ren_pos => ren_pos, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, data_out_ready => 
        data_out_ready, AHB_slave_dummy_0_read_en => 
        AHB_slave_dummy_0_read_en, start_wen => start_wen, 
        SHA256_Module_0_error_o => \SHA256_Module_0_error_o\, 
        SHA256_Module_0_di_req_o => \SHA256_Module_0_di_req_o\, 
        SHA256_Module_0_do_valid_o => 
        \SHA256_Module_0_do_valid_o\);
    
    reg1_highonly_0 : reg1_highonly
      port map(CertificationSystem_sb_0_GPIO_9_M2F => 
        CertificationSystem_sb_0_GPIO_9_M2F, 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0 => 
        CertificationSystem_sb_0_GPIO_9_M2F_i_0, start_wen => 
        start_wen, CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, 
        SHA256_BLOCK_0_start_o => SHA256_BLOCK_0_start_o);
    
    AND2_0 : AND2
      port map(A => start_wen, B => SHA256_BLOCK_0_do_valid_o, Y
         => \SHA256_Module_0_do_valid_o\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_FABOSC_0_OSC is

    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );

end CertificationSystem_sb_FABOSC_0_OSC;

architecture DEF_ARCH of CertificationSystem_sb_FABOSC_0_OSC is 

  component RCOSC_25_50MHZ
    generic (FREQUENCY:real := 50.0);

    port( CLKOUT : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    I_RCOSC_25_50MHZ : RCOSC_25_50MHZ
      generic map(FREQUENCY => 50.0)

      port map(CLKOUT => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreResetP is

    port( MSS_READY                                             : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic;
          CertificationSystem_sb_0_POWER_ON_RESET_N             : in    std_logic
        );

end CoreResetP;

architecture DEF_ARCH of CoreResetP is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \MSS_HPMS_READY_int\, \mss_ready_select\, VCC_net_1, 
        \POWER_ON_RESET_N_clk_base\, 
        \un6_fic_2_apb_m_preset_n_clk_base\, GND_net_1, 
        \mss_ready_state\, \RESET_N_M2F_clk_base\, 
        \RESET_N_M2F_q1\, \FIC_2_APB_M_PRESET_N_q1\, 
        \POWER_ON_RESET_N_q1\, \FIC_2_APB_M_PRESET_N_clk_base\, 
        \MSS_HPMS_READY_int_3\ : std_logic;

begin 


    RESET_N_M2F_clk_base : SLE
      port map(D => \RESET_N_M2F_q1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RESET_N_M2F_clk_base\);
    
    POWER_ON_RESET_N_clk_base : SLE
      port map(D => \POWER_ON_RESET_N_q1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \POWER_ON_RESET_N_clk_base\);
    
    mss_ready_select : SLE
      port map(D => VCC_net_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \un6_fic_2_apb_m_preset_n_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_select\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    mss_ready_state : SLE
      port map(D => VCC_net_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        \RESET_N_M2F_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_state\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    un6_fic_2_apb_m_preset_n_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \FIC_2_APB_M_PRESET_N_clk_base\, B => 
        \mss_ready_state\, Y => 
        \un6_fic_2_apb_m_preset_n_clk_base\);
    
    RESET_N_M2F_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RESET_N_M2F_q1\);
    
    FIC_2_APB_M_PRESET_N_clk_base : SLE
      port map(D => \FIC_2_APB_M_PRESET_N_q1\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \FIC_2_APB_M_PRESET_N_clk_base\);
    
    POWER_ON_RESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \POWER_ON_RESET_N_q1\);
    
    MSS_HPMS_READY_int_RNIRS5B : CLKINT
      port map(A => \MSS_HPMS_READY_int\, Y => MSS_READY);
    
    FIC_2_APB_M_PRESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \FIC_2_APB_M_PRESET_N_q1\);
    
    MSS_HPMS_READY_int_3 : CFG3
      generic map(INIT => x"E0")

      port map(A => \RESET_N_M2F_clk_base\, B => 
        \mss_ready_select\, C => \FIC_2_APB_M_PRESET_N_clk_base\, 
        Y => \MSS_HPMS_READY_int_3\);
    
    MSS_HPMS_READY_int : SLE
      port map(D => \MSS_HPMS_READY_int_3\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \MSS_HPMS_READY_int\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVEARBITER_1_0 is

    port( arbRegSMCurrentState_ns_i_0                             : out   std_logic_vector(1 to 1);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR : in    std_logic_vector(5 downto 3);
          regHADDR                                                : in    std_logic_vector(5 downto 3);
          MSS_READY                                               : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                    : in    std_logic;
          N_127                                                   : in    std_logic;
          N_120                                                   : in    std_logic;
          N_226                                                   : out   std_logic;
          N_226_i_0                                               : out   std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY              : in    std_logic;
          masterRegAddrSel                                        : in    std_logic;
          N_218_i_0                                               : out   std_logic;
          N_217_i_0                                               : out   std_logic;
          N_203_i_0                                               : out   std_logic
        );

end COREAHBLITE_SLAVEARBITER_1_0;

architecture DEF_ARCH of COREAHBLITE_SLAVEARBITER_1_0 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \arbRegSMCurrentState[15]_net_1\, VCC_net_1, 
        N_109_i_0, GND_net_1, \arbRegSMCurrentState[14]_net_1\, 
        N_111_i_0, \arbRegSMCurrentState[10]_net_1\, N_81_i_0, 
        \arbRegSMCurrentState[6]_net_1\, N_79_i_0, 
        \arbRegSMCurrentState[2]_net_1\, N_220_i_0, 
        \arbRegSMCurrentState_ns_i_0_a2_1[1]_net_1\, N_306, N_188, 
        N_280, \N_226\ : std_logic;

begin 

    N_226 <= \N_226\;

    \arbRegSMCurrentState_RNO[2]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \arbRegSMCurrentState[2]_net_1\, B => N_120, 
        C => N_127, Y => N_220_i_0);
    
    \arbRegSMCurrentState_ns_i_0_a2_RNIOO6J[0]\ : CFG4
      generic map(INIT => x"3022")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(4), 
        B => \N_226\, C => regHADDR(4), D => masterRegAddrSel, Y
         => N_217_i_0);
    
    \arbRegSMCurrentState[10]\ : SLE
      port map(D => N_81_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[10]_net_1\);
    
    \arbRegSMCurrentState_RNO[10]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \arbRegSMCurrentState[10]_net_1\, B => N_120, 
        C => N_127, Y => N_81_i_0);
    
    \arbRegSMCurrentState[14]\ : SLE
      port map(D => N_111_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[14]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \arbRegSMCurrentState_ns_i_0_a2[0]\ : CFG4
      generic map(INIT => x"0F0E")

      port map(A => N_120, B => N_127, C => 
        \arbRegSMCurrentState[15]_net_1\, D => N_188, Y => 
        \N_226\);
    
    \arbRegSMCurrentState[15]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[15]_net_1\);
    
    \arbRegSMCurrentState_RNO[14]\ : CFG3
      generic map(INIT => x"0D")

      port map(A => N_280, B => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, C => N_306, Y
         => N_111_i_0);
    
    \arbRegSMCurrentState_ns_i_0_a2_RNIPP6J[0]\ : CFG4
      generic map(INIT => x"3022")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(5), 
        B => \N_226\, C => regHADDR(5), D => masterRegAddrSel, Y
         => N_218_i_0);
    
    \arbRegSMCurrentState_ns_i_0_a2_0[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \arbRegSMCurrentState[14]_net_1\, B => 
        \arbRegSMCurrentState[10]_net_1\, C => 
        \arbRegSMCurrentState[6]_net_1\, D => 
        \arbRegSMCurrentState[2]_net_1\, Y => N_188);
    
    \arbRegSMCurrentState_ns_i_0[1]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => N_280, B => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, C => N_306, Y
         => arbRegSMCurrentState_ns_i_0(1));
    
    \arbRegSMCurrentState_RNO[15]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \N_226\, B => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, Y => 
        N_109_i_0);
    
    \arbRegSMCurrentState_RNO[6]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \arbRegSMCurrentState[6]_net_1\, B => N_120, 
        C => N_127, Y => N_79_i_0);
    
    \arbRegSMCurrentState_ns_i_0_a2_RNINN6J[0]\ : CFG4
      generic map(INIT => x"3022")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(3), 
        B => \N_226\, C => regHADDR(3), D => masterRegAddrSel, Y
         => N_203_i_0);
    
    \arbRegSMCurrentState[6]\ : SLE
      port map(D => N_79_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[6]_net_1\);
    
    \arbRegSMCurrentState_ns_i_0_a2[1]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => \arbRegSMCurrentState[14]_net_1\, B => 
        \arbRegSMCurrentState[15]_net_1\, C => N_127, D => 
        \arbRegSMCurrentState_ns_i_0_a2_1[1]_net_1\, Y => N_306);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \arbRegSMCurrentState_ns_i_0_a2_1[1]\ : CFG4
      generic map(INIT => x"3332")

      port map(A => \arbRegSMCurrentState[2]_net_1\, B => N_120, 
        C => \arbRegSMCurrentState[10]_net_1\, D => 
        \arbRegSMCurrentState[6]_net_1\, Y => 
        \arbRegSMCurrentState_ns_i_0_a2_1[1]_net_1\);
    
    \arbRegSMCurrentState[2]\ : SLE
      port map(D => N_220_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[2]_net_1\);
    
    \arbRegSMCurrentState_ns_i_0_a2_0_RNIVU8H[0]\ : CFG4
      generic map(INIT => x"F0F1")

      port map(A => N_120, B => N_127, C => 
        \arbRegSMCurrentState[15]_net_1\, D => N_188, Y => 
        N_226_i_0);
    
    \arbRegSMCurrentState_ns_i_0_o3[1]\ : CFG3
      generic map(INIT => x"57")

      port map(A => \arbRegSMCurrentState[14]_net_1\, B => N_120, 
        C => N_127, Y => N_280);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVESTAGE_0 is

    port( masterDataInProg                                         : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA : in    std_logic_vector(31 downto 0);
          arbRegSMCurrentState_ns_i_0                              : out   std_logic_vector(1 to 1);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR  : in    std_logic_vector(5 downto 3);
          regHADDR                                                 : in    std_logic_vector(5 downto 3);
          MSS_READY                                                : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                     : in    std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY               : in    std_logic;
          N_65_i_0                                                 : out   std_logic;
          N_67_i_0                                                 : out   std_logic;
          N_110_i_0                                                : out   std_logic;
          N_112_i_0                                                : out   std_logic;
          N_114_i_0                                                : out   std_logic;
          N_116_i_0                                                : out   std_logic;
          N_69_i_0                                                 : out   std_logic;
          N_71_i_0                                                 : out   std_logic;
          N_73_i_0                                                 : out   std_logic;
          N_75_i_0                                                 : out   std_logic;
          N_77_i_0                                                 : out   std_logic;
          N_83_i_0                                                 : out   std_logic;
          N_85_i_0                                                 : out   std_logic;
          N_133_i_0                                                : out   std_logic;
          N_87_i_0                                                 : out   std_logic;
          N_89_i_0                                                 : out   std_logic;
          N_140_i_0                                                : out   std_logic;
          N_91_i_0                                                 : out   std_logic;
          N_93_i_0                                                 : out   std_logic;
          N_95_i_0                                                 : out   std_logic;
          N_97_i_0                                                 : out   std_logic;
          N_99_i_0                                                 : out   std_logic;
          N_152_i_0                                                : out   std_logic;
          N_101_i_0                                                : out   std_logic;
          N_156_i_0                                                : out   std_logic;
          N_158_i_0                                                : out   std_logic;
          N_103_i_0                                                : out   std_logic;
          N_105_i_0                                                : out   std_logic;
          N_107_i_0                                                : out   std_logic;
          N_168_i_0                                                : out   std_logic;
          N_109_i_0                                                : out   std_logic;
          N_111_i_0                                                : out   std_logic;
          N_127                                                    : in    std_logic;
          N_120                                                    : in    std_logic;
          N_226                                                    : out   std_logic;
          masterRegAddrSel                                         : in    std_logic;
          N_218_i_0                                                : out   std_logic;
          N_217_i_0                                                : out   std_logic;
          N_203_i_0                                                : out   std_logic
        );

end COREAHBLITE_SLAVESTAGE_0;

architecture DEF_ARCH of COREAHBLITE_SLAVESTAGE_0 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVEARBITER_1_0
    port( arbRegSMCurrentState_ns_i_0                             : out   std_logic_vector(1 to 1);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR : in    std_logic_vector(5 downto 3) := (others => 'U');
          regHADDR                                                : in    std_logic_vector(5 downto 3) := (others => 'U');
          MSS_READY                                               : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                    : in    std_logic := 'U';
          N_127                                                   : in    std_logic := 'U';
          N_120                                                   : in    std_logic := 'U';
          N_226                                                   : out   std_logic;
          N_226_i_0                                               : out   std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY              : in    std_logic := 'U';
          masterRegAddrSel                                        : in    std_logic := 'U';
          N_218_i_0                                               : out   std_logic;
          N_217_i_0                                               : out   std_logic;
          N_203_i_0                                               : out   std_logic
        );
  end component;

    signal \masterDataInProg[0]_net_1\, VCC_net_1, N_226_i_0, 
        GND_net_1 : std_logic;

    for all : COREAHBLITE_SLAVEARBITER_1_0
	Use entity work.COREAHBLITE_SLAVEARBITER_1_0(DEF_ARCH);
begin 

    masterDataInProg(0) <= \masterDataInProg[0]_net_1\;

    \masterDataInProg_RNIEMMC_3[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        B => \masterDataInProg[0]_net_1\, Y => N_168_i_0);
    
    \masterDataInProg_RNIEMMC_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        B => \masterDataInProg[0]_net_1\, Y => N_107_i_0);
    
    \masterDataInProg_RNIEMMC_14[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        B => \masterDataInProg[0]_net_1\, Y => N_110_i_0);
    
    \masterDataInProg_RNIEMMC_22[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        B => \masterDataInProg[0]_net_1\, Y => N_93_i_0);
    
    \masterDataInProg_RNIEMMC_15[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        B => \masterDataInProg[0]_net_1\, Y => N_105_i_0);
    
    \masterDataInProg_RNIEMMC_16[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        B => \masterDataInProg[0]_net_1\, Y => N_103_i_0);
    
    \masterDataInProg_RNIEMMC_18[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        B => \masterDataInProg[0]_net_1\, Y => N_156_i_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \masterDataInProg_RNIEMMC_27[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        B => \masterDataInProg[0]_net_1\, Y => N_133_i_0);
    
    \masterDataInProg_RNIEMMC_23[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        B => \masterDataInProg[0]_net_1\, Y => N_91_i_0);
    
    \masterDataInProg_RNIEMMC_29[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        B => \masterDataInProg[0]_net_1\, Y => N_83_i_0);
    
    \masterDataInProg_RNIEMMC_11[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        B => \masterDataInProg[0]_net_1\, Y => N_116_i_0);
    
    \masterDataInProg_RNIEMMC_9[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        B => \masterDataInProg[0]_net_1\, Y => N_71_i_0);
    
    \masterDataInProg_RNIEMMC_10[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        B => \masterDataInProg[0]_net_1\, Y => N_69_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \masterDataInProg[0]\ : SLE
      port map(D => N_226_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \masterDataInProg[0]_net_1\);
    
    \masterDataInProg_RNIEMMC_7[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        B => \masterDataInProg[0]_net_1\, Y => N_75_i_0);
    
    \masterDataInProg_RNIEMMC_30[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        B => \masterDataInProg[0]_net_1\, Y => N_77_i_0);
    
    \masterDataInProg_RNIEMMC_24[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        B => \masterDataInProg[0]_net_1\, Y => N_140_i_0);
    
    \masterDataInProg_RNIEMMC[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        B => \masterDataInProg[0]_net_1\, Y => N_67_i_0);
    
    \masterDataInProg_RNIEMMC_25[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        B => \masterDataInProg[0]_net_1\, Y => N_89_i_0);
    
    \masterDataInProg_RNIEMMC_26[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        B => \masterDataInProg[0]_net_1\, Y => N_87_i_0);
    
    \masterDataInProg_RNIEMMC_28[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        B => \masterDataInProg[0]_net_1\, Y => N_85_i_0);
    
    \masterDataInProg_RNIEMMC_1[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        B => \masterDataInProg[0]_net_1\, Y => N_111_i_0);
    
    \masterDataInProg_RNIEMMC_6[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        B => \masterDataInProg[0]_net_1\, Y => N_97_i_0);
    
    \masterDataInProg_RNIEMMC_12[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        B => \masterDataInProg[0]_net_1\, Y => N_114_i_0);
    
    slave_arbiter : COREAHBLITE_SLAVEARBITER_1_0
      port map(arbRegSMCurrentState_ns_i_0(1) => 
        arbRegSMCurrentState_ns_i_0(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(5)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(5), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(4)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(4), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(3)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(3), 
        regHADDR(5) => regHADDR(5), regHADDR(4) => regHADDR(4), 
        regHADDR(3) => regHADDR(3), MSS_READY => MSS_READY, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, N_127 => N_127, 
        N_120 => N_120, N_226 => N_226, N_226_i_0 => N_226_i_0, 
        CertificationSystem_sb_0_AHBmslave5_HREADY => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, 
        masterRegAddrSel => masterRegAddrSel, N_218_i_0 => 
        N_218_i_0, N_217_i_0 => N_217_i_0, N_203_i_0 => N_203_i_0);
    
    \masterDataInProg_RNIEMMC_8[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        B => \masterDataInProg[0]_net_1\, Y => N_73_i_0);
    
    \masterDataInProg_RNIEMMC_21[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        B => \masterDataInProg[0]_net_1\, Y => N_95_i_0);
    
    \masterDataInProg_RNIEMMC_20[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        B => \masterDataInProg[0]_net_1\, Y => N_152_i_0);
    
    \masterDataInProg_RNIEMMC_2[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        B => \masterDataInProg[0]_net_1\, Y => N_109_i_0);
    
    \masterDataInProg_RNIEMMC_5[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        B => \masterDataInProg[0]_net_1\, Y => N_99_i_0);
    
    \masterDataInProg_RNIEMMC_17[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        B => \masterDataInProg[0]_net_1\, Y => N_158_i_0);
    
    \masterDataInProg_RNIEMMC_13[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        B => \masterDataInProg[0]_net_1\, Y => N_112_i_0);
    
    \masterDataInProg_RNIEMMC_19[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        B => \masterDataInProg[0]_net_1\, Y => N_101_i_0);
    
    \masterDataInProg_RNIEMMC_0[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        B => \masterDataInProg[0]_net_1\, Y => N_65_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVEARBITER_1 is

    port( xhdl1221                                                  : in    std_logic_vector(3 to 3);
          CoreAHBLite_0_AHBmslave3_HADDR                            : out   std_logic_vector(11 to 11);
          arbRegSMCurrentState_13                                   : out   std_logic;
          arbRegSMCurrentState_12                                   : out   std_logic;
          arbRegSMCurrentState_8                                    : out   std_logic;
          arbRegSMCurrentState_4                                    : out   std_logic;
          arbRegSMCurrentState_0                                    : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 : in    std_logic;
          regHADDR_8                                                : in    std_logic;
          regHADDR_2                                                : in    std_logic;
          regHADDR_1                                                : in    std_logic;
          regHADDR_0                                                : in    std_logic;
          MSS_READY                                                 : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                      : in    std_logic;
          N_271                                                     : in    std_logic;
          N_120                                                     : in    std_logic;
          N_225                                                     : in    std_logic;
          N_157_i_i_o2_0                                            : out   std_logic;
          N_148                                                     : in    std_logic;
          N_138                                                     : in    std_logic;
          N_149                                                     : in    std_logic;
          N_157_i_i_o2_0_out                                        : out   std_logic;
          hsel2_i_4                                                 : out   std_logic;
          N_135                                                     : in    std_logic;
          masterRegAddrSel                                          : in    std_logic;
          hsel2_i_4_i_0                                             : out   std_logic;
          N_196_i_0                                                 : out   std_logic;
          N_195_i_0                                                 : out   std_logic;
          N_194_i_0                                                 : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                       : in    std_logic
        );

end COREAHBLITE_SLAVEARBITER_1;

architecture DEF_ARCH of COREAHBLITE_SLAVEARBITER_1 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \arbRegSMCurrentState_13\, VCC_net_1, N_109_i_0, 
        GND_net_1, \arbRegSMCurrentState_12\, 
        \arbRegSMCurrentState_ns_i_i[1]_net_1\, 
        \arbRegSMCurrentState_8\, N_104_i_0, 
        \arbRegSMCurrentState_4\, N_102_i_0, 
        \arbRegSMCurrentState_0\, N_100_i_0, \N_157_i_i_o2_0\, 
        \N_157_i_i_o2_0_out\, \hsel2_i_4\ : std_logic;

begin 

    arbRegSMCurrentState_13 <= \arbRegSMCurrentState_13\;
    arbRegSMCurrentState_12 <= \arbRegSMCurrentState_12\;
    arbRegSMCurrentState_8 <= \arbRegSMCurrentState_8\;
    arbRegSMCurrentState_4 <= \arbRegSMCurrentState_4\;
    arbRegSMCurrentState_0 <= \arbRegSMCurrentState_0\;
    N_157_i_i_o2_0 <= \N_157_i_i_o2_0\;
    N_157_i_i_o2_0_out <= \N_157_i_i_o2_0_out\;
    hsel2_i_4 <= \hsel2_i_4\;

    N_157_i_i_o2_0_0 : CFG2
      generic map(INIT => x"B")

      port map(A => N_120, B => N_225, Y => \N_157_i_i_o2_0\);
    
    \arbRegSMCurrentState_RNO[2]\ : CFG4
      generic map(INIT => x"CCC8")

      port map(A => N_120, B => \arbRegSMCurrentState_0\, C => 
        N_135, D => N_148, Y => N_100_i_0);
    
    \arbRegSMCurrentState[10]\ : SLE
      port map(D => N_104_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_8\);
    
    \arbRegSMCurrentState_RNO[10]\ : CFG4
      generic map(INIT => x"CCC8")

      port map(A => N_120, B => \arbRegSMCurrentState_8\, C => 
        N_135, D => N_148, Y => N_104_i_0);
    
    \arbRegSMCurrentState[14]\ : SLE
      port map(D => \arbRegSMCurrentState_ns_i_i[1]_net_1\, CLK
         => CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_12\);
    
    \arbRegSMCurrentState_ns_i_0_a2_RNILNJC[0]\ : CFG4
      generic map(INIT => x"3022")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        B => \hsel2_i_4\, C => regHADDR_0, D => masterRegAddrSel, 
        Y => N_194_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \arbRegSMCurrentState_ns_i_0_a2[0]\ : CFG4
      generic map(INIT => x"3331")

      port map(A => N_225, B => \arbRegSMCurrentState_13\, C => 
        \N_157_i_i_o2_0_out\, D => N_120, Y => \hsel2_i_4\);
    
    \arbRegSMCurrentState_ns_i_0_a2_RNINPJC[0]\ : CFG4
      generic map(INIT => x"3022")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        B => \hsel2_i_4\, C => regHADDR_2, D => masterRegAddrSel, 
        Y => N_196_i_0);
    
    \arbRegSMCurrentState[15]\ : SLE
      port map(D => N_109_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_13\);
    
    \arbRegSMCurrentState_RNO[15]\ : CFG4
      generic map(INIT => x"888C")

      port map(A => \arbRegSMCurrentState_13\, B => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, C => 
        \N_157_i_i_o2_0\, D => \N_157_i_i_o2_0_out\, Y => 
        N_109_i_0);
    
    \arbRegSMCurrentState_RNO[6]\ : CFG4
      generic map(INIT => x"CCC8")

      port map(A => N_120, B => \arbRegSMCurrentState_4\, C => 
        N_135, D => N_148, Y => N_102_i_0);
    
    \arbRegSMCurrentState[6]\ : SLE
      port map(D => N_102_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_4\);
    
    N_157_i_i_o2_0_s : CFG3
      generic map(INIT => x"BF")

      port map(A => N_148, B => N_138, C => N_149, Y => 
        \N_157_i_i_o2_0_out\);
    
    \arbRegSMCurrentState_ns_i_0_a2_RNI41UH[0]\ : CFG4
      generic map(INIT => x"3022")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        B => \hsel2_i_4\, C => regHADDR_8, D => masterRegAddrSel, 
        Y => CoreAHBLite_0_AHBmslave3_HADDR(11));
    
    hsel2_i_4_i : CFG4
      generic map(INIT => x"CCCE")

      port map(A => N_225, B => \arbRegSMCurrentState_13\, C => 
        \N_157_i_i_o2_0_out\, D => N_120, Y => hsel2_i_4_i_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \arbRegSMCurrentState_ns_i_i[1]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \arbRegSMCurrentState_12\, B => xhdl1221(3), 
        C => N_271, Y => \arbRegSMCurrentState_ns_i_i[1]_net_1\);
    
    \arbRegSMCurrentState[2]\ : SLE
      port map(D => N_100_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState_0\);
    
    \arbRegSMCurrentState_ns_i_0_a2_RNIMOJC[0]\ : CFG4
      generic map(INIT => x"3022")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        B => \hsel2_i_4\, C => regHADDR_1, D => masterRegAddrSel, 
        Y => N_195_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVESTAGE_1 is

    port( masterDataInProg                                          : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA  : in    std_logic_vector(31 downto 0);
          xhdl1221                                                  : in    std_logic_vector(3 to 3);
          CoreAHBLite_0_AHBmslave3_HADDR                            : out   std_logic_vector(11 to 11);
          arbRegSMCurrentState_13                                   : out   std_logic;
          arbRegSMCurrentState_12                                   : out   std_logic;
          arbRegSMCurrentState_8                                    : out   std_logic;
          arbRegSMCurrentState_4                                    : out   std_logic;
          arbRegSMCurrentState_0                                    : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 : in    std_logic;
          regHADDR_8                                                : in    std_logic;
          regHADDR_2                                                : in    std_logic;
          regHADDR_1                                                : in    std_logic;
          regHADDR_0                                                : in    std_logic;
          MSS_READY                                                 : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                      : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                   : in    std_logic;
          N_63_i_0                                                  : out   std_logic;
          N_62_i_0                                                  : out   std_logic;
          N_60_i_0                                                  : out   std_logic;
          N_98_i_0                                                  : out   std_logic;
          N_96_i_0                                                  : out   std_logic;
          N_94_i_0                                                  : out   std_logic;
          N_92_i_0                                                  : out   std_logic;
          N_90_i_0                                                  : out   std_logic;
          N_88_i_0                                                  : out   std_logic;
          N_86_i_0                                                  : out   std_logic;
          N_84_i_0                                                  : out   std_logic;
          N_82_i_0                                                  : out   std_logic;
          N_80_i_0                                                  : out   std_logic;
          N_78_i_0                                                  : out   std_logic;
          N_76_i_0                                                  : out   std_logic;
          N_74_i_0                                                  : out   std_logic;
          N_72_i_0                                                  : out   std_logic;
          N_70_i_0                                                  : out   std_logic;
          N_68_i_0                                                  : out   std_logic;
          N_66_i_0                                                  : out   std_logic;
          N_64_i_0                                                  : out   std_logic;
          N_58_i_0                                                  : out   std_logic;
          N_56_i_0                                                  : out   std_logic;
          N_54_i_0                                                  : out   std_logic;
          N_52_i_0                                                  : out   std_logic;
          N_50_i_0                                                  : out   std_logic;
          N_48_i_0                                                  : out   std_logic;
          N_46_i_0                                                  : out   std_logic;
          N_44_i_0                                                  : out   std_logic;
          N_42_i_0                                                  : out   std_logic;
          N_40_i_0                                                  : out   std_logic;
          N_38_i_0                                                  : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                       : in    std_logic;
          hready_m_xhdl345                                          : in    std_logic;
          un1_SDATASELInt_1                                         : in    std_logic;
          HTRANS_i_a2_0_0                                           : out   std_logic;
          N_271                                                     : in    std_logic;
          N_120                                                     : in    std_logic;
          N_225                                                     : in    std_logic;
          N_157_i_i_o2_0                                            : out   std_logic;
          N_148                                                     : in    std_logic;
          N_138                                                     : in    std_logic;
          N_149                                                     : in    std_logic;
          N_157_i_i_o2_0_out                                        : out   std_logic;
          hsel2_i_4                                                 : out   std_logic;
          N_135                                                     : in    std_logic;
          masterRegAddrSel                                          : in    std_logic;
          N_196_i_0                                                 : out   std_logic;
          N_195_i_0                                                 : out   std_logic;
          N_194_i_0                                                 : out   std_logic
        );

end COREAHBLITE_SLAVESTAGE_1;

architecture DEF_ARCH of COREAHBLITE_SLAVESTAGE_1 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVEARBITER_1
    port( xhdl1221                                                  : in    std_logic_vector(3 to 3) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HADDR                            : out   std_logic_vector(11 to 11);
          arbRegSMCurrentState_13                                   : out   std_logic;
          arbRegSMCurrentState_12                                   : out   std_logic;
          arbRegSMCurrentState_8                                    : out   std_logic;
          arbRegSMCurrentState_4                                    : out   std_logic;
          arbRegSMCurrentState_0                                    : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 : in    std_logic := 'U';
          regHADDR_8                                                : in    std_logic := 'U';
          regHADDR_2                                                : in    std_logic := 'U';
          regHADDR_1                                                : in    std_logic := 'U';
          regHADDR_0                                                : in    std_logic := 'U';
          MSS_READY                                                 : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                      : in    std_logic := 'U';
          N_271                                                     : in    std_logic := 'U';
          N_120                                                     : in    std_logic := 'U';
          N_225                                                     : in    std_logic := 'U';
          N_157_i_i_o2_0                                            : out   std_logic;
          N_148                                                     : in    std_logic := 'U';
          N_138                                                     : in    std_logic := 'U';
          N_149                                                     : in    std_logic := 'U';
          N_157_i_i_o2_0_out                                        : out   std_logic;
          hsel2_i_4                                                 : out   std_logic;
          N_135                                                     : in    std_logic := 'U';
          masterRegAddrSel                                          : in    std_logic := 'U';
          hsel2_i_4_i_0                                             : out   std_logic;
          N_196_i_0                                                 : out   std_logic;
          N_195_i_0                                                 : out   std_logic;
          N_194_i_0                                                 : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                       : in    std_logic := 'U'
        );
  end component;

    signal \masterDataInProg[0]_net_1\, VCC_net_1, hsel2_i_4_i_0, 
        GND_net_1, \arbRegSMCurrentState_13\ : std_logic;

    for all : COREAHBLITE_SLAVEARBITER_1
	Use entity work.COREAHBLITE_SLAVEARBITER_1(DEF_ARCH);
begin 

    masterDataInProg(0) <= \masterDataInProg[0]_net_1\;
    arbRegSMCurrentState_13 <= \arbRegSMCurrentState_13\;

    \masterDataInProg_RNICEPO_6[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        B => \masterDataInProg[0]_net_1\, Y => N_40_i_0);
    
    \masterDataInProg_RNICEPO_8[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        B => \masterDataInProg[0]_net_1\, Y => N_56_i_0);
    
    \masterDataInProg_RNICEPO_23[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        B => \masterDataInProg[0]_net_1\, Y => N_88_i_0);
    
    \masterDataInProg_RNICEPO_17[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        B => \masterDataInProg[0]_net_1\, Y => N_60_i_0);
    
    \masterDataInProg_RNICEPO_15[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        B => \masterDataInProg[0]_net_1\, Y => N_63_i_0);
    
    \masterDataInProg_RNICEPO_12[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        B => \masterDataInProg[0]_net_1\, Y => N_66_i_0);
    
    \masterDataInProg_RNICEPO_20[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        B => \masterDataInProg[0]_net_1\, Y => N_94_i_0);
    
    \masterDataInProg_RNICEPO_24[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        B => \masterDataInProg[0]_net_1\, Y => N_86_i_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \masterDataInProg_RNICEPO_21[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        B => \masterDataInProg[0]_net_1\, Y => N_92_i_0);
    
    \masterDataInProg_RNICEPO[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        B => \masterDataInProg[0]_net_1\, Y => N_54_i_0);
    
    \masterDataInProg_RNICEPO_1[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        B => \masterDataInProg[0]_net_1\, Y => N_50_i_0);
    
    \masterDataInProg_RNICEPO_7[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        B => \masterDataInProg[0]_net_1\, Y => N_38_i_0);
    
    \masterDataInProg_RNICEPO_18[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        B => \masterDataInProg[0]_net_1\, Y => N_98_i_0);
    
    \masterDataInProg_RNICEPO_26[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        B => \masterDataInProg[0]_net_1\, Y => N_82_i_0);
    
    \HTRANS_i_a2_0_0\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \arbRegSMCurrentState_13\, B => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, C => 
        hready_m_xhdl345, D => un1_SDATASELInt_1, Y => 
        HTRANS_i_a2_0_0);
    
    \masterDataInProg_RNICEPO_13[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        B => \masterDataInProg[0]_net_1\, Y => N_64_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \masterDataInProg_RNICEPO_30[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        B => \masterDataInProg[0]_net_1\, Y => N_74_i_0);
    
    \masterDataInProg[0]\ : SLE
      port map(D => hsel2_i_4_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \masterDataInProg[0]_net_1\);
    
    \masterDataInProg_RNICEPO_29[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        B => \masterDataInProg[0]_net_1\, Y => N_76_i_0);
    
    \masterDataInProg_RNICEPO_10[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        B => \masterDataInProg[0]_net_1\, Y => N_70_i_0);
    
    \masterDataInProg_RNICEPO_14[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        B => \masterDataInProg[0]_net_1\, Y => N_58_i_0);
    
    \masterDataInProg_RNICEPO_3[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        B => \masterDataInProg[0]_net_1\, Y => N_46_i_0);
    
    \masterDataInProg_RNICEPO_11[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        B => \masterDataInProg[0]_net_1\, Y => N_68_i_0);
    
    \masterDataInProg_RNICEPO_9[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        B => \masterDataInProg[0]_net_1\, Y => N_72_i_0);
    
    \masterDataInProg_RNICEPO_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        B => \masterDataInProg[0]_net_1\, Y => N_44_i_0);
    
    \masterDataInProg_RNICEPO_27[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        B => \masterDataInProg[0]_net_1\, Y => N_80_i_0);
    
    \masterDataInProg_RNICEPO_25[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        B => \masterDataInProg[0]_net_1\, Y => N_84_i_0);
    
    \masterDataInProg_RNICEPO_22[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        B => \masterDataInProg[0]_net_1\, Y => N_90_i_0);
    
    slave_arbiter : COREAHBLITE_SLAVEARBITER_1
      port map(xhdl1221(3) => xhdl1221(3), 
        CoreAHBLite_0_AHBmslave3_HADDR(11) => 
        CoreAHBLite_0_AHBmslave3_HADDR(11), 
        arbRegSMCurrentState_13 => \arbRegSMCurrentState_13\, 
        arbRegSMCurrentState_12 => arbRegSMCurrentState_12, 
        arbRegSMCurrentState_8 => arbRegSMCurrentState_8, 
        arbRegSMCurrentState_4 => arbRegSMCurrentState_4, 
        arbRegSMCurrentState_0 => arbRegSMCurrentState_0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        regHADDR_8 => regHADDR_8, regHADDR_2 => regHADDR_2, 
        regHADDR_1 => regHADDR_1, regHADDR_0 => regHADDR_0, 
        MSS_READY => MSS_READY, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, N_271 => N_271, 
        N_120 => N_120, N_225 => N_225, N_157_i_i_o2_0 => 
        N_157_i_i_o2_0, N_148 => N_148, N_138 => N_138, N_149 => 
        N_149, N_157_i_i_o2_0_out => N_157_i_i_o2_0_out, 
        hsel2_i_4 => hsel2_i_4, N_135 => N_135, masterRegAddrSel
         => masterRegAddrSel, hsel2_i_4_i_0 => hsel2_i_4_i_0, 
        N_196_i_0 => N_196_i_0, N_195_i_0 => N_195_i_0, N_194_i_0
         => N_194_i_0, CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1);
    
    \masterDataInProg_RNICEPO_0[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        B => \masterDataInProg[0]_net_1\, Y => N_52_i_0);
    
    \masterDataInProg_RNICEPO_2[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        B => \masterDataInProg[0]_net_1\, Y => N_48_i_0);
    
    \masterDataInProg_RNICEPO_16[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        B => \masterDataInProg[0]_net_1\, Y => N_62_i_0);
    
    \masterDataInProg_RNICEPO_19[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        B => \masterDataInProg[0]_net_1\, Y => N_96_i_0);
    
    \masterDataInProg_RNICEPO_5[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        B => \masterDataInProg[0]_net_1\, Y => N_42_i_0);
    
    \masterDataInProg_RNICEPO_28[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        B => \masterDataInProg[0]_net_1\, Y => N_78_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_DEFAULTSLAVESM_0 is

    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP : in    std_logic_vector(0 to 0);
          MSS_READY                                               : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                    : in    std_logic;
          defSlaveSMNextState                                     : out   std_logic;
          N_321                                                   : in    std_logic;
          N_126                                                   : in    std_logic;
          hready_m_xhdl345                                        : in    std_logic;
          N_129                                                   : out   std_logic
        );

end COREAHBLITE_DEFAULTSLAVESM_0;

architecture DEF_ARCH of COREAHBLITE_DEFAULTSLAVESM_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal \defSlaveSMCurrentState\, VCC_net_1, 
        defSlaveSMNextState_net_1, GND_net_1 : std_logic;

begin 

    defSlaveSMNextState <= defSlaveSMNextState_net_1;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    defSlaveSMNextState_RNICC2O3 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_126, B => defSlaveSMNextState_net_1, C => 
        hready_m_xhdl345, D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        Y => N_129);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \defSlaveSMNextState\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_321, B => \defSlaveSMCurrentState\, Y => 
        defSlaveSMNextState_net_1);
    
    defSlaveSMCurrentState : SLE
      port map(D => defSlaveSMNextState_net_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \defSlaveSMCurrentState\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MASTERSTAGE_1_1_0_40_0 is

    port( xhdl1221                                                    : out   std_logic_vector(3 to 3);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE     : in    std_logic_vector(1 downto 0);
          masterDataInProg                                            : in    std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS    : in    std_logic_vector(1 to 1);
          result_addr_net_0                                           : in    std_logic_vector(3 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP     : out   std_logic_vector(0 to 0);
          masterDataInProg_0                                          : in    std_logic_vector(0 to 0);
          CoreAHBLite_0_AHBmslave3_HRDATA                             : in    std_logic_vector(31 downto 0);
          line_7                                                      : in    std_logic_vector(2 downto 1);
          arbRegSMCurrentState_ns_i_0                                 : in    std_logic_vector(1 to 1);
          xhdl1222_0                                                  : out   std_logic;
          xhdl1222_2                                                  : out   std_logic;
          SDATASELInt_0                                               : out   std_logic;
          SDATASELInt_1                                               : out   std_logic;
          SDATASELInt_2                                               : out   std_logic;
          SDATASELInt_4                                               : out   std_logic;
          SDATASELInt_6                                               : out   std_logic;
          SDATASELInt_7                                               : out   std_logic;
          SDATASELInt_8                                               : out   std_logic;
          SDATASELInt_9                                               : out   std_logic;
          SDATASELInt_10                                              : out   std_logic;
          SDATASELInt_11                                              : out   std_logic;
          SDATASELInt_12                                              : out   std_logic;
          SDATASELInt_13                                              : out   std_logic;
          regHADDR_11                                                 : out   std_logic;
          regHADDR_3                                                  : out   std_logic;
          regHADDR_4                                                  : out   std_logic;
          regHADDR_5                                                  : out   std_logic;
          arbRegSMCurrentState_13                                     : in    std_logic;
          arbRegSMCurrentState_12                                     : in    std_logic;
          arbRegSMCurrentState_8                                      : in    std_logic;
          arbRegSMCurrentState_4                                      : in    std_logic;
          arbRegSMCurrentState_0                                      : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31  : in    std_logic;
          line_13                                                     : in    std_logic;
          line_10                                                     : in    std_logic;
          line_21                                                     : in    std_logic;
          line_24                                                     : in    std_logic;
          line_18                                                     : in    std_logic;
          line_23                                                     : in    std_logic;
          line_16                                                     : in    std_logic;
          line_28                                                     : in    std_logic;
          line_9                                                      : in    std_logic;
          line_3_d0                                                   : in    std_logic;
          line_5_d0                                                   : in    std_logic;
          line_15                                                     : in    std_logic;
          line_26                                                     : in    std_logic;
          line_14                                                     : in    std_logic;
          line_20                                                     : in    std_logic;
          line_2_d0                                                   : in    std_logic;
          line_25                                                     : in    std_logic;
          line_29                                                     : in    std_logic;
          line_19                                                     : in    std_logic;
          line_27                                                     : in    std_logic;
          line_30                                                     : in    std_logic;
          line_17                                                     : in    std_logic;
          line_8                                                      : in    std_logic;
          line_0_d0                                                   : in    std_logic;
          line_6_d0                                                   : in    std_logic;
          line_1_d0                                                   : in    std_logic;
          line_0_10                                                   : in    std_logic;
          line_0_21                                                   : in    std_logic;
          line_0_24                                                   : in    std_logic;
          line_0_18                                                   : in    std_logic;
          line_0_23                                                   : in    std_logic;
          line_0_16                                                   : in    std_logic;
          line_0_28                                                   : in    std_logic;
          line_0_9                                                    : in    std_logic;
          line_0_3                                                    : in    std_logic;
          line_0_5                                                    : in    std_logic;
          line_0_15                                                   : in    std_logic;
          line_0_26                                                   : in    std_logic;
          line_0_14                                                   : in    std_logic;
          line_0_20                                                   : in    std_logic;
          line_0_2                                                    : in    std_logic;
          line_0_25                                                   : in    std_logic;
          line_0_29                                                   : in    std_logic;
          line_0_19                                                   : in    std_logic;
          line_0_27                                                   : in    std_logic;
          line_0_30                                                   : in    std_logic;
          line_0_17                                                   : in    std_logic;
          line_0_8                                                    : in    std_logic;
          line_0_0                                                    : in    std_logic;
          line_0_1                                                    : in    std_logic;
          line_0_6                                                    : in    std_logic;
          line_0_13                                                   : in    std_logic;
          line_1_10                                                   : in    std_logic;
          line_1_21                                                   : in    std_logic;
          line_1_24                                                   : in    std_logic;
          line_1_18                                                   : in    std_logic;
          line_1_23                                                   : in    std_logic;
          line_1_16                                                   : in    std_logic;
          line_1_28                                                   : in    std_logic;
          line_1_9                                                    : in    std_logic;
          line_1_3                                                    : in    std_logic;
          line_1_5                                                    : in    std_logic;
          line_1_15                                                   : in    std_logic;
          line_1_26                                                   : in    std_logic;
          line_1_14                                                   : in    std_logic;
          line_1_20                                                   : in    std_logic;
          line_1_2                                                    : in    std_logic;
          line_1_25                                                   : in    std_logic;
          line_1_29                                                   : in    std_logic;
          line_1_19                                                   : in    std_logic;
          line_1_27                                                   : in    std_logic;
          line_1_30                                                   : in    std_logic;
          line_1_17                                                   : in    std_logic;
          line_1_8                                                    : in    std_logic;
          line_1_0                                                    : in    std_logic;
          line_1_1                                                    : in    std_logic;
          line_1_6                                                    : in    std_logic;
          line_1_13                                                   : in    std_logic;
          line_2_19                                                   : in    std_logic;
          line_2_27                                                   : in    std_logic;
          line_2_30                                                   : in    std_logic;
          line_2_17                                                   : in    std_logic;
          line_2_8                                                    : in    std_logic;
          line_2_10                                                   : in    std_logic;
          line_2_15                                                   : in    std_logic;
          line_2_26                                                   : in    std_logic;
          line_2_20                                                   : in    std_logic;
          line_2_0                                                    : in    std_logic;
          line_2_1                                                    : in    std_logic;
          line_2_29                                                   : in    std_logic;
          line_2_25                                                   : in    std_logic;
          line_2_2                                                    : in    std_logic;
          line_2_6                                                    : in    std_logic;
          line_2_13                                                   : in    std_logic;
          line_2_14                                                   : in    std_logic;
          line_2_5                                                    : in    std_logic;
          line_2_3                                                    : in    std_logic;
          line_2_9                                                    : in    std_logic;
          line_2_28                                                   : in    std_logic;
          line_2_16                                                   : in    std_logic;
          line_2_23                                                   : in    std_logic;
          line_2_18                                                   : in    std_logic;
          line_2_24                                                   : in    std_logic;
          line_2_21                                                   : in    std_logic;
          line_3_19                                                   : in    std_logic;
          line_3_17                                                   : in    std_logic;
          line_3_8                                                    : in    std_logic;
          line_3_0                                                    : in    std_logic;
          line_3_1                                                    : in    std_logic;
          line_3_29                                                   : in    std_logic;
          line_3_25                                                   : in    std_logic;
          line_3_2                                                    : in    std_logic;
          line_3_20                                                   : in    std_logic;
          line_3_6                                                    : in    std_logic;
          line_3_13                                                   : in    std_logic;
          line_3_14                                                   : in    std_logic;
          line_3_26                                                   : in    std_logic;
          line_3_15                                                   : in    std_logic;
          line_3_5                                                    : in    std_logic;
          line_3_3                                                    : in    std_logic;
          line_3_9                                                    : in    std_logic;
          line_3_28                                                   : in    std_logic;
          line_3_16                                                   : in    std_logic;
          line_3_23                                                   : in    std_logic;
          line_3_18                                                   : in    std_logic;
          line_3_24                                                   : in    std_logic;
          line_3_21                                                   : in    std_logic;
          line_3_10                                                   : in    std_logic;
          SHA256_Module_0_data_out_5                                  : in    std_logic;
          SHA256_Module_0_data_out_13                                 : in    std_logic;
          SHA256_Module_0_data_out_12                                 : in    std_logic;
          SHA256_Module_0_data_out_8                                  : in    std_logic;
          SHA256_Module_0_data_out_23                                 : in    std_logic;
          SHA256_Module_0_data_out_0                                  : in    std_logic;
          line_4_19                                                   : in    std_logic;
          line_4_17                                                   : in    std_logic;
          line_4_8                                                    : in    std_logic;
          line_4_0                                                    : in    std_logic;
          line_4_1                                                    : in    std_logic;
          line_4_29                                                   : in    std_logic;
          line_4_25                                                   : in    std_logic;
          line_4_2                                                    : in    std_logic;
          line_4_20                                                   : in    std_logic;
          line_4_14                                                   : in    std_logic;
          line_4_26                                                   : in    std_logic;
          line_4_15                                                   : in    std_logic;
          line_4_5                                                    : in    std_logic;
          line_4_3                                                    : in    std_logic;
          line_4_9                                                    : in    std_logic;
          line_4_28                                                   : in    std_logic;
          line_4_16                                                   : in    std_logic;
          line_4_23                                                   : in    std_logic;
          line_4_18                                                   : in    std_logic;
          line_4_24                                                   : in    std_logic;
          line_4_21                                                   : in    std_logic;
          line_4_10                                                   : in    std_logic;
          line_4_6                                                    : in    std_logic;
          line_4_13                                                   : in    std_logic;
          line_5_19                                                   : in    std_logic;
          line_5_17                                                   : in    std_logic;
          line_5_8                                                    : in    std_logic;
          line_5_0                                                    : in    std_logic;
          line_5_1                                                    : in    std_logic;
          line_5_29                                                   : in    std_logic;
          line_5_25                                                   : in    std_logic;
          line_5_2                                                    : in    std_logic;
          line_5_20                                                   : in    std_logic;
          line_5_6                                                    : in    std_logic;
          line_5_13                                                   : in    std_logic;
          line_5_14                                                   : in    std_logic;
          line_5_26                                                   : in    std_logic;
          line_5_15                                                   : in    std_logic;
          line_5_5                                                    : in    std_logic;
          line_5_3                                                    : in    std_logic;
          line_5_9                                                    : in    std_logic;
          line_5_28                                                   : in    std_logic;
          line_5_16                                                   : in    std_logic;
          line_5_23                                                   : in    std_logic;
          line_5_18                                                   : in    std_logic;
          line_5_24                                                   : in    std_logic;
          line_5_21                                                   : in    std_logic;
          line_5_10                                                   : in    std_logic;
          line_6_19                                                   : in    std_logic;
          line_6_17                                                   : in    std_logic;
          line_6_8                                                    : in    std_logic;
          line_6_0                                                    : in    std_logic;
          line_6_1                                                    : in    std_logic;
          line_6_29                                                   : in    std_logic;
          line_6_25                                                   : in    std_logic;
          line_6_2                                                    : in    std_logic;
          line_6_20                                                   : in    std_logic;
          line_6_6                                                    : in    std_logic;
          line_6_13                                                   : in    std_logic;
          line_6_14                                                   : in    std_logic;
          line_6_26                                                   : in    std_logic;
          line_6_15                                                   : in    std_logic;
          line_6_5                                                    : in    std_logic;
          line_6_3                                                    : in    std_logic;
          line_6_9                                                    : in    std_logic;
          line_6_28                                                   : in    std_logic;
          line_6_16                                                   : in    std_logic;
          line_6_23                                                   : in    std_logic;
          line_6_18                                                   : in    std_logic;
          line_6_24                                                   : in    std_logic;
          line_6_21                                                   : in    std_logic;
          line_6_10                                                   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11 : out   std_logic;
          MSS_READY                                                   : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                        : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE    : in    std_logic;
          masterRegAddrSel                                            : out   std_logic;
          N_138                                                       : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                         : in    std_logic;
          N_148                                                       : out   std_logic;
          N_135                                                       : out   std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY                  : in    std_logic;
          hready_m_xhdl344_7                                          : out   std_logic;
          N_225                                                       : out   std_logic;
          N_149                                                       : out   std_logic;
          N_276                                                       : out   std_logic;
          N_259                                                       : out   std_logic;
          N_243                                                       : out   std_logic;
          N_236                                                       : out   std_logic;
          N_235                                                       : out   std_logic;
          N_277                                                       : out   std_logic;
          N_255                                                       : out   std_logic;
          N_241                                                       : out   std_logic;
          N_242                                                       : out   std_logic;
          N_244                                                       : out   std_logic;
          N_246                                                       : out   std_logic;
          N_247                                                       : out   std_logic;
          N_256                                                       : out   std_logic;
          N_257                                                       : out   std_logic;
          N_258                                                       : out   std_logic;
          ren_pos                                                     : in    std_logic;
          hready_m_xhdl343_10                                         : out   std_logic;
          hready_m_xhdl343_11                                         : out   std_logic;
          N_120                                                       : out   std_logic;
          N_127                                                       : out   std_logic;
          N_216                                                       : in    std_logic;
          N_215                                                       : in    std_logic;
          hready_m_xhdl345                                            : out   std_logic;
          un1_SDATASELInt_1                                           : out   std_logic;
          N_335                                                       : in    std_logic;
          N_214                                                       : in    std_logic;
          N_305                                                       : in    std_logic;
          N_206                                                       : out   std_logic;
          N_508                                                       : in    std_logic;
          N_478_i_0                                                   : out   std_logic;
          N_507                                                       : in    std_logic;
          N_477_i_0                                                   : out   std_logic;
          N_479_i_0                                                   : out   std_logic;
          N_480_i_0                                                   : out   std_logic;
          N_481_i_0                                                   : out   std_logic;
          un8_hreadyin_i_0                                            : in    std_logic;
          N_9_i_0                                                     : out   std_logic;
          N_226                                                       : in    std_logic;
          defSlaveSMNextState                                         : out   std_logic
        );

end COREAHBLITE_MASTERSTAGE_1_1_0_40_0;

architecture DEF_ARCH of COREAHBLITE_MASTERSTAGE_1_1_0_40_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component COREAHBLITE_DEFAULTSLAVESM_0
    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP : in    std_logic_vector(0 to 0) := (others => 'U');
          MSS_READY                                               : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                    : in    std_logic := 'U';
          defSlaveSMNextState                                     : out   std_logic;
          N_321                                                   : in    std_logic := 'U';
          N_126                                                   : in    std_logic := 'U';
          hready_m_xhdl345                                        : in    std_logic := 'U';
          N_129                                                   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \SDATASELInt[15]_net_1\, VCC_net_1, N_61_i_0, 
        N_27_i_0, GND_net_1, \SDATASELInt_0\, N_35_i_0, 
        \SDATASELInt_1\, N_37_i_0, \SDATASELInt_2\, N_39_i_0, 
        \xhdl1222_0\, \xhdl1221[3]\, \SDATASELInt_4\, N_41_i_0, 
        \xhdl1222_2\, N_249_i_0, \SDATASELInt_6\, N_43_i_0, 
        \SDATASELInt_7\, N_45_i_1, \SDATASELInt_8\, N_47_i_0, 
        \SDATASELInt_9\, N_49_i_0, \SDATASELInt_10\, N_51_i_0, 
        \SDATASELInt_11\, N_53_i_0, \SDATASELInt_12\, N_55_i_0, 
        \SDATASELInt_13\, N_57_i_1, \SDATASELInt[14]_net_1\, 
        N_59_i_0, N_106_i_0, \regHADDR[12]_net_1\, 
        \regHADDR[13]_net_1\, \regHADDR[14]_net_1\, 
        \regHADDR[15]_net_1\, \regHADDR[29]_net_1\, 
        \regHADDR[30]_net_1\, \regHSIZE[0]_net_1\, 
        \regHSIZE[1]_net_1\, \regHADDR[0]_net_1\, 
        \regHADDR[1]_net_1\, \regHADDR[2]_net_1\, 
        \regHADDR[6]_net_1\, \regHADDR[7]_net_1\, 
        \regHADDR[8]_net_1\, \regHADDR[9]_net_1\, 
        \regHADDR[10]_net_1\, \regHWRITE\, \regHTRANS\, 
        masterRegAddrSel_net_1, N_108_i_0, \N_138\, \N_148\, 
        N_178, N_737, N_550, N_742, \HRDATA_1_4_1[11]_net_1\, 
        \HRDATA_1_4[11]_net_1\, N_740, N_739, 
        \HRDATA_1_4_1[22]_net_1\, \HRDATA_1_4[22]_net_1\, 
        \HRDATA_1_4_1[25]_net_1\, \HRDATA_1_4[25]_net_1\, 
        \HRDATA_1_4_1[19]_net_1\, \HRDATA_1_4[19]_net_1\, 
        \HRDATA_1_4_1[24]_net_1\, \HRDATA_1_4[24]_net_1\, 
        \HRDATA_1_4_1[17]_net_1\, \HRDATA_1_4[17]_net_1\, 
        \HRDATA_1_4_1[29]_net_1\, \HRDATA_1_4[29]_net_1\, 
        \HRDATA_1_4_1[10]_net_1\, \HRDATA_1_4[10]_net_1\, 
        \HRDATA_1_4_1[4]_net_1\, \HRDATA_1_4[4]_net_1\, 
        \HRDATA_1_4_1[6]_net_1\, \HRDATA_1_4[6]_net_1\, 
        \HRDATA_1_4_1[16]_net_1\, \HRDATA_1_4[16]_net_1\, 
        \HRDATA_1_4_1[27]_net_1\, \HRDATA_1_4[27]_net_1\, 
        \HRDATA_1_4_1[15]_net_1\, \HRDATA_1_4[15]_net_1\, 
        \HRDATA_1_4_1[21]_net_1\, \HRDATA_1_4[21]_net_1\, 
        \HRDATA_1_4_1[3]_net_1\, \HRDATA_1_4[3]_net_1\, 
        \HRDATA_1_4_1[26]_net_1\, \HRDATA_1_4[26]_net_1\, 
        \HRDATA_1_4_1[30]_net_1\, \HRDATA_1_4[30]_net_1\, 
        \HRDATA_1_m5_0_i_m3_1_1[20]\, N_511, 
        \HRDATA_i_m3_1_1[28]\, N_501, 
        \HRDATA_1_m5_i_m3_1_1[20]_net_1\, N_514, 
        \HRDATA_i_m3_1_1[31]\, N_502, 
        \HRDATA_1_m5_0_i_m3_1_1[18]\, N_517, 
        \HRDATA_1_m5_i_m3_1_1[9]_net_1\, N_264, 
        \HRDATA_1_m5_i_m3_1_1[18]_net_1\, N_520, 
        \HRDATA_1_m5_0_i_m3_1_1[9]\, N_523, \N_135\, N_144, N_738, 
        N_741, N_126, N_320, \hready_m_xhdl344_7\, \N_225\, 
        \N_149\, \HRDATA_1_a3_7_0[11]_net_1\, 
        \HRDATA_1_a3_17_0[11]_net_1\, N_318, N_681, 
        \hready_m_xhdl343_10\, \hready_m_xhdl343_11\, 
        \SADDRSEL_i_0[8]\, \SADDRSEL_i_0[4]\, N_142_i, N_146, 
        \N_120\, N_143, N_151, un1_hready_m_xhdl343_1_i_0_a2_1, 
        N_321, N_249, un1_hready_m_xhdl343_1_i_0_o2_1_tz, 
        \hready_m_xhdl345\, \un1_SDATASELInt_1\, N_602, N_436, 
        N_733, N_485, N_755, un1_hready_m_xhdl343_1_i_0_o2_0, 
        N_750, N_298, N_308, N_555, N_572, N_582, N_592, N_415, 
        N_425, N_439, N_449, N_469, N_607, N_617, N_627, N_637, 
        N_647, N_657, N_667, N_678, N_687, N_751, N_757, N_758, 
        \N_206\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        \HRDATA_i_1[31]_net_1\, \HRDATA_1_i_1[18]_net_1\, 
        \HRDATA_1_i_1[9]_net_1\, \HRDATA_1_i_1[20]_net_1\, 
        \HRDATA_i_1[28]_net_1\, \d_masterRegAddrSel_i_o2_0\, 
        N_536, N_543, N_556, N_558, N_559, N_564, N_587, N_461, 
        N_629, N_631, N_632, N_746, N_748, N_207, 
        \HRDATA_1_2[1]_net_1\, \HRDATA_1_1[1]_net_1\, 
        \HRDATA_1_0[1]_net_1\, \HRDATA_1_2[2]_net_1\, 
        \HRDATA_1_1[2]_net_1\, \HRDATA_1_0[2]_net_1\, 
        \HRDATA_1_1[30]_net_1\, \HRDATA_1_0[30]_net_1\, 
        \HRDATA_1_1[26]_net_1\, \HRDATA_1_0[26]_net_1\, 
        \HRDATA_1_1[3]_net_1\, \HRDATA_1_0[3]_net_1\, 
        \HRDATA_1_1[21]_net_1\, \HRDATA_1_0[21]_net_1\, 
        \HRDATA_1_2[7]_net_1\, \HRDATA_1_1[7]_net_1\, 
        \HRDATA_1_0[7]_net_1\, \HRDATA_1_2[14]_net_1\, 
        \HRDATA_1_1[14]_net_1\, \HRDATA_1_0[14]_net_1\, 
        \HRDATA_1_1[15]_net_1\, \HRDATA_1_0[15]_net_1\, 
        \HRDATA_1_1[27]_net_1\, \HRDATA_1_0[27]_net_1\, 
        \HRDATA_1_1[16]_net_1\, \HRDATA_1_0[16]_net_1\, 
        \HRDATA_1_1[6]_net_1\, \HRDATA_1_0[6]_net_1\, 
        \HRDATA_1_1[4]_net_1\, \HRDATA_1_0[4]_net_1\, 
        \HRDATA_1_1[10]_net_1\, \HRDATA_1_0[10]_net_1\, 
        \HRDATA_1_1[29]_net_1\, \HRDATA_1_0[29]_net_1\, 
        \HRDATA_1_1[17]_net_1\, \HRDATA_1_0[17]_net_1\, 
        \HRDATA_1_1[24]_net_1\, \HRDATA_1_0[24]_net_1\, 
        \HRDATA_1_1[19]_net_1\, \HRDATA_1_0[19]_net_1\, 
        \HRDATA_1_1[25]_net_1\, \HRDATA_1_0[25]_net_1\, 
        \HRDATA_1_1[22]_net_1\, \HRDATA_1_0[22]_net_1\, 
        \HRDATA_1_1[11]_net_1\, \HRDATA_1_0[11]_net_1\, 
        \HRDATA_1_5[1]_net_1\, \HRDATA_1_5[2]_net_1\, 
        \HRDATA_1_5[30]_net_1\, \HRDATA_1_5[26]_net_1\, 
        \HRDATA_1_5[3]_net_1\, \HRDATA_1_5[21]_net_1\, 
        \HRDATA_1_5[7]_net_1\, \HRDATA_1_4[7]_net_1\, 
        \HRDATA_1_5[14]_net_1\, \HRDATA_1_4[14]_net_1\, 
        \HRDATA_1_5[15]_net_1\, \HRDATA_1_5[27]_net_1\, 
        \HRDATA_1_5[16]_net_1\, \HRDATA_1_5[6]_net_1\, 
        \HRDATA_1_5[4]_net_1\, \HRDATA_1_5[10]_net_1\, 
        \HRDATA_1_5[29]_net_1\, \HRDATA_1_5[17]_net_1\, 
        \HRDATA_1_5[24]_net_1\, \HRDATA_1_5[19]_net_1\, 
        \HRDATA_1_5[25]_net_1\, \HRDATA_1_5[22]_net_1\, 
        \HRDATA_1_5[11]_net_1\, N_129, 
        \masterAddrClockEnable_i_2\, \HRDATA_1_6[1]_net_1\, 
        \HRDATA_1_6[2]_net_1\, \d_masterRegAddrSel_i_0\, 
        \masterAddrClockEnable_i_5\ : std_logic;

    for all : COREAHBLITE_DEFAULTSLAVESM_0
	Use entity work.COREAHBLITE_DEFAULTSLAVESM_0(DEF_ARCH);
begin 

    xhdl1221(3) <= \xhdl1221[3]\;
    CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0) <= 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\;
    xhdl1222_0 <= \xhdl1222_0\;
    xhdl1222_2 <= \xhdl1222_2\;
    SDATASELInt_0 <= \SDATASELInt_0\;
    SDATASELInt_1 <= \SDATASELInt_1\;
    SDATASELInt_2 <= \SDATASELInt_2\;
    SDATASELInt_4 <= \SDATASELInt_4\;
    SDATASELInt_6 <= \SDATASELInt_6\;
    SDATASELInt_7 <= \SDATASELInt_7\;
    SDATASELInt_8 <= \SDATASELInt_8\;
    SDATASELInt_9 <= \SDATASELInt_9\;
    SDATASELInt_10 <= \SDATASELInt_10\;
    SDATASELInt_11 <= \SDATASELInt_11\;
    SDATASELInt_12 <= \SDATASELInt_12\;
    SDATASELInt_13 <= \SDATASELInt_13\;
    masterRegAddrSel <= masterRegAddrSel_net_1;
    N_138 <= \N_138\;
    N_148 <= \N_148\;
    N_135 <= \N_135\;
    hready_m_xhdl344_7 <= \hready_m_xhdl344_7\;
    N_225 <= \N_225\;
    N_149 <= \N_149\;
    hready_m_xhdl343_10 <= \hready_m_xhdl343_10\;
    hready_m_xhdl343_11 <= \hready_m_xhdl343_11\;
    N_120 <= \N_120\;
    hready_m_xhdl345 <= \hready_m_xhdl345\;
    un1_SDATASELInt_1 <= \un1_SDATASELInt_1\;
    N_206 <= \N_206\;

    \SADDRSEL_i_o2[1]\ : CFG4
      generic map(INIT => x"7277")

      port map(A => masterRegAddrSel_net_1, B => \regHTRANS\, C
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        Y => \N_120\);
    
    hready_m_xhdl345_0_a2_0 : CFG2
      generic map(INIT => x"2")

      port map(A => \xhdl1222_2\, B => \xhdl1222_0\, Y => N_320);
    
    \HRDATA_1_a2_4[14]\ : CFG4
      generic map(INIT => x"0040")

      port map(A => result_addr_net_0(2), B => N_737, C => 
        line_13, D => result_addr_net_0(1), Y => N_550);
    
    \HRDATA_1_i_a2_0[9]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => N_523, B => N_321, C => result_addr_net_0(0), 
        D => N_320, Y => N_687);
    
    \regHADDR[30]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[30]_net_1\);
    
    \HRDATA_1_a3_7_0[11]\ : CFG3
      generic map(INIT => x"10")

      port map(A => result_addr_net_0(2), B => 
        result_addr_net_0(3), C => result_addr_net_0(1), Y => 
        \HRDATA_1_a3_7_0[11]_net_1\);
    
    \HRDATA_1_2[14]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => line_0_13, B => N_740, C => N_737, D => N_550, 
        Y => \HRDATA_1_2[14]_net_1\);
    
    \HRDATA_1_1[17]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_16, B => line_3_16, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[17]_net_1\);
    
    hready_m_xhdl343_1_0_0_a2_0_RNIRFT71 : CFG4
      generic map(INIT => x"1000")

      port map(A => \xhdl1222_0\, B => \xhdl1222_2\, C => N_216, 
        D => N_318, Y => un1_hready_m_xhdl343_1_i_0_a2_1);
    
    \HRDATA_1_5[15]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_14, B => line_6_14, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[15]_net_1\);
    
    \HRDATA_1_0[7]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_3_6, C => N_737, D => N_582, 
        Y => \HRDATA_1_0[7]_net_1\);
    
    hready_m_xhdl340_11_0_a2_0_a2 : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt_13\, B => \SDATASELInt_12\, C
         => \SDATASELInt_11\, D => \SDATASELInt_10\, Y => 
        \hready_m_xhdl343_11\);
    
    \SDATASELInt[7]\ : SLE
      port map(D => N_45_i_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_7\);
    
    \HRDATA_1_1[11]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_3_10, B => line_4_10, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[11]_net_1\);
    
    \SDATASELInt_RNIBDNP[14]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \SDATASELInt[14]_net_1\, B => 
        \SDATASELInt[15]_net_1\, Y => \hready_m_xhdl344_7\);
    
    \HRDATA_1_1[19]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_18, B => line_3_18, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[19]_net_1\);
    
    \HRDATA_1_a2_1[2]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_1_d0, B => N_738, C => N_737, Y => N_629);
    
    \regHADDR[15]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[15]_net_1\);
    
    \GATEDHSIZE_i_m2[0]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHSIZE[0]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0), 
        Y => N_236);
    
    \HRDATA_1_0[24]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_23, C => N_737, D => N_449, 
        Y => \HRDATA_1_0[24]_net_1\);
    
    \HRDATA_1_a2[24]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(24), C => N_321, D => 
        \xhdl1222_2\, Y => N_449);
    
    \HRDATA_1_a3_8[11]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => N_741, B => result_addr_net_0(0), C => N_321, 
        D => \HRDATA_1_a3_17_0[11]_net_1\, Y => N_751);
    
    \PREGATEDHADDR_i_m2[14]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[14]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14, 
        Y => N_242);
    
    masterRegAddrSel_RNO : CFG4
      generic map(INIT => x"0A0E")

      port map(A => \d_masterRegAddrSel_i_o2_0\, B => 
        arbRegSMCurrentState_ns_i_0(1), C => 
        \d_masterRegAddrSel_i_0\, D => N_249, Y => N_108_i_0);
    
    \HRDATA_i_1_RNO[31]\ : CFG4
      generic map(INIT => x"46CE")

      port map(A => result_addr_net_0(1), B => 
        \HRDATA_i_m3_1_1[31]\, C => line_30, D => line_0_30, Y
         => N_502);
    
    \HRDATA_1[30]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[30]_net_1\, B => 
        \HRDATA_1_1[30]_net_1\, C => \HRDATA_1_4[30]_net_1\, D
         => \HRDATA_1_5[30]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30);
    
    \HRDATA_1_5[6]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_5, B => line_6_5, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[6]_net_1\);
    
    \HRDATA_1_4_1[22]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_21, B => line_1_21, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[22]_net_1\);
    
    \HRDATA_1[25]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[25]_net_1\, B => 
        \HRDATA_1_1[25]_net_1\, C => \HRDATA_1_4[25]_net_1\, D
         => \HRDATA_1_5[25]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25);
    
    \HRDATA_1[15]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[15]_net_1\, B => 
        \HRDATA_1_1[15]_net_1\, C => \HRDATA_1_4[15]_net_1\, D
         => \HRDATA_1_5[15]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15);
    
    \HRDATA_1_1[25]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_24, B => line_3_24, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[25]_net_1\);
    
    \SDATASELInt[13]\ : SLE
      port map(D => N_57_i_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_13\);
    
    \regHSIZE[0]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0), 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHSIZE[0]_net_1\);
    
    default_slave_sm : COREAHBLITE_DEFAULTSLAVESM_0
      port map(
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        MSS_READY => MSS_READY, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, defSlaveSMNextState
         => defSlaveSMNextState, N_321 => N_321, N_126 => N_126, 
        hready_m_xhdl345 => \hready_m_xhdl345\, N_129 => N_129);
    
    \HRDATA_1_4_1[16]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_15, B => line_1_15, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[16]_net_1\);
    
    \HRDATA_1_a3_13[11]\ : CFG2
      generic map(INIT => x"1")

      port map(A => result_addr_net_0(2), B => 
        result_addr_net_0(1), Y => N_739);
    
    \HRDATA_1_a2[10]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(10), C => N_321, D => 
        \xhdl1222_2\, Y => N_657);
    
    \HRDATA_i_1[31]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_755, B => N_502, C => N_485, D => N_602, Y
         => \HRDATA_i_1[31]_net_1\);
    
    \HRDATA_1_a3_3[11]\ : CFG3
      generic map(INIT => x"40")

      port map(A => result_addr_net_0(3), B => N_738, C => N_733, 
        Y => N_746);
    
    \SDATASELInt_RNO[9]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \N_149\, B => \N_148\, C => N_146, D => 
        \N_225\, Y => N_49_i_0);
    
    \HRDATA_1_4_1[29]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_28, B => line_1_28, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[29]_net_1\);
    
    \HRDATA_1_0[3]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_2, C => N_737, D => N_667, 
        Y => \HRDATA_1_0[3]_net_1\);
    
    \HRDATA_1_1[16]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => line_3_15, B => N_750, C => N_543, Y => 
        \HRDATA_1_1[16]_net_1\);
    
    \HRDATA_i_1[28]\ : CFG4
      generic map(INIT => x"B100")

      port map(A => result_addr_net_0(0), B => N_508, C => N_501, 
        D => \hready_m_xhdl345\, Y => \HRDATA_i_1[28]_net_1\);
    
    \HRDATA_1_a2[15]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(15), C => N_321, D => 
        \xhdl1222_2\, Y => N_617);
    
    \HRDATA_1_4_1[24]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_23, B => line_1_23, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[24]_net_1\);
    
    \HRDATA[13]\ : CFG4
      generic map(INIT => x"88C0")

      port map(A => SHA256_Module_0_data_out_13, B => 
        \un1_SDATASELInt_1\, C => 
        CoreAHBLite_0_AHBmslave3_HRDATA(13), D => \xhdl1222_2\, Y
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13);
    
    \SADDRSEL_i_o2[9]\ : CFG3
      generic map(INIT => x"DF")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        B => masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        Y => N_146);
    
    masterAddrClockEnable_i_2 : CFG4
      generic map(INIT => x"FFEF")

      port map(A => N_207, B => masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        D => N_129, Y => \masterAddrClockEnable_i_2\);
    
    \SDATASELInt[0]\ : SLE
      port map(D => N_35_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_0\);
    
    \HRDATA_1_a2_3[1]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_0_0, B => N_740, C => N_737, Y => N_558);
    
    \regHADDR[2]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[2]_net_1\);
    
    \HRDATA_1_a2_3[2]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_0_1, B => N_740, C => N_737, Y => N_631);
    
    \HRDATA_1_0[14]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_3_13, C => N_737, D => N_308, 
        Y => \HRDATA_1_0[14]_net_1\);
    
    d_masterRegAddrSel_i_0 : CFG3
      generic map(INIT => x"32")

      port map(A => N_129, B => masterRegAddrSel_net_1, C => 
        N_207, Y => \d_masterRegAddrSel_i_0\);
    
    \HRDATA_1_4_1[15]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_14, B => line_1_14, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[15]_net_1\);
    
    \SADDRSEL_i_o2[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \N_135\, B => \N_120\, Y => N_151);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SDATASELInt[9]\ : SLE
      port map(D => N_49_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_9\);
    
    \PREGATEDHADDR_i_m2[13]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[13]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13, 
        Y => N_243);
    
    \HRDATA_1_4_1[17]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_16, B => line_1_16, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[17]_net_1\);
    
    \HRDATA_1_4[14]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => line_6_13, B => N_742, C => 
        \HRDATA_1_2[14]_net_1\, Y => \HRDATA_1_4[14]_net_1\);
    
    \SDATASELInt_RNO[2]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_144, B => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        C => \N_148\, Y => N_39_i_0);
    
    \HRDATA_1_0[6]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_5, C => N_737, D => N_647, 
        Y => \HRDATA_1_0[6]_net_1\);
    
    \HRDATA_1_i_a2_0_RNO[9]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => result_addr_net_0(1), B => 
        \HRDATA_1_m5_0_i_m3_1_1[9]\, C => line_3_8, D => line_4_8, 
        Y => N_523);
    
    \HRDATA_1_0[2]\ : CFG4
      generic map(INIT => x"F8F0")

      port map(A => line_4_1, B => result_addr_net_0(3), C => 
        N_627, D => N_733, Y => \HRDATA_1_0[2]_net_1\);
    
    \HRDATA_1[26]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[26]_net_1\, B => 
        \HRDATA_1_1[26]_net_1\, C => \HRDATA_1_4[26]_net_1\, D
         => \HRDATA_1_5[26]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26);
    
    \HRDATA_1[16]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[16]_net_1\, B => 
        \HRDATA_1_4[16]_net_1\, C => \HRDATA_1_1[16]_net_1\, D
         => \HRDATA_1_5[16]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16);
    
    \HRDATA_i_a2_0[28]\ : CFG3
      generic map(INIT => x"15")

      port map(A => CoreAHBLite_0_AHBmslave3_HRDATA(28), B => 
        N_320, C => N_321, Y => N_436);
    
    \HRDATA_1_4[24]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_23, D => 
        \HRDATA_1_4_1[24]_net_1\, Y => \HRDATA_1_4[24]_net_1\);
    
    \SDATASELInt_RNO[1]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \N_149\, B => \N_225\, C => \N_148\, D => 
        \N_120\, Y => N_37_i_0);
    
    hready_m_xhdl340_10_0_a2_0_a2 : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt_9\, B => \SDATASELInt_8\, C => 
        \SDATASELInt_7\, D => \SDATASELInt_6\, Y => 
        \hready_m_xhdl343_10\);
    
    \HRDATA_i_1_RNO_0[28]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_27, B => line_2_27, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \HRDATA_i_m3_1_1[28]\);
    
    \HRDATA_1_4_1[4]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_3, B => line_1_3, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[4]_net_1\);
    
    \HRDATA_i_1_RNO[28]\ : CFG4
      generic map(INIT => x"46CE")

      port map(A => result_addr_net_0(1), B => 
        \HRDATA_i_m3_1_1[28]\, C => line_27, D => line_0_27, Y
         => N_501);
    
    \HRDATA[5]\ : CFG4
      generic map(INIT => x"88C0")

      port map(A => SHA256_Module_0_data_out_5, B => 
        \un1_SDATASELInt_1\, C => 
        CoreAHBLite_0_AHBmslave3_HRDATA(5), D => \xhdl1222_2\, Y
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5);
    
    masterAddrClockEnable_i_o2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \N_138\, B => arbRegSMCurrentState_13, Y => 
        N_143);
    
    \HRDATA_1_m5_i_m3_1_1[20]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_19, B => line_6_19, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \HRDATA_1_m5_i_m3_1_1[20]_net_1\);
    
    \HRDATA_1_a2_4[2]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_1_1, B => N_739, C => N_737, Y => N_632);
    
    \regHADDR[9]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[9]_net_1\);
    
    \HRDATA_1_i_1[9]\ : CFG4
      generic map(INIT => x"FFAB")

      port map(A => N_687, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(9), C => 
        \hready_m_xhdl345\, D => N_485, Y => 
        \HRDATA_1_i_1[9]_net_1\);
    
    \regHADDR[0]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[0]_net_1\);
    
    \SDATASELInt[6]\ : SLE
      port map(D => N_43_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_6\);
    
    masterAddrClockEnable_i_o2_1 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => arbRegSMCurrentState_12, B => 
        arbRegSMCurrentState_8, C => arbRegSMCurrentState_4, D
         => arbRegSMCurrentState_0, Y => \N_138\);
    
    \HRDATA_1_a2[1]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(1), C => N_321, D => 
        \xhdl1222_2\, Y => N_555);
    
    \HRDATA[12]\ : CFG4
      generic map(INIT => x"88C0")

      port map(A => SHA256_Module_0_data_out_12, B => 
        \un1_SDATASELInt_1\, C => 
        CoreAHBLite_0_AHBmslave3_HRDATA(12), D => N_320, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12);
    
    \HRDATA_1_1[4]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_3, B => line_3_3, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[4]_net_1\);
    
    \HRDATA_1_0[10]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_9, C => N_737, D => N_657, 
        Y => \HRDATA_1_0[10]_net_1\);
    
    GATEDHTRANS_i_i2_1_m3 : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHTRANS\, B => masterRegAddrSel_net_1, C
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        Y => \N_225\);
    
    \HRDATA_1_5[14]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_4_13, B => line_5_13, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[14]_net_1\);
    
    \HRDATA_1_2[1]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => line_2_0, B => N_751, C => N_558, Y => 
        \HRDATA_1_2[1]_net_1\);
    
    \regHADDR[5]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        regHADDR_5);
    
    \HRDATA_1_4[10]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_9, D => 
        \HRDATA_1_4_1[10]_net_1\, Y => \HRDATA_1_4[10]_net_1\);
    
    \HRDATA_1_5[2]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => line_5_1, B => line_6_1, C => N_746, D => 
        N_742, Y => \HRDATA_1_5[2]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \HRDATA_1_m5_i_m3[20]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => result_addr_net_0(1), B => 
        \HRDATA_1_m5_i_m3_1_1[20]_net_1\, C => line_3_19, D => 
        line_4_19, Y => N_514);
    
    \HRDATA_1_a3[11]\ : CFG3
      generic map(INIT => x"40")

      port map(A => result_addr_net_0(3), B => N_739, C => N_733, 
        Y => N_742);
    
    \HRDATA_1_1[15]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_14, B => line_3_14, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[15]_net_1\);
    
    \SDATASELInt_RNO[4]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \N_149\, B => \N_148\, C => \SADDRSEL_i_0[4]\, 
        D => \N_225\, Y => N_41_i_0);
    
    \regHADDR[13]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[13]_net_1\);
    
    \HRDATA_1_m5_i_m3_1_1[9]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_8, B => line_2_8, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \HRDATA_1_m5_i_m3_1_1[9]_net_1\);
    
    \HRDATA_1_a3_14[11]\ : CFG2
      generic map(INIT => x"4")

      port map(A => result_addr_net_0(2), B => 
        result_addr_net_0(1), Y => N_740);
    
    \PREGATEDHADDR_i_m2[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[1]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        Y => N_246);
    
    \SDATASELInt_RNO[5]\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \N_149\, B => \N_225\, C => \N_148\, D => 
        \N_120\, Y => N_249_i_0);
    
    \regHADDR[29]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[29]_net_1\);
    
    \HRDATA_i_1_RNO_0[31]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_30, B => line_2_30, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \HRDATA_i_m3_1_1[31]\);
    
    \HRDATA_1_5[27]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_26, B => line_6_26, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[27]_net_1\);
    
    regHWRITE : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHWRITE\);
    
    \regHADDR[4]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        regHADDR_4);
    
    \SDATASELInt_RNO[14]\ : CFG3
      generic map(INIT => x"40")

      port map(A => N_144, B => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        C => \N_148\, Y => N_59_i_0);
    
    \PREGATEDHADDR_i_m3[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[2]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        Y => N_276);
    
    \HRDATA_1_5[21]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_20, B => line_6_20, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[21]_net_1\);
    
    \HRDATA_1_1[24]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_23, B => line_3_23, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[24]_net_1\);
    
    \HRDATA_1_5[29]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_28, B => line_6_28, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[29]_net_1\);
    
    \SADDRSEL_i_o2[11]\ : CFG4
      generic map(INIT => x"3F77")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        B => \N_225\, C => \regHADDR[29]_net_1\, D => 
        masterRegAddrSel_net_1, Y => \N_135\);
    
    \HRDATA_1_i_1_RNO_0[18]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_17, B => line_2_17, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \HRDATA_1_m5_0_i_m3_1_1[18]\);
    
    \HRDATA_1_a2[29]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(29), C => N_321, D => 
        \xhdl1222_2\, Y => N_425);
    
    \HRDATA_1_a2[16]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(16), C => N_321, D => 
        \xhdl1222_2\, Y => N_298);
    
    \HRDATA_1[21]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[21]_net_1\, B => 
        \HRDATA_1_5[21]_net_1\, C => \HRDATA_1_1[21]_net_1\, D
         => \HRDATA_1_4[21]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21);
    
    \HRDATA_1[11]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[11]_net_1\, B => 
        \HRDATA_1_5[11]_net_1\, C => \HRDATA_1_1[11]_net_1\, D
         => \HRDATA_1_4[11]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11);
    
    \SADDRSEL_i_0[12]\ : CFG3
      generic map(INIT => x"FD")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        B => masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        Y => \SADDRSEL_i_0[8]\);
    
    \HRDATA_1_4_1[11]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_10, B => line_1_10, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[11]_net_1\);
    
    \HRDATA_1_i_1_RNIC58O2[9]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => N_758, B => \HRDATA_1_i_1[9]_net_1\, C => 
        N_264, D => N_757, Y => N_481_i_0);
    
    \HRDATA_1_0[27]\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => \hready_m_xhdl345\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(27), C => N_564, D => 
        \un1_SDATASELInt_1\, Y => \HRDATA_1_0[27]_net_1\);
    
    \HRDATA_1[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_2[2]_net_1\, B => 
        \HRDATA_1_6[2]_net_1\, C => \HRDATA_1_5[2]_net_1\, D => 
        \HRDATA_1_1[2]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2);
    
    \HRDATA_i_a2_0[31]\ : CFG3
      generic map(INIT => x"15")

      port map(A => CoreAHBLite_0_AHBmslave3_HRDATA(31), B => 
        N_320, C => N_321, Y => N_602);
    
    \HRDATA_i_a3_0[31]\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_321, B => result_addr_net_0(0), C => N_320, 
        Y => N_755);
    
    \HRDATA_1_5[10]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_9, B => line_6_9, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[10]_net_1\);
    
    \HRDATA_1_0[21]\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => \hready_m_xhdl345\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(21), C => N_461, D => 
        \un1_SDATASELInt_1\, Y => \HRDATA_1_0[21]_net_1\);
    
    GATEDHWRITE_i_m3 : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHWRITE\, B => masterRegAddrSel_net_1, C
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        Y => N_277);
    
    \HRDATA_1_2[2]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => line_2_1, B => N_751, C => N_631, Y => 
        \HRDATA_1_2[2]_net_1\);
    
    \HRDATA_1_0[29]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_28, C => N_737, D => N_425, 
        Y => \HRDATA_1_0[29]_net_1\);
    
    \HRDATA_1_a2[6]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(6), C => N_321, D => 
        \xhdl1222_2\, Y => N_647);
    
    \SDATASELInt_RNO[0]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \N_149\, B => \N_148\, C => \SADDRSEL_i_0[4]\, 
        D => \N_225\, Y => N_35_i_0);
    
    \SDATASELInt_RNO[15]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \N_149\, B => \N_148\, C => N_146, D => 
        \N_225\, Y => N_61_i_0);
    
    \regHADDR[8]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[8]_net_1\);
    
    \SDATASELInt[11]\ : SLE
      port map(D => N_53_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_11\);
    
    \HRDATA_1_5[26]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_25, B => line_6_25, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[26]_net_1\);
    
    \HRDATA_1_a2_1[21]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_2_20, B => N_738, C => N_737, Y => N_461);
    
    \PREGATEDHADDR_i_m2[12]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[12]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12, 
        Y => N_244);
    
    \HRDATA_1_0[1]\ : CFG4
      generic map(INIT => x"F8F0")

      port map(A => line_4_0, B => result_addr_net_0(3), C => 
        N_555, D => N_733, Y => \HRDATA_1_0[1]_net_1\);
    
    \SDATASELInt[10]\ : SLE
      port map(D => N_51_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_10\);
    
    hready_m_xhdl345_0_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => N_321, B => N_320, Y => \hready_m_xhdl345\);
    
    \HRDATA_1_i_1_RNO[18]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => result_addr_net_0(1), B => 
        \HRDATA_1_m5_0_i_m3_1_1[18]\, C => line_17, D => 
        line_0_17, Y => N_517);
    
    \SDATASELInt[3]\ : SLE
      port map(D => \xhdl1221[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \xhdl1222_0\);
    
    \SDATASELInt_RNO[8]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \N_149\, B => \N_148\, C => \SADDRSEL_i_0[8]\, 
        D => \N_225\, Y => N_47_i_0);
    
    \SDATASELInt[5]\ : SLE
      port map(D => N_249_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \xhdl1222_2\);
    
    \HRDATA_1_a3_12[11]\ : CFG2
      generic map(INIT => x"8")

      port map(A => result_addr_net_0(2), B => 
        result_addr_net_0(1), Y => N_738);
    
    d_masterRegAddrSel_i_o2_0 : CFG4
      generic map(INIT => x"000B")

      port map(A => CoreAHBLite_0_AHBmslave3_HREADY_i_1, B => 
        N_143, C => N_151, D => \N_148\, Y => 
        \d_masterRegAddrSel_i_o2_0\);
    
    hready_m_xhdl343_1_0_0_a2_0 : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt_4\, B => \SDATASELInt_2\, C => 
        \SDATASELInt_1\, D => \SDATASELInt_0\, Y => N_318);
    
    \HRDATA_1_a2_4[7]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_6_d0, B => N_739, C => N_737, Y => N_587);
    
    \SADDRSEL_i_0[0]\ : CFG4
      generic map(INIT => x"DDD8")

      port map(A => masterRegAddrSel_net_1, B => \regHTRANS\, C
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        Y => \SADDRSEL_i_0[4]\);
    
    \HRDATA_1[3]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[3]_net_1\, B => 
        \HRDATA_1_1[3]_net_1\, C => \HRDATA_1_4[3]_net_1\, D => 
        \HRDATA_1_5[3]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3);
    
    \HRDATA_1_4_1[26]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_25, B => line_1_25, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[26]_net_1\);
    
    \HRDATA_1_i_1[18]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => N_755, B => N_485, C => N_681, D => N_517, Y
         => \HRDATA_1_i_1[18]_net_1\);
    
    \HRDATA_1_5[22]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_21, B => line_6_21, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[22]_net_1\);
    
    hready_m_xhdl343_1_0_0_a2_0_RNIHM4M1 : CFG4
      generic map(INIT => x"A8A0")

      port map(A => N_335, B => N_214, C => 
        un1_hready_m_xhdl343_1_i_0_a2_1, D => N_305, Y => 
        un1_hready_m_xhdl343_1_i_0_o2_0);
    
    \HRDATA_1_4[30]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_29, D => 
        \HRDATA_1_4_1[30]_net_1\, Y => \HRDATA_1_4[30]_net_1\);
    
    \SDATASELInt_RNO[7]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \N_135\, B => \N_120\, C => \N_148\, Y => 
        N_45_i_1);
    
    \HRDATA_1_4[3]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_2_d0, D => 
        \HRDATA_1_4_1[3]_net_1\, Y => \HRDATA_1_4[3]_net_1\);
    
    \SADDRSEL_i_o2_1_o2[4]\ : CFG3
      generic map(INIT => x"DF")

      port map(A => \N_225\, B => \N_149\, C => \N_148\, Y => 
        N_127);
    
    \HRDATA_1_4_1[3]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_2, B => line_1_2, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[3]_net_1\);
    
    \HRDATA_1_0[26]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_25, C => N_737, D => N_439, 
        Y => \HRDATA_1_0[26]_net_1\);
    
    \HRDATA_1_0[17]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_16, C => N_737, D => N_607, 
        Y => \HRDATA_1_0[17]_net_1\);
    
    \PREGATEDHADDR_i_m3[8]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[8]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        Y => N_257);
    
    \HRDATA_1_6[2]\ : CFG4
      generic map(INIT => x"FFEA")

      port map(A => N_632, B => N_748, C => line_7(2), D => 
        \HRDATA_1_0[2]_net_1\, Y => \HRDATA_1_6[2]_net_1\);
    
    \HRDATA_1_m5_i_m3_1_1[18]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_17, B => line_6_17, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \HRDATA_1_m5_i_m3_1_1[18]_net_1\);
    
    \HRDATA_1_0[11]\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => \hready_m_xhdl345\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(11), C => N_536, D => 
        \un1_SDATASELInt_1\, Y => \HRDATA_1_0[11]_net_1\);
    
    \HRDATA_1_a2[25]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(25), C => N_321, D => 
        \xhdl1222_2\, Y => N_637);
    
    \HRDATA_1_4[6]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_5_d0, D => 
        \HRDATA_1_4_1[6]_net_1\, Y => \HRDATA_1_4[6]_net_1\);
    
    \HRDATA_1_1[30]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_29, B => line_3_29, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[30]_net_1\);
    
    \HRDATA_1_0[19]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_18, C => N_737, D => N_469, 
        Y => \HRDATA_1_0[19]_net_1\);
    
    hready_m_xhdl345_0_a2_RNICTNV7 : CFG2
      generic map(INIT => x"1")

      port map(A => N_129, B => N_207, Y => N_9_i_0);
    
    \HRDATA_1_4[17]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_16, D => 
        \HRDATA_1_4_1[17]_net_1\, Y => \HRDATA_1_4[17]_net_1\);
    
    \HRDATA_1_i_1_RNIPTLS2[20]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => N_758, B => \HRDATA_1_i_1[20]_net_1\, C => 
        N_514, D => N_757, Y => N_479_i_0);
    
    \HRDATA_1_4_1[25]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_24, B => line_1_24, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[25]_net_1\);
    
    \HRDATA_1_4[11]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_10, D => 
        \HRDATA_1_4_1[11]_net_1\, Y => \HRDATA_1_4[11]_net_1\);
    
    \HRDATA_1_a2[7]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(7), C => N_321, D => 
        \xhdl1222_2\, Y => N_582);
    
    \PREGATEDHADDR_i_m2[30]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[30]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        Y => \N_148\);
    
    \HRDATA_1_4[19]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_18, D => 
        \HRDATA_1_4_1[19]_net_1\, Y => \HRDATA_1_4[19]_net_1\);
    
    \HRDATA_1_4_1[27]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_26, B => line_1_26, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[27]_net_1\);
    
    \HRDATA_1_0[22]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_21, C => N_737, D => N_572, 
        Y => \HRDATA_1_0[22]_net_1\);
    
    \HRDATA_1_i_a2_0_RNO[20]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => result_addr_net_0(1), B => 
        \HRDATA_1_m5_0_i_m3_1_1[20]\, C => line_19, D => 
        line_0_19, Y => N_511);
    
    \HRDATA_1_4[27]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_26, D => 
        \HRDATA_1_4_1[27]_net_1\, Y => \HRDATA_1_4[27]_net_1\);
    
    \SDATASELInt_RNIDUN21[14]\ : CFG4
      generic map(INIT => x"7610")

      port map(A => \SDATASELInt[15]_net_1\, B => 
        \SDATASELInt[14]_net_1\, C => N_215, D => 
        \hready_m_xhdl343_10\, Y => 
        un1_hready_m_xhdl343_1_i_0_o2_1_tz);
    
    \HRDATA_1_a2_1[11]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_2_10, B => N_738, C => N_737, Y => N_536);
    
    \HRDATA_1_4[7]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => line_6_6, B => N_742, C => 
        \HRDATA_1_2[7]_net_1\, Y => \HRDATA_1_4[7]_net_1\);
    
    \HRDATA_1_a2[14]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(14), C => N_321, D => 
        \xhdl1222_2\, Y => N_308);
    
    \HRDATA_1_4[21]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_20, D => 
        \HRDATA_1_4_1[21]_net_1\, Y => \HRDATA_1_4[21]_net_1\);
    
    \HRDATA_1_4[29]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_28, D => 
        \HRDATA_1_4_1[29]_net_1\, Y => \HRDATA_1_4[29]_net_1\);
    
    hready_m_xhdl345_0_a2_RNI0HL74 : CFG4
      generic map(INIT => x"0D00")

      port map(A => masterDataInProg_0(0), B => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, C => 
        \hready_m_xhdl345\, D => \un1_SDATASELInt_1\, Y => N_207);
    
    \HRDATA_1_1[14]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_1_13, B => line_2_13, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[14]_net_1\);
    
    \PREGATEDHADDR_i_m2[0]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[0]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        Y => N_247);
    
    \HRDATA_1[6]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[6]_net_1\, B => 
        \HRDATA_1_1[6]_net_1\, C => \HRDATA_1_4[6]_net_1\, D => 
        \HRDATA_1_5[6]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6);
    
    \HRDATA_1_1[7]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_1_6, B => line_2_6, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[7]_net_1\);
    
    \HRDATA_1_m5_i_m3[9]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => result_addr_net_0(1), B => 
        \HRDATA_1_m5_i_m3_1_1[9]_net_1\, C => line_8, D => 
        line_0_8, Y => N_264);
    
    \SADDRSEL_i_o2[2]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        B => \N_135\, C => masterRegAddrSel_net_1, Y => N_144);
    
    masterAddrClockEnable_i_5_RNIU9KI1 : CFG4
      generic map(INIT => x"0F0D")

      port map(A => CertificationSystem_sb_0_AHBmslave5_HREADY, B
         => N_249, C => \masterAddrClockEnable_i_5\, D => N_226, 
        Y => N_106_i_0);
    
    \HRDATA_1_i_1_RNISSHS2[18]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => N_758, B => \HRDATA_1_i_1[18]_net_1\, C => 
        N_520, D => N_757, Y => N_480_i_0);
    
    \SDATASELInt[15]\ : SLE
      port map(D => N_61_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[15]_net_1\);
    
    \HRDATA_1_0[16]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_741, B => line_4_15, C => N_737, D => N_298, 
        Y => \HRDATA_1_0[16]_net_1\);
    
    \HRDATA_1_a2[17]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(17), C => N_321, D => 
        \xhdl1222_2\, Y => N_607);
    
    \HRDATA_i_o2[31]\ : CFG4
      generic map(INIT => x"B7BF")

      port map(A => \xhdl1222_2\, B => N_321, C => \xhdl1222_0\, 
        D => ren_pos, Y => N_485);
    
    \HRDATA_1_5[30]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_29, B => line_6_29, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[30]_net_1\);
    
    \HRDATA_1_5[25]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_24, B => line_6_24, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[25]_net_1\);
    
    \HRDATA_1_4[16]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_15, D => 
        \HRDATA_1_4_1[16]_net_1\, Y => \HRDATA_1_4[16]_net_1\);
    
    un1_SDATASELInt_1_0_a2 : CFG3
      generic map(INIT => x"60")

      port map(A => \xhdl1222_0\, B => \xhdl1222_2\, C => N_321, 
        Y => \un1_SDATASELInt_1\);
    
    \HRDATA_1_1[1]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => line_3_0, B => N_750, C => N_556, Y => 
        \HRDATA_1_1[1]_net_1\);
    
    \HRDATA_1_5[1]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => line_5_0, B => line_6_0, C => N_748, D => 
        N_742, Y => \HRDATA_1_5[1]_net_1\);
    
    \HRDATA_1_a2_1[1]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_0_d0, B => N_738, C => N_737, Y => N_556);
    
    \HRDATA_1_0[30]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_29, C => N_737, D => N_415, 
        Y => \HRDATA_1_0[30]_net_1\);
    
    \HRDATA_1_5[17]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_16, B => line_6_16, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[17]_net_1\);
    
    \PREGATEDHADDR_i_m3[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[7]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7, 
        Y => N_258);
    
    \PREGATEDHADDR_i_m2_RNI1D521[29]\ : CFG4
      generic map(INIT => x"FFBF")

      port map(A => \N_149\, B => \N_225\, C => \N_148\, D => 
        \N_120\, Y => N_249);
    
    \HRDATA_1_4_1[19]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_18, B => line_1_18, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[19]_net_1\);
    
    \HRDATA_1_4[26]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_25, D => 
        \HRDATA_1_4_1[26]_net_1\, Y => \HRDATA_1_4[26]_net_1\);
    
    \HRDATA_1[10]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[10]_net_1\, B => 
        \HRDATA_1_1[10]_net_1\, C => \HRDATA_1_4[10]_net_1\, D
         => \HRDATA_1_5[10]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10);
    
    \regHADDR[6]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[6]_net_1\);
    
    \HRDATA_1_5[11]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_10, B => line_6_10, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[11]_net_1\);
    
    \HRDATA_1_5[19]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_18, B => line_6_18, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[19]_net_1\);
    
    \HRDATA_i_a3_2[31]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => result_addr_net_0(0), B => 
        result_addr_net_0(3), C => N_321, D => N_320, Y => N_758);
    
    \masterRegAddrSel\ : SLE
      port map(D => N_108_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        masterRegAddrSel_net_1);
    
    hready_m_xhdl343_1_0_0_a2_0_RNIATE83 : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_318, B => N_305, C => 
        un1_hready_m_xhdl343_1_i_0_o2_1_tz, D => 
        un1_hready_m_xhdl343_1_i_0_o2_0, Y => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\);
    
    \HRDATA_1_a3_5[11]\ : CFG3
      generic map(INIT => x"40")

      port map(A => result_addr_net_0(3), B => N_741, C => N_733, 
        Y => N_748);
    
    \HRDATA_1_a2_4[1]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_1_0, B => N_739, C => N_737, Y => N_559);
    
    \HRDATA_1[4]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[4]_net_1\, B => 
        \HRDATA_1_1[4]_net_1\, C => \HRDATA_1_4[4]_net_1\, D => 
        \HRDATA_1_5[4]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4);
    
    \HRDATA_1_m5_i_m3[18]\ : CFG4
      generic map(INIT => x"B931")

      port map(A => result_addr_net_0(1), B => 
        \HRDATA_1_m5_i_m3_1_1[18]_net_1\, C => line_3_17, D => 
        line_4_17, Y => N_520);
    
    \HRDATA_1_i_a2[18]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \xhdl1222_2\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(18), C => \xhdl1222_0\, Y
         => N_681);
    
    \HRDATA_1_1[6]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_5, B => line_3_5, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[6]_net_1\);
    
    \HRDATA[0]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => \hready_m_xhdl345\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(0), C => 
        SHA256_Module_0_data_out_0, D => \un1_SDATASELInt_1\, Y
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0);
    
    \HRDATA_1_a2_1[16]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_2_15, B => N_738, C => N_737, Y => N_543);
    
    \HRDATA_i_1_RNIJ96R2[31]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => N_758, B => \HRDATA_i_1[31]_net_1\, C => 
        N_507, D => N_757, Y => N_477_i_0);
    
    \SDATASELInt_RNIJDUB4[3]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un8_hreadyin_i_0, B => \N_206\, Y => N_27_i_0);
    
    \HRDATA_1_4[22]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_21, D => 
        \HRDATA_1_4_1[22]_net_1\, Y => \HRDATA_1_4[22]_net_1\);
    
    \HRDATA_1_0[25]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_24, C => N_737, D => N_637, 
        Y => \HRDATA_1_0[25]_net_1\);
    
    \regHADDR[14]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[14]_net_1\);
    
    \HRDATA_1_a2_1[27]\ : CFG3
      generic map(INIT => x"80")

      port map(A => line_2_26, B => N_738, C => N_737, Y => N_564);
    
    \SDATASELInt_RNO[13]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \N_149\, B => \N_148\, C => N_146, D => 
        \N_225\, Y => N_57_i_1);
    
    \HRDATA_1_1[10]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_9, B => line_3_9, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[10]_net_1\);
    
    DEFSLAVEDATASEL_i_a2 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_318, B => \hready_m_xhdl343_10\, C => 
        \hready_m_xhdl344_7\, D => \hready_m_xhdl343_11\, Y => 
        N_321);
    
    \HRDATA_1_1[27]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_3_26, B => line_4_26, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[27]_net_1\);
    
    \SADDRSEL_i_o2_RNIB5R01[11]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \N_135\, B => \N_120\, C => \N_148\, Y => 
        \xhdl1221[3]\);
    
    \regHADDR[10]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[10]_net_1\);
    
    \HRDATA_1_1[21]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_3_20, B => line_4_20, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[21]_net_1\);
    
    \HRDATA_1_5[4]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_3, B => line_6_3, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[4]_net_1\);
    
    \HRDATA_1_4_1[10]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_9, B => line_1_9, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[10]_net_1\);
    
    \HRDATA_1_1[29]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_28, B => line_3_28, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[29]_net_1\);
    
    \SDATASELInt[1]\ : SLE
      port map(D => N_37_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_1\);
    
    \PREGATEDHADDR_i_m2[15]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[15]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15, 
        Y => N_241);
    
    \HRDATA_1_4[4]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_3_d0, D => 
        \HRDATA_1_4_1[4]_net_1\, Y => \HRDATA_1_4[4]_net_1\);
    
    \HRDATA_1[24]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[24]_net_1\, B => 
        \HRDATA_1_1[24]_net_1\, C => \HRDATA_1_4[24]_net_1\, D
         => \HRDATA_1_5[24]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24);
    
    \HRDATA_1[14]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_1[14]_net_1\, B => 
        \HRDATA_1_0[14]_net_1\, C => \HRDATA_1_4[14]_net_1\, D
         => \HRDATA_1_5[14]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14);
    
    \HRDATA_1_a3_15[11]\ : CFG2
      generic map(INIT => x"2")

      port map(A => result_addr_net_0(2), B => 
        result_addr_net_0(1), Y => N_741);
    
    \HRDATA_1_i_a2_0_RNO_0[20]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_1_19, B => line_2_19, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \HRDATA_1_m5_0_i_m3_1_1[20]\);
    
    \HRDATA_1_a3_9[11]\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_321, B => result_addr_net_0(0), C => 
        \HRDATA_1_a3_17_0[11]_net_1\, Y => N_733);
    
    \HRDATA_1_a3_17_0[11]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \xhdl1222_2\, B => \xhdl1222_0\, C => ren_pos, 
        Y => \HRDATA_1_a3_17_0[11]_net_1\);
    
    \HRDATA_1_5[16]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_15, B => line_6_15, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[16]_net_1\);
    
    \regHADDR[11]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        regHADDR_11);
    
    \HRDATA_1_4_1[6]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_5, B => line_1_5, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[6]_net_1\);
    
    \PREGATEDHADDR_i_m3[9]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[9]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9, 
        Y => N_256);
    
    \HRDATA_1[22]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[22]_net_1\, B => 
        \HRDATA_1_1[22]_net_1\, C => \HRDATA_1_4[22]_net_1\, D
         => \HRDATA_1_5[22]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22);
    
    \HRDATA_1_5[7]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_4_6, B => line_5_6, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[7]_net_1\);
    
    \HRDATA_1_2[7]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => line_0_6, B => N_740, C => N_737, D => N_587, 
        Y => \HRDATA_1_2[7]_net_1\);
    
    \regHADDR[7]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[7]_net_1\);
    
    \GATEDHSIZE_i_m2[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHSIZE[1]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1), 
        Y => N_235);
    
    \SDATASELInt[14]\ : SLE
      port map(D => N_59_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt[14]_net_1\);
    
    \HRDATA_1_i_a2_0_RNO_0[9]\ : CFG4
      generic map(INIT => x"0F35")

      port map(A => line_5_8, B => line_6_8, C => 
        result_addr_net_0(2), D => result_addr_net_0(1), Y => 
        \HRDATA_1_m5_0_i_m3_1_1[9]\);
    
    \PREGATEDHADDR_i_m2[29]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[29]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        Y => \N_149\);
    
    \regHADDR[3]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        regHADDR_3);
    
    \HRDATA_1_5[3]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_2, B => line_6_2, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[3]_net_1\);
    
    \HRDATA_1_4_1[21]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_20, B => line_1_20, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[21]_net_1\);
    
    \HRDATA_1_a2[26]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(26), C => N_321, D => 
        \xhdl1222_2\, Y => N_439);
    
    regHTRANS : SLE
      port map(D => VCC_net_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_106_i_0, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \regHTRANS\);
    
    \PREGATEDHADDR_i_m3[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[6]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        Y => N_259);
    
    masterAddrClockEnable_i_a2 : CFG4
      generic map(INIT => x"000E")

      port map(A => arbRegSMCurrentState_13, B => \N_138\, C => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, D => \N_148\, Y => 
        N_178);
    
    \HRDATA_1_0[4]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_3, C => N_737, D => N_592, 
        Y => \HRDATA_1_0[4]_net_1\);
    
    \SDATASELInt_RNO[6]\ : CFG3
      generic map(INIT => x"10")

      port map(A => N_144, B => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        C => \N_148\, Y => N_43_i_0);
    
    \HRDATA_1_4_1[30]\ : CFG4
      generic map(INIT => x"153F")

      port map(A => line_0_29, B => line_1_29, C => N_740, D => 
        N_739, Y => \HRDATA_1_4_1[30]_net_1\);
    
    \SDATASELInt_RNO[10]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_144, B => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        C => \N_148\, Y => N_51_i_0);
    
    \HRDATA[8]\ : CFG4
      generic map(INIT => x"88C0")

      port map(A => SHA256_Module_0_data_out_8, B => 
        \un1_SDATASELInt_1\, C => 
        CoreAHBLite_0_AHBmslave3_HRDATA(8), D => N_320, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8);
    
    masterAddrClockEnable_i_x2 : CFG4
      generic map(INIT => x"3C66")

      port map(A => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        B => \N_149\, C => \regHADDR[30]_net_1\, D => 
        masterRegAddrSel_net_1, Y => N_142_i);
    
    \SDATASELInt[12]\ : SLE
      port map(D => N_55_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_12\);
    
    \regHADDR[1]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[1]_net_1\);
    
    \HRDATA_1_0[15]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_738, B => line_4_14, C => N_737, D => N_617, 
        Y => \HRDATA_1_0[15]_net_1\);
    
    masterAddrClockEnable_i_5 : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \masterAddrClockEnable_i_2\, B => \N_120\, C
         => N_142_i, D => N_178, Y => \masterAddrClockEnable_i_5\);
    
    \HRDATA_1_1[26]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_25, B => line_3_25, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[26]_net_1\);
    
    \HRDATA_1_a3_7[11]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \HRDATA_1_a3_17_0[11]_net_1\, B => N_321, C
         => result_addr_net_0(0), D => 
        \HRDATA_1_a3_7_0[11]_net_1\, Y => N_750);
    
    \HRDATA_1_1[2]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => line_3_1, B => N_750, C => N_629, Y => 
        \HRDATA_1_1[2]_net_1\);
    
    \PREGATEDHADDR_i_m3[10]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[10]_net_1\, B => 
        masterRegAddrSel_net_1, C => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10, 
        Y => N_255);
    
    \HRDATA_1_4[15]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_14, D => 
        \HRDATA_1_4_1[15]_net_1\, Y => \HRDATA_1_4[15]_net_1\);
    
    HREADY_M_iv_i_i_o2_1 : CFG2
      generic map(INIT => x"7")

      port map(A => masterDataInProg(0), B => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, Y => N_126);
    
    \HRDATA_1[29]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[29]_net_1\, B => 
        \HRDATA_1_1[29]_net_1\, C => \HRDATA_1_4[29]_net_1\, D
         => \HRDATA_1_5[29]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29);
    
    \HRDATA_1[19]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[19]_net_1\, B => 
        \HRDATA_1_1[19]_net_1\, C => \HRDATA_1_4[19]_net_1\, D
         => \HRDATA_1_5[19]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19);
    
    \HRDATA_1_a2[22]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(22), C => N_321, D => 
        \xhdl1222_2\, Y => N_572);
    
    \HRDATA_1_6[1]\ : CFG4
      generic map(INIT => x"FFEA")

      port map(A => N_559, B => N_746, C => line_7(1), D => 
        \HRDATA_1_0[1]_net_1\, Y => \HRDATA_1_6[1]_net_1\);
    
    \HRDATA_1_a3_11[11]\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_321, B => result_addr_net_0(0), C => 
        \HRDATA_1_a3_17_0[11]_net_1\, Y => N_737);
    
    \SDATASELInt_RNO[11]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \N_149\, B => \N_148\, C => N_146, D => 
        \N_225\, Y => N_53_i_0);
    
    \HRDATA_1_4[25]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_737, B => N_742, C => line_24, D => 
        \HRDATA_1_4_1[25]_net_1\, Y => \HRDATA_1_4[25]_net_1\);
    
    \HRDATA_1[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_2[1]_net_1\, B => 
        \HRDATA_1_6[1]_net_1\, C => \HRDATA_1_5[1]_net_1\, D => 
        \HRDATA_1_1[1]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1);
    
    \HRDATA_i_a3_1[31]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => result_addr_net_0(0), B => 
        result_addr_net_0(3), C => N_321, D => N_320, Y => N_757);
    
    \HRDATA_1_i_1[20]\ : CFG4
      generic map(INIT => x"FFAB")

      port map(A => N_678, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(20), C => 
        \hready_m_xhdl345\, D => N_485, Y => 
        \HRDATA_1_i_1[20]_net_1\);
    
    \HRDATA_1_1[22]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_21, B => line_3_21, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[22]_net_1\);
    
    \HRDATA_1[7]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_1[7]_net_1\, B => 
        \HRDATA_1_0[7]_net_1\, C => \HRDATA_1_4[7]_net_1\, D => 
        \HRDATA_1_5[7]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7);
    
    \HRDATA_1_i_a2_0[20]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => N_511, B => N_321, C => result_addr_net_0(0), 
        D => N_320, Y => N_678);
    
    \regHADDR[12]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12, 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHADDR[12]_net_1\);
    
    \HRDATA_1_a2[2]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(2), C => N_321, D => 
        \xhdl1222_2\, Y => N_627);
    
    \SDATASELInt[8]\ : SLE
      port map(D => N_47_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_8\);
    
    \SDATASELInt[2]\ : SLE
      port map(D => N_39_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_2\);
    
    \HRDATA_1_a2[30]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(30), C => N_321, D => 
        \xhdl1222_2\, Y => N_415);
    
    \HRDATA_1_1[3]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_2_2, B => line_3_2, C => N_751, D => 
        N_750, Y => \HRDATA_1_1[3]_net_1\);
    
    \regHSIZE[1]\ : SLE
      port map(D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1), 
        CLK => CertificationSystem_sb_0_FAB_CCC_GL0, EN => 
        N_106_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \regHSIZE[1]_net_1\);
    
    \HRDATA_1[27]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[27]_net_1\, B => 
        \HRDATA_1_5[27]_net_1\, C => \HRDATA_1_1[27]_net_1\, D
         => \HRDATA_1_4[27]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27);
    
    \HRDATA_1[17]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \HRDATA_1_0[17]_net_1\, B => 
        \HRDATA_1_1[17]_net_1\, C => \HRDATA_1_4[17]_net_1\, D
         => \HRDATA_1_5[17]_net_1\, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17);
    
    \HRDATA_1_a2[4]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(4), C => N_321, D => 
        \xhdl1222_2\, Y => N_592);
    
    \SDATASELInt_RNIE2CB4[3]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \xhdl1222_2\, B => \xhdl1222_0\, C => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, D => N_321, Y => 
        \N_206\);
    
    \SDATASELInt[4]\ : SLE
      port map(D => N_41_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_27_i_0, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \SDATASELInt_4\);
    
    \HRDATA_i_1_RNIHH261[28]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => N_758, B => \HRDATA_i_1[28]_net_1\, C => 
        N_436, D => N_485, Y => N_478_i_0);
    
    \HRDATA[23]\ : CFG4
      generic map(INIT => x"88C0")

      port map(A => SHA256_Module_0_data_out_23, B => 
        \un1_SDATASELInt_1\, C => 
        CoreAHBLite_0_AHBmslave3_HRDATA(23), D => N_320, Y => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23);
    
    \SDATASELInt_RNO[12]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \N_149\, B => \N_148\, C => \SADDRSEL_i_0[8]\, 
        D => \N_225\, Y => N_55_i_0);
    
    \HRDATA_1_a2[19]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(19), C => N_321, D => 
        \xhdl1222_2\, Y => N_469);
    
    \HRDATA_1_a2[3]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \xhdl1222_0\, B => 
        CoreAHBLite_0_AHBmslave3_HRDATA(3), C => N_321, D => 
        \xhdl1222_2\, Y => N_667);
    
    \HRDATA_1_5[24]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => line_5_23, B => line_6_23, C => N_748, D => 
        N_746, Y => \HRDATA_1_5[24]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MATRIX4X16 is

    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE     : in    std_logic_vector(1 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS    : in    std_logic_vector(1 to 1);
          result_addr_net_0                                           : in    std_logic_vector(3 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP     : out   std_logic_vector(0 to 0);
          CoreAHBLite_0_AHBmslave3_HRDATA                             : in    std_logic_vector(31 downto 0);
          line_7                                                      : in    std_logic_vector(2 downto 1);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA    : in    std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave3_HADDR                              : out   std_logic_vector(11 to 11);
          xhdl1222_0                                                  : out   std_logic;
          xhdl1222_2                                                  : out   std_logic;
          SDATASELInt_0                                               : out   std_logic;
          SDATASELInt_1                                               : out   std_logic;
          SDATASELInt_2                                               : out   std_logic;
          SDATASELInt_4                                               : out   std_logic;
          SDATASELInt_6                                               : out   std_logic;
          SDATASELInt_7                                               : out   std_logic;
          SDATASELInt_8                                               : out   std_logic;
          SDATASELInt_9                                               : out   std_logic;
          SDATASELInt_10                                              : out   std_logic;
          SDATASELInt_11                                              : out   std_logic;
          SDATASELInt_12                                              : out   std_logic;
          SDATASELInt_13                                              : out   std_logic;
          arbRegSMCurrentState_13                                     : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31  : in    std_logic;
          line_13                                                     : in    std_logic;
          line_10                                                     : in    std_logic;
          line_21                                                     : in    std_logic;
          line_24                                                     : in    std_logic;
          line_18                                                     : in    std_logic;
          line_23                                                     : in    std_logic;
          line_16                                                     : in    std_logic;
          line_28                                                     : in    std_logic;
          line_9                                                      : in    std_logic;
          line_3_d0                                                   : in    std_logic;
          line_5_d0                                                   : in    std_logic;
          line_15                                                     : in    std_logic;
          line_26                                                     : in    std_logic;
          line_14                                                     : in    std_logic;
          line_20                                                     : in    std_logic;
          line_2_d0                                                   : in    std_logic;
          line_25                                                     : in    std_logic;
          line_29                                                     : in    std_logic;
          line_19                                                     : in    std_logic;
          line_27                                                     : in    std_logic;
          line_30                                                     : in    std_logic;
          line_17                                                     : in    std_logic;
          line_8                                                      : in    std_logic;
          line_0_d0                                                   : in    std_logic;
          line_6_d0                                                   : in    std_logic;
          line_1_d0                                                   : in    std_logic;
          line_0_10                                                   : in    std_logic;
          line_0_21                                                   : in    std_logic;
          line_0_24                                                   : in    std_logic;
          line_0_18                                                   : in    std_logic;
          line_0_23                                                   : in    std_logic;
          line_0_16                                                   : in    std_logic;
          line_0_28                                                   : in    std_logic;
          line_0_9                                                    : in    std_logic;
          line_0_3                                                    : in    std_logic;
          line_0_5                                                    : in    std_logic;
          line_0_15                                                   : in    std_logic;
          line_0_26                                                   : in    std_logic;
          line_0_14                                                   : in    std_logic;
          line_0_20                                                   : in    std_logic;
          line_0_2                                                    : in    std_logic;
          line_0_25                                                   : in    std_logic;
          line_0_29                                                   : in    std_logic;
          line_0_19                                                   : in    std_logic;
          line_0_27                                                   : in    std_logic;
          line_0_30                                                   : in    std_logic;
          line_0_17                                                   : in    std_logic;
          line_0_8                                                    : in    std_logic;
          line_0_0                                                    : in    std_logic;
          line_0_1                                                    : in    std_logic;
          line_0_6                                                    : in    std_logic;
          line_0_13                                                   : in    std_logic;
          line_1_10                                                   : in    std_logic;
          line_1_21                                                   : in    std_logic;
          line_1_24                                                   : in    std_logic;
          line_1_18                                                   : in    std_logic;
          line_1_23                                                   : in    std_logic;
          line_1_16                                                   : in    std_logic;
          line_1_28                                                   : in    std_logic;
          line_1_9                                                    : in    std_logic;
          line_1_3                                                    : in    std_logic;
          line_1_5                                                    : in    std_logic;
          line_1_15                                                   : in    std_logic;
          line_1_26                                                   : in    std_logic;
          line_1_14                                                   : in    std_logic;
          line_1_20                                                   : in    std_logic;
          line_1_2                                                    : in    std_logic;
          line_1_25                                                   : in    std_logic;
          line_1_29                                                   : in    std_logic;
          line_1_19                                                   : in    std_logic;
          line_1_27                                                   : in    std_logic;
          line_1_30                                                   : in    std_logic;
          line_1_17                                                   : in    std_logic;
          line_1_8                                                    : in    std_logic;
          line_1_0                                                    : in    std_logic;
          line_1_1                                                    : in    std_logic;
          line_1_6                                                    : in    std_logic;
          line_1_13                                                   : in    std_logic;
          line_2_19                                                   : in    std_logic;
          line_2_27                                                   : in    std_logic;
          line_2_30                                                   : in    std_logic;
          line_2_17                                                   : in    std_logic;
          line_2_8                                                    : in    std_logic;
          line_2_10                                                   : in    std_logic;
          line_2_15                                                   : in    std_logic;
          line_2_26                                                   : in    std_logic;
          line_2_20                                                   : in    std_logic;
          line_2_0                                                    : in    std_logic;
          line_2_1                                                    : in    std_logic;
          line_2_29                                                   : in    std_logic;
          line_2_25                                                   : in    std_logic;
          line_2_2                                                    : in    std_logic;
          line_2_6                                                    : in    std_logic;
          line_2_13                                                   : in    std_logic;
          line_2_14                                                   : in    std_logic;
          line_2_5                                                    : in    std_logic;
          line_2_3                                                    : in    std_logic;
          line_2_9                                                    : in    std_logic;
          line_2_28                                                   : in    std_logic;
          line_2_16                                                   : in    std_logic;
          line_2_23                                                   : in    std_logic;
          line_2_18                                                   : in    std_logic;
          line_2_24                                                   : in    std_logic;
          line_2_21                                                   : in    std_logic;
          line_3_19                                                   : in    std_logic;
          line_3_17                                                   : in    std_logic;
          line_3_8                                                    : in    std_logic;
          line_3_0                                                    : in    std_logic;
          line_3_1                                                    : in    std_logic;
          line_3_29                                                   : in    std_logic;
          line_3_25                                                   : in    std_logic;
          line_3_2                                                    : in    std_logic;
          line_3_20                                                   : in    std_logic;
          line_3_6                                                    : in    std_logic;
          line_3_13                                                   : in    std_logic;
          line_3_14                                                   : in    std_logic;
          line_3_26                                                   : in    std_logic;
          line_3_15                                                   : in    std_logic;
          line_3_5                                                    : in    std_logic;
          line_3_3                                                    : in    std_logic;
          line_3_9                                                    : in    std_logic;
          line_3_28                                                   : in    std_logic;
          line_3_16                                                   : in    std_logic;
          line_3_23                                                   : in    std_logic;
          line_3_18                                                   : in    std_logic;
          line_3_24                                                   : in    std_logic;
          line_3_21                                                   : in    std_logic;
          line_3_10                                                   : in    std_logic;
          SHA256_Module_0_data_out_5                                  : in    std_logic;
          SHA256_Module_0_data_out_13                                 : in    std_logic;
          SHA256_Module_0_data_out_12                                 : in    std_logic;
          SHA256_Module_0_data_out_8                                  : in    std_logic;
          SHA256_Module_0_data_out_23                                 : in    std_logic;
          SHA256_Module_0_data_out_0                                  : in    std_logic;
          line_4_19                                                   : in    std_logic;
          line_4_17                                                   : in    std_logic;
          line_4_8                                                    : in    std_logic;
          line_4_0                                                    : in    std_logic;
          line_4_1                                                    : in    std_logic;
          line_4_29                                                   : in    std_logic;
          line_4_25                                                   : in    std_logic;
          line_4_2                                                    : in    std_logic;
          line_4_20                                                   : in    std_logic;
          line_4_14                                                   : in    std_logic;
          line_4_26                                                   : in    std_logic;
          line_4_15                                                   : in    std_logic;
          line_4_5                                                    : in    std_logic;
          line_4_3                                                    : in    std_logic;
          line_4_9                                                    : in    std_logic;
          line_4_28                                                   : in    std_logic;
          line_4_16                                                   : in    std_logic;
          line_4_23                                                   : in    std_logic;
          line_4_18                                                   : in    std_logic;
          line_4_24                                                   : in    std_logic;
          line_4_21                                                   : in    std_logic;
          line_4_10                                                   : in    std_logic;
          line_4_6                                                    : in    std_logic;
          line_4_13                                                   : in    std_logic;
          line_5_19                                                   : in    std_logic;
          line_5_17                                                   : in    std_logic;
          line_5_8                                                    : in    std_logic;
          line_5_0                                                    : in    std_logic;
          line_5_1                                                    : in    std_logic;
          line_5_29                                                   : in    std_logic;
          line_5_25                                                   : in    std_logic;
          line_5_2                                                    : in    std_logic;
          line_5_20                                                   : in    std_logic;
          line_5_6                                                    : in    std_logic;
          line_5_13                                                   : in    std_logic;
          line_5_14                                                   : in    std_logic;
          line_5_26                                                   : in    std_logic;
          line_5_15                                                   : in    std_logic;
          line_5_5                                                    : in    std_logic;
          line_5_3                                                    : in    std_logic;
          line_5_9                                                    : in    std_logic;
          line_5_28                                                   : in    std_logic;
          line_5_16                                                   : in    std_logic;
          line_5_23                                                   : in    std_logic;
          line_5_18                                                   : in    std_logic;
          line_5_24                                                   : in    std_logic;
          line_5_21                                                   : in    std_logic;
          line_5_10                                                   : in    std_logic;
          line_6_19                                                   : in    std_logic;
          line_6_17                                                   : in    std_logic;
          line_6_8                                                    : in    std_logic;
          line_6_0                                                    : in    std_logic;
          line_6_1                                                    : in    std_logic;
          line_6_29                                                   : in    std_logic;
          line_6_25                                                   : in    std_logic;
          line_6_2                                                    : in    std_logic;
          line_6_20                                                   : in    std_logic;
          line_6_6                                                    : in    std_logic;
          line_6_13                                                   : in    std_logic;
          line_6_14                                                   : in    std_logic;
          line_6_26                                                   : in    std_logic;
          line_6_15                                                   : in    std_logic;
          line_6_5                                                    : in    std_logic;
          line_6_3                                                    : in    std_logic;
          line_6_9                                                    : in    std_logic;
          line_6_28                                                   : in    std_logic;
          line_6_16                                                   : in    std_logic;
          line_6_23                                                   : in    std_logic;
          line_6_18                                                   : in    std_logic;
          line_6_24                                                   : in    std_logic;
          line_6_21                                                   : in    std_logic;
          line_6_10                                                   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11 : out   std_logic;
          MSS_READY                                                   : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                        : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE    : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                         : in    std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY                  : in    std_logic;
          hready_m_xhdl344_7                                          : out   std_logic;
          N_225                                                       : out   std_logic;
          N_276                                                       : out   std_logic;
          N_259                                                       : out   std_logic;
          N_243                                                       : out   std_logic;
          N_236                                                       : out   std_logic;
          N_235                                                       : out   std_logic;
          N_277                                                       : out   std_logic;
          N_255                                                       : out   std_logic;
          N_241                                                       : out   std_logic;
          N_242                                                       : out   std_logic;
          N_244                                                       : out   std_logic;
          N_246                                                       : out   std_logic;
          N_247                                                       : out   std_logic;
          N_256                                                       : out   std_logic;
          N_257                                                       : out   std_logic;
          N_258                                                       : out   std_logic;
          ren_pos                                                     : in    std_logic;
          hready_m_xhdl343_10                                         : out   std_logic;
          hready_m_xhdl343_11                                         : out   std_logic;
          N_120                                                       : out   std_logic;
          N_216                                                       : in    std_logic;
          N_215                                                       : in    std_logic;
          hready_m_xhdl345                                            : out   std_logic;
          N_335                                                       : in    std_logic;
          N_214                                                       : in    std_logic;
          N_305                                                       : in    std_logic;
          N_206                                                       : out   std_logic;
          N_508                                                       : in    std_logic;
          N_478_i_0                                                   : out   std_logic;
          N_507                                                       : in    std_logic;
          N_477_i_0                                                   : out   std_logic;
          N_479_i_0                                                   : out   std_logic;
          N_480_i_0                                                   : out   std_logic;
          N_481_i_0                                                   : out   std_logic;
          un8_hreadyin_i_0                                            : in    std_logic;
          N_9_i_0                                                     : out   std_logic;
          N_226                                                       : out   std_logic;
          defSlaveSMNextState                                         : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                     : in    std_logic;
          N_63_i_0                                                    : out   std_logic;
          N_62_i_0                                                    : out   std_logic;
          N_60_i_0                                                    : out   std_logic;
          N_98_i_0                                                    : out   std_logic;
          N_96_i_0                                                    : out   std_logic;
          N_94_i_0                                                    : out   std_logic;
          N_92_i_0                                                    : out   std_logic;
          N_90_i_0                                                    : out   std_logic;
          N_88_i_0                                                    : out   std_logic;
          N_86_i_0                                                    : out   std_logic;
          N_84_i_0                                                    : out   std_logic;
          N_82_i_0                                                    : out   std_logic;
          N_80_i_0                                                    : out   std_logic;
          N_78_i_0                                                    : out   std_logic;
          N_76_i_0                                                    : out   std_logic;
          N_74_i_0                                                    : out   std_logic;
          N_72_i_0                                                    : out   std_logic;
          N_70_i_0                                                    : out   std_logic;
          N_68_i_0                                                    : out   std_logic;
          N_66_i_0                                                    : out   std_logic;
          N_64_i_0                                                    : out   std_logic;
          N_58_i_0                                                    : out   std_logic;
          N_56_i_0                                                    : out   std_logic;
          N_54_i_0                                                    : out   std_logic;
          N_52_i_0                                                    : out   std_logic;
          N_50_i_0                                                    : out   std_logic;
          N_48_i_0                                                    : out   std_logic;
          N_46_i_0                                                    : out   std_logic;
          N_44_i_0                                                    : out   std_logic;
          N_42_i_0                                                    : out   std_logic;
          N_40_i_0                                                    : out   std_logic;
          N_38_i_0                                                    : out   std_logic;
          HTRANS_i_a2_0_0                                             : out   std_logic;
          N_271                                                       : in    std_logic;
          N_157_i_i_o2_0                                              : out   std_logic;
          N_157_i_i_o2_0_out                                          : out   std_logic;
          hsel2_i_4                                                   : out   std_logic;
          N_196_i_0                                                   : out   std_logic;
          N_195_i_0                                                   : out   std_logic;
          N_194_i_0                                                   : out   std_logic;
          N_65_i_0                                                    : out   std_logic;
          N_67_i_0                                                    : out   std_logic;
          N_110_i_0                                                   : out   std_logic;
          N_112_i_0                                                   : out   std_logic;
          N_114_i_0                                                   : out   std_logic;
          N_116_i_0                                                   : out   std_logic;
          N_69_i_0                                                    : out   std_logic;
          N_71_i_0                                                    : out   std_logic;
          N_73_i_0                                                    : out   std_logic;
          N_75_i_0                                                    : out   std_logic;
          N_77_i_0                                                    : out   std_logic;
          N_83_i_0                                                    : out   std_logic;
          N_85_i_0                                                    : out   std_logic;
          N_133_i_0                                                   : out   std_logic;
          N_87_i_0                                                    : out   std_logic;
          N_89_i_0                                                    : out   std_logic;
          N_140_i_0                                                   : out   std_logic;
          N_91_i_0                                                    : out   std_logic;
          N_93_i_0                                                    : out   std_logic;
          N_95_i_0                                                    : out   std_logic;
          N_97_i_0                                                    : out   std_logic;
          N_99_i_0                                                    : out   std_logic;
          N_152_i_0                                                   : out   std_logic;
          N_101_i_0                                                   : out   std_logic;
          N_156_i_0                                                   : out   std_logic;
          N_158_i_0                                                   : out   std_logic;
          N_103_i_0                                                   : out   std_logic;
          N_105_i_0                                                   : out   std_logic;
          N_107_i_0                                                   : out   std_logic;
          N_168_i_0                                                   : out   std_logic;
          N_109_i_0                                                   : out   std_logic;
          N_111_i_0                                                   : out   std_logic;
          N_218_i_0                                                   : out   std_logic;
          N_217_i_0                                                   : out   std_logic;
          N_203_i_0                                                   : out   std_logic
        );

end COREAHBLITE_MATRIX4X16;

architecture DEF_ARCH of COREAHBLITE_MATRIX4X16 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVESTAGE_0
    port( masterDataInProg                                         : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA : in    std_logic_vector(31 downto 0) := (others => 'U');
          arbRegSMCurrentState_ns_i_0                              : out   std_logic_vector(1 to 1);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR  : in    std_logic_vector(5 downto 3) := (others => 'U');
          regHADDR                                                 : in    std_logic_vector(5 downto 3) := (others => 'U');
          MSS_READY                                                : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                     : in    std_logic := 'U';
          CertificationSystem_sb_0_AHBmslave5_HREADY               : in    std_logic := 'U';
          N_65_i_0                                                 : out   std_logic;
          N_67_i_0                                                 : out   std_logic;
          N_110_i_0                                                : out   std_logic;
          N_112_i_0                                                : out   std_logic;
          N_114_i_0                                                : out   std_logic;
          N_116_i_0                                                : out   std_logic;
          N_69_i_0                                                 : out   std_logic;
          N_71_i_0                                                 : out   std_logic;
          N_73_i_0                                                 : out   std_logic;
          N_75_i_0                                                 : out   std_logic;
          N_77_i_0                                                 : out   std_logic;
          N_83_i_0                                                 : out   std_logic;
          N_85_i_0                                                 : out   std_logic;
          N_133_i_0                                                : out   std_logic;
          N_87_i_0                                                 : out   std_logic;
          N_89_i_0                                                 : out   std_logic;
          N_140_i_0                                                : out   std_logic;
          N_91_i_0                                                 : out   std_logic;
          N_93_i_0                                                 : out   std_logic;
          N_95_i_0                                                 : out   std_logic;
          N_97_i_0                                                 : out   std_logic;
          N_99_i_0                                                 : out   std_logic;
          N_152_i_0                                                : out   std_logic;
          N_101_i_0                                                : out   std_logic;
          N_156_i_0                                                : out   std_logic;
          N_158_i_0                                                : out   std_logic;
          N_103_i_0                                                : out   std_logic;
          N_105_i_0                                                : out   std_logic;
          N_107_i_0                                                : out   std_logic;
          N_168_i_0                                                : out   std_logic;
          N_109_i_0                                                : out   std_logic;
          N_111_i_0                                                : out   std_logic;
          N_127                                                    : in    std_logic := 'U';
          N_120                                                    : in    std_logic := 'U';
          N_226                                                    : out   std_logic;
          masterRegAddrSel                                         : in    std_logic := 'U';
          N_218_i_0                                                : out   std_logic;
          N_217_i_0                                                : out   std_logic;
          N_203_i_0                                                : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVESTAGE_1
    port( masterDataInProg                                          : out   std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA  : in    std_logic_vector(31 downto 0) := (others => 'U');
          xhdl1221                                                  : in    std_logic_vector(3 to 3) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HADDR                            : out   std_logic_vector(11 to 11);
          arbRegSMCurrentState_13                                   : out   std_logic;
          arbRegSMCurrentState_12                                   : out   std_logic;
          arbRegSMCurrentState_8                                    : out   std_logic;
          arbRegSMCurrentState_4                                    : out   std_logic;
          arbRegSMCurrentState_0                                    : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0 : in    std_logic := 'U';
          regHADDR_8                                                : in    std_logic := 'U';
          regHADDR_2                                                : in    std_logic := 'U';
          regHADDR_1                                                : in    std_logic := 'U';
          regHADDR_0                                                : in    std_logic := 'U';
          MSS_READY                                                 : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                      : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                   : in    std_logic := 'U';
          N_63_i_0                                                  : out   std_logic;
          N_62_i_0                                                  : out   std_logic;
          N_60_i_0                                                  : out   std_logic;
          N_98_i_0                                                  : out   std_logic;
          N_96_i_0                                                  : out   std_logic;
          N_94_i_0                                                  : out   std_logic;
          N_92_i_0                                                  : out   std_logic;
          N_90_i_0                                                  : out   std_logic;
          N_88_i_0                                                  : out   std_logic;
          N_86_i_0                                                  : out   std_logic;
          N_84_i_0                                                  : out   std_logic;
          N_82_i_0                                                  : out   std_logic;
          N_80_i_0                                                  : out   std_logic;
          N_78_i_0                                                  : out   std_logic;
          N_76_i_0                                                  : out   std_logic;
          N_74_i_0                                                  : out   std_logic;
          N_72_i_0                                                  : out   std_logic;
          N_70_i_0                                                  : out   std_logic;
          N_68_i_0                                                  : out   std_logic;
          N_66_i_0                                                  : out   std_logic;
          N_64_i_0                                                  : out   std_logic;
          N_58_i_0                                                  : out   std_logic;
          N_56_i_0                                                  : out   std_logic;
          N_54_i_0                                                  : out   std_logic;
          N_52_i_0                                                  : out   std_logic;
          N_50_i_0                                                  : out   std_logic;
          N_48_i_0                                                  : out   std_logic;
          N_46_i_0                                                  : out   std_logic;
          N_44_i_0                                                  : out   std_logic;
          N_42_i_0                                                  : out   std_logic;
          N_40_i_0                                                  : out   std_logic;
          N_38_i_0                                                  : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                       : in    std_logic := 'U';
          hready_m_xhdl345                                          : in    std_logic := 'U';
          un1_SDATASELInt_1                                         : in    std_logic := 'U';
          HTRANS_i_a2_0_0                                           : out   std_logic;
          N_271                                                     : in    std_logic := 'U';
          N_120                                                     : in    std_logic := 'U';
          N_225                                                     : in    std_logic := 'U';
          N_157_i_i_o2_0                                            : out   std_logic;
          N_148                                                     : in    std_logic := 'U';
          N_138                                                     : in    std_logic := 'U';
          N_149                                                     : in    std_logic := 'U';
          N_157_i_i_o2_0_out                                        : out   std_logic;
          hsel2_i_4                                                 : out   std_logic;
          N_135                                                     : in    std_logic := 'U';
          masterRegAddrSel                                          : in    std_logic := 'U';
          N_196_i_0                                                 : out   std_logic;
          N_195_i_0                                                 : out   std_logic;
          N_194_i_0                                                 : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MASTERSTAGE_1_1_0_40_0
    port( xhdl1221                                                    : out   std_logic_vector(3 to 3);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE     : in    std_logic_vector(1 downto 0) := (others => 'U');
          masterDataInProg                                            : in    std_logic_vector(0 to 0) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS    : in    std_logic_vector(1 to 1) := (others => 'U');
          result_addr_net_0                                           : in    std_logic_vector(3 downto 0) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP     : out   std_logic_vector(0 to 0);
          masterDataInProg_0                                          : in    std_logic_vector(0 to 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HRDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          line_7                                                      : in    std_logic_vector(2 downto 1) := (others => 'U');
          arbRegSMCurrentState_ns_i_0                                 : in    std_logic_vector(1 to 1) := (others => 'U');
          xhdl1222_0                                                  : out   std_logic;
          xhdl1222_2                                                  : out   std_logic;
          SDATASELInt_0                                               : out   std_logic;
          SDATASELInt_1                                               : out   std_logic;
          SDATASELInt_2                                               : out   std_logic;
          SDATASELInt_4                                               : out   std_logic;
          SDATASELInt_6                                               : out   std_logic;
          SDATASELInt_7                                               : out   std_logic;
          SDATASELInt_8                                               : out   std_logic;
          SDATASELInt_9                                               : out   std_logic;
          SDATASELInt_10                                              : out   std_logic;
          SDATASELInt_11                                              : out   std_logic;
          SDATASELInt_12                                              : out   std_logic;
          SDATASELInt_13                                              : out   std_logic;
          regHADDR_11                                                 : out   std_logic;
          regHADDR_3                                                  : out   std_logic;
          regHADDR_4                                                  : out   std_logic;
          regHADDR_5                                                  : out   std_logic;
          arbRegSMCurrentState_13                                     : in    std_logic := 'U';
          arbRegSMCurrentState_12                                     : in    std_logic := 'U';
          arbRegSMCurrentState_8                                      : in    std_logic := 'U';
          arbRegSMCurrentState_4                                      : in    std_logic := 'U';
          arbRegSMCurrentState_0                                      : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31  : in    std_logic := 'U';
          line_13                                                     : in    std_logic := 'U';
          line_10                                                     : in    std_logic := 'U';
          line_21                                                     : in    std_logic := 'U';
          line_24                                                     : in    std_logic := 'U';
          line_18                                                     : in    std_logic := 'U';
          line_23                                                     : in    std_logic := 'U';
          line_16                                                     : in    std_logic := 'U';
          line_28                                                     : in    std_logic := 'U';
          line_9                                                      : in    std_logic := 'U';
          line_3_d0                                                   : in    std_logic := 'U';
          line_5_d0                                                   : in    std_logic := 'U';
          line_15                                                     : in    std_logic := 'U';
          line_26                                                     : in    std_logic := 'U';
          line_14                                                     : in    std_logic := 'U';
          line_20                                                     : in    std_logic := 'U';
          line_2_d0                                                   : in    std_logic := 'U';
          line_25                                                     : in    std_logic := 'U';
          line_29                                                     : in    std_logic := 'U';
          line_19                                                     : in    std_logic := 'U';
          line_27                                                     : in    std_logic := 'U';
          line_30                                                     : in    std_logic := 'U';
          line_17                                                     : in    std_logic := 'U';
          line_8                                                      : in    std_logic := 'U';
          line_0_d0                                                   : in    std_logic := 'U';
          line_6_d0                                                   : in    std_logic := 'U';
          line_1_d0                                                   : in    std_logic := 'U';
          line_0_10                                                   : in    std_logic := 'U';
          line_0_21                                                   : in    std_logic := 'U';
          line_0_24                                                   : in    std_logic := 'U';
          line_0_18                                                   : in    std_logic := 'U';
          line_0_23                                                   : in    std_logic := 'U';
          line_0_16                                                   : in    std_logic := 'U';
          line_0_28                                                   : in    std_logic := 'U';
          line_0_9                                                    : in    std_logic := 'U';
          line_0_3                                                    : in    std_logic := 'U';
          line_0_5                                                    : in    std_logic := 'U';
          line_0_15                                                   : in    std_logic := 'U';
          line_0_26                                                   : in    std_logic := 'U';
          line_0_14                                                   : in    std_logic := 'U';
          line_0_20                                                   : in    std_logic := 'U';
          line_0_2                                                    : in    std_logic := 'U';
          line_0_25                                                   : in    std_logic := 'U';
          line_0_29                                                   : in    std_logic := 'U';
          line_0_19                                                   : in    std_logic := 'U';
          line_0_27                                                   : in    std_logic := 'U';
          line_0_30                                                   : in    std_logic := 'U';
          line_0_17                                                   : in    std_logic := 'U';
          line_0_8                                                    : in    std_logic := 'U';
          line_0_0                                                    : in    std_logic := 'U';
          line_0_1                                                    : in    std_logic := 'U';
          line_0_6                                                    : in    std_logic := 'U';
          line_0_13                                                   : in    std_logic := 'U';
          line_1_10                                                   : in    std_logic := 'U';
          line_1_21                                                   : in    std_logic := 'U';
          line_1_24                                                   : in    std_logic := 'U';
          line_1_18                                                   : in    std_logic := 'U';
          line_1_23                                                   : in    std_logic := 'U';
          line_1_16                                                   : in    std_logic := 'U';
          line_1_28                                                   : in    std_logic := 'U';
          line_1_9                                                    : in    std_logic := 'U';
          line_1_3                                                    : in    std_logic := 'U';
          line_1_5                                                    : in    std_logic := 'U';
          line_1_15                                                   : in    std_logic := 'U';
          line_1_26                                                   : in    std_logic := 'U';
          line_1_14                                                   : in    std_logic := 'U';
          line_1_20                                                   : in    std_logic := 'U';
          line_1_2                                                    : in    std_logic := 'U';
          line_1_25                                                   : in    std_logic := 'U';
          line_1_29                                                   : in    std_logic := 'U';
          line_1_19                                                   : in    std_logic := 'U';
          line_1_27                                                   : in    std_logic := 'U';
          line_1_30                                                   : in    std_logic := 'U';
          line_1_17                                                   : in    std_logic := 'U';
          line_1_8                                                    : in    std_logic := 'U';
          line_1_0                                                    : in    std_logic := 'U';
          line_1_1                                                    : in    std_logic := 'U';
          line_1_6                                                    : in    std_logic := 'U';
          line_1_13                                                   : in    std_logic := 'U';
          line_2_19                                                   : in    std_logic := 'U';
          line_2_27                                                   : in    std_logic := 'U';
          line_2_30                                                   : in    std_logic := 'U';
          line_2_17                                                   : in    std_logic := 'U';
          line_2_8                                                    : in    std_logic := 'U';
          line_2_10                                                   : in    std_logic := 'U';
          line_2_15                                                   : in    std_logic := 'U';
          line_2_26                                                   : in    std_logic := 'U';
          line_2_20                                                   : in    std_logic := 'U';
          line_2_0                                                    : in    std_logic := 'U';
          line_2_1                                                    : in    std_logic := 'U';
          line_2_29                                                   : in    std_logic := 'U';
          line_2_25                                                   : in    std_logic := 'U';
          line_2_2                                                    : in    std_logic := 'U';
          line_2_6                                                    : in    std_logic := 'U';
          line_2_13                                                   : in    std_logic := 'U';
          line_2_14                                                   : in    std_logic := 'U';
          line_2_5                                                    : in    std_logic := 'U';
          line_2_3                                                    : in    std_logic := 'U';
          line_2_9                                                    : in    std_logic := 'U';
          line_2_28                                                   : in    std_logic := 'U';
          line_2_16                                                   : in    std_logic := 'U';
          line_2_23                                                   : in    std_logic := 'U';
          line_2_18                                                   : in    std_logic := 'U';
          line_2_24                                                   : in    std_logic := 'U';
          line_2_21                                                   : in    std_logic := 'U';
          line_3_19                                                   : in    std_logic := 'U';
          line_3_17                                                   : in    std_logic := 'U';
          line_3_8                                                    : in    std_logic := 'U';
          line_3_0                                                    : in    std_logic := 'U';
          line_3_1                                                    : in    std_logic := 'U';
          line_3_29                                                   : in    std_logic := 'U';
          line_3_25                                                   : in    std_logic := 'U';
          line_3_2                                                    : in    std_logic := 'U';
          line_3_20                                                   : in    std_logic := 'U';
          line_3_6                                                    : in    std_logic := 'U';
          line_3_13                                                   : in    std_logic := 'U';
          line_3_14                                                   : in    std_logic := 'U';
          line_3_26                                                   : in    std_logic := 'U';
          line_3_15                                                   : in    std_logic := 'U';
          line_3_5                                                    : in    std_logic := 'U';
          line_3_3                                                    : in    std_logic := 'U';
          line_3_9                                                    : in    std_logic := 'U';
          line_3_28                                                   : in    std_logic := 'U';
          line_3_16                                                   : in    std_logic := 'U';
          line_3_23                                                   : in    std_logic := 'U';
          line_3_18                                                   : in    std_logic := 'U';
          line_3_24                                                   : in    std_logic := 'U';
          line_3_21                                                   : in    std_logic := 'U';
          line_3_10                                                   : in    std_logic := 'U';
          SHA256_Module_0_data_out_5                                  : in    std_logic := 'U';
          SHA256_Module_0_data_out_13                                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_12                                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_8                                  : in    std_logic := 'U';
          SHA256_Module_0_data_out_23                                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_0                                  : in    std_logic := 'U';
          line_4_19                                                   : in    std_logic := 'U';
          line_4_17                                                   : in    std_logic := 'U';
          line_4_8                                                    : in    std_logic := 'U';
          line_4_0                                                    : in    std_logic := 'U';
          line_4_1                                                    : in    std_logic := 'U';
          line_4_29                                                   : in    std_logic := 'U';
          line_4_25                                                   : in    std_logic := 'U';
          line_4_2                                                    : in    std_logic := 'U';
          line_4_20                                                   : in    std_logic := 'U';
          line_4_14                                                   : in    std_logic := 'U';
          line_4_26                                                   : in    std_logic := 'U';
          line_4_15                                                   : in    std_logic := 'U';
          line_4_5                                                    : in    std_logic := 'U';
          line_4_3                                                    : in    std_logic := 'U';
          line_4_9                                                    : in    std_logic := 'U';
          line_4_28                                                   : in    std_logic := 'U';
          line_4_16                                                   : in    std_logic := 'U';
          line_4_23                                                   : in    std_logic := 'U';
          line_4_18                                                   : in    std_logic := 'U';
          line_4_24                                                   : in    std_logic := 'U';
          line_4_21                                                   : in    std_logic := 'U';
          line_4_10                                                   : in    std_logic := 'U';
          line_4_6                                                    : in    std_logic := 'U';
          line_4_13                                                   : in    std_logic := 'U';
          line_5_19                                                   : in    std_logic := 'U';
          line_5_17                                                   : in    std_logic := 'U';
          line_5_8                                                    : in    std_logic := 'U';
          line_5_0                                                    : in    std_logic := 'U';
          line_5_1                                                    : in    std_logic := 'U';
          line_5_29                                                   : in    std_logic := 'U';
          line_5_25                                                   : in    std_logic := 'U';
          line_5_2                                                    : in    std_logic := 'U';
          line_5_20                                                   : in    std_logic := 'U';
          line_5_6                                                    : in    std_logic := 'U';
          line_5_13                                                   : in    std_logic := 'U';
          line_5_14                                                   : in    std_logic := 'U';
          line_5_26                                                   : in    std_logic := 'U';
          line_5_15                                                   : in    std_logic := 'U';
          line_5_5                                                    : in    std_logic := 'U';
          line_5_3                                                    : in    std_logic := 'U';
          line_5_9                                                    : in    std_logic := 'U';
          line_5_28                                                   : in    std_logic := 'U';
          line_5_16                                                   : in    std_logic := 'U';
          line_5_23                                                   : in    std_logic := 'U';
          line_5_18                                                   : in    std_logic := 'U';
          line_5_24                                                   : in    std_logic := 'U';
          line_5_21                                                   : in    std_logic := 'U';
          line_5_10                                                   : in    std_logic := 'U';
          line_6_19                                                   : in    std_logic := 'U';
          line_6_17                                                   : in    std_logic := 'U';
          line_6_8                                                    : in    std_logic := 'U';
          line_6_0                                                    : in    std_logic := 'U';
          line_6_1                                                    : in    std_logic := 'U';
          line_6_29                                                   : in    std_logic := 'U';
          line_6_25                                                   : in    std_logic := 'U';
          line_6_2                                                    : in    std_logic := 'U';
          line_6_20                                                   : in    std_logic := 'U';
          line_6_6                                                    : in    std_logic := 'U';
          line_6_13                                                   : in    std_logic := 'U';
          line_6_14                                                   : in    std_logic := 'U';
          line_6_26                                                   : in    std_logic := 'U';
          line_6_15                                                   : in    std_logic := 'U';
          line_6_5                                                    : in    std_logic := 'U';
          line_6_3                                                    : in    std_logic := 'U';
          line_6_9                                                    : in    std_logic := 'U';
          line_6_28                                                   : in    std_logic := 'U';
          line_6_16                                                   : in    std_logic := 'U';
          line_6_23                                                   : in    std_logic := 'U';
          line_6_18                                                   : in    std_logic := 'U';
          line_6_24                                                   : in    std_logic := 'U';
          line_6_21                                                   : in    std_logic := 'U';
          line_6_10                                                   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11 : out   std_logic;
          MSS_READY                                                   : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                        : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE    : in    std_logic := 'U';
          masterRegAddrSel                                            : out   std_logic;
          N_138                                                       : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                         : in    std_logic := 'U';
          N_148                                                       : out   std_logic;
          N_135                                                       : out   std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY                  : in    std_logic := 'U';
          hready_m_xhdl344_7                                          : out   std_logic;
          N_225                                                       : out   std_logic;
          N_149                                                       : out   std_logic;
          N_276                                                       : out   std_logic;
          N_259                                                       : out   std_logic;
          N_243                                                       : out   std_logic;
          N_236                                                       : out   std_logic;
          N_235                                                       : out   std_logic;
          N_277                                                       : out   std_logic;
          N_255                                                       : out   std_logic;
          N_241                                                       : out   std_logic;
          N_242                                                       : out   std_logic;
          N_244                                                       : out   std_logic;
          N_246                                                       : out   std_logic;
          N_247                                                       : out   std_logic;
          N_256                                                       : out   std_logic;
          N_257                                                       : out   std_logic;
          N_258                                                       : out   std_logic;
          ren_pos                                                     : in    std_logic := 'U';
          hready_m_xhdl343_10                                         : out   std_logic;
          hready_m_xhdl343_11                                         : out   std_logic;
          N_120                                                       : out   std_logic;
          N_127                                                       : out   std_logic;
          N_216                                                       : in    std_logic := 'U';
          N_215                                                       : in    std_logic := 'U';
          hready_m_xhdl345                                            : out   std_logic;
          un1_SDATASELInt_1                                           : out   std_logic;
          N_335                                                       : in    std_logic := 'U';
          N_214                                                       : in    std_logic := 'U';
          N_305                                                       : in    std_logic := 'U';
          N_206                                                       : out   std_logic;
          N_508                                                       : in    std_logic := 'U';
          N_478_i_0                                                   : out   std_logic;
          N_507                                                       : in    std_logic := 'U';
          N_477_i_0                                                   : out   std_logic;
          N_479_i_0                                                   : out   std_logic;
          N_480_i_0                                                   : out   std_logic;
          N_481_i_0                                                   : out   std_logic;
          un8_hreadyin_i_0                                            : in    std_logic := 'U';
          N_9_i_0                                                     : out   std_logic;
          N_226                                                       : in    std_logic := 'U';
          defSlaveSMNextState                                         : out   std_logic
        );
  end component;

    signal \xhdl1221[3]\, \regHADDR[11]\, \regHADDR[3]\, 
        \regHADDR[4]\, \regHADDR[5]\, \arbRegSMCurrentState_13\, 
        \arbRegSMCurrentState[14]\, \arbRegSMCurrentState[10]\, 
        \arbRegSMCurrentState[6]\, \arbRegSMCurrentState[2]\, 
        \masterDataInProg[0]\, \masterDataInProg_0[0]\, 
        \arbRegSMCurrentState_ns_i_0[1]\, masterRegAddrSel, N_138, 
        N_148, N_135, \N_225\, N_149, \N_120\, N_127, 
        \hready_m_xhdl345\, un1_SDATASELInt_1, \N_226\, GND_net_1, 
        VCC_net_1 : std_logic;

    for all : COREAHBLITE_SLAVESTAGE_0
	Use entity work.COREAHBLITE_SLAVESTAGE_0(DEF_ARCH);
    for all : COREAHBLITE_SLAVESTAGE_1
	Use entity work.COREAHBLITE_SLAVESTAGE_1(DEF_ARCH);
    for all : COREAHBLITE_MASTERSTAGE_1_1_0_40_0
	Use entity work.COREAHBLITE_MASTERSTAGE_1_1_0_40_0(DEF_ARCH);
begin 

    arbRegSMCurrentState_13 <= \arbRegSMCurrentState_13\;
    N_225 <= \N_225\;
    N_120 <= \N_120\;
    hready_m_xhdl345 <= \hready_m_xhdl345\;
    N_226 <= \N_226\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    slavestage_5 : COREAHBLITE_SLAVESTAGE_0
      port map(masterDataInProg(0) => \masterDataInProg[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        arbRegSMCurrentState_ns_i_0(1) => 
        \arbRegSMCurrentState_ns_i_0[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(5)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(4)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR(3)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        regHADDR(5) => \regHADDR[5]\, regHADDR(4) => 
        \regHADDR[4]\, regHADDR(3) => \regHADDR[3]\, MSS_READY
         => MSS_READY, CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, 
        CertificationSystem_sb_0_AHBmslave5_HREADY => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, N_65_i_0 => 
        N_65_i_0, N_67_i_0 => N_67_i_0, N_110_i_0 => N_110_i_0, 
        N_112_i_0 => N_112_i_0, N_114_i_0 => N_114_i_0, N_116_i_0
         => N_116_i_0, N_69_i_0 => N_69_i_0, N_71_i_0 => N_71_i_0, 
        N_73_i_0 => N_73_i_0, N_75_i_0 => N_75_i_0, N_77_i_0 => 
        N_77_i_0, N_83_i_0 => N_83_i_0, N_85_i_0 => N_85_i_0, 
        N_133_i_0 => N_133_i_0, N_87_i_0 => N_87_i_0, N_89_i_0
         => N_89_i_0, N_140_i_0 => N_140_i_0, N_91_i_0 => 
        N_91_i_0, N_93_i_0 => N_93_i_0, N_95_i_0 => N_95_i_0, 
        N_97_i_0 => N_97_i_0, N_99_i_0 => N_99_i_0, N_152_i_0 => 
        N_152_i_0, N_101_i_0 => N_101_i_0, N_156_i_0 => N_156_i_0, 
        N_158_i_0 => N_158_i_0, N_103_i_0 => N_103_i_0, N_105_i_0
         => N_105_i_0, N_107_i_0 => N_107_i_0, N_168_i_0 => 
        N_168_i_0, N_109_i_0 => N_109_i_0, N_111_i_0 => N_111_i_0, 
        N_127 => N_127, N_120 => \N_120\, N_226 => \N_226\, 
        masterRegAddrSel => masterRegAddrSel, N_218_i_0 => 
        N_218_i_0, N_217_i_0 => N_217_i_0, N_203_i_0 => N_203_i_0);
    
    slavestage_3 : COREAHBLITE_SLAVESTAGE_1
      port map(masterDataInProg(0) => \masterDataInProg_0[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        xhdl1221(3) => \xhdl1221[3]\, 
        CoreAHBLite_0_AHBmslave3_HADDR(11) => 
        CoreAHBLite_0_AHBmslave3_HADDR(11), 
        arbRegSMCurrentState_13 => \arbRegSMCurrentState_13\, 
        arbRegSMCurrentState_12 => \arbRegSMCurrentState[14]\, 
        arbRegSMCurrentState_8 => \arbRegSMCurrentState[10]\, 
        arbRegSMCurrentState_4 => \arbRegSMCurrentState[6]\, 
        arbRegSMCurrentState_0 => \arbRegSMCurrentState[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        regHADDR_8 => \regHADDR[11]\, regHADDR_2 => \regHADDR[5]\, 
        regHADDR_1 => \regHADDR[4]\, regHADDR_0 => \regHADDR[3]\, 
        MSS_READY => MSS_READY, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, N_63_i_0 => 
        N_63_i_0, N_62_i_0 => N_62_i_0, N_60_i_0 => N_60_i_0, 
        N_98_i_0 => N_98_i_0, N_96_i_0 => N_96_i_0, N_94_i_0 => 
        N_94_i_0, N_92_i_0 => N_92_i_0, N_90_i_0 => N_90_i_0, 
        N_88_i_0 => N_88_i_0, N_86_i_0 => N_86_i_0, N_84_i_0 => 
        N_84_i_0, N_82_i_0 => N_82_i_0, N_80_i_0 => N_80_i_0, 
        N_78_i_0 => N_78_i_0, N_76_i_0 => N_76_i_0, N_74_i_0 => 
        N_74_i_0, N_72_i_0 => N_72_i_0, N_70_i_0 => N_70_i_0, 
        N_68_i_0 => N_68_i_0, N_66_i_0 => N_66_i_0, N_64_i_0 => 
        N_64_i_0, N_58_i_0 => N_58_i_0, N_56_i_0 => N_56_i_0, 
        N_54_i_0 => N_54_i_0, N_52_i_0 => N_52_i_0, N_50_i_0 => 
        N_50_i_0, N_48_i_0 => N_48_i_0, N_46_i_0 => N_46_i_0, 
        N_44_i_0 => N_44_i_0, N_42_i_0 => N_42_i_0, N_40_i_0 => 
        N_40_i_0, N_38_i_0 => N_38_i_0, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, hready_m_xhdl345 => 
        \hready_m_xhdl345\, un1_SDATASELInt_1 => 
        un1_SDATASELInt_1, HTRANS_i_a2_0_0 => HTRANS_i_a2_0_0, 
        N_271 => N_271, N_120 => \N_120\, N_225 => \N_225\, 
        N_157_i_i_o2_0 => N_157_i_i_o2_0, N_148 => N_148, N_138
         => N_138, N_149 => N_149, N_157_i_i_o2_0_out => 
        N_157_i_i_o2_0_out, hsel2_i_4 => hsel2_i_4, N_135 => 
        N_135, masterRegAddrSel => masterRegAddrSel, N_196_i_0
         => N_196_i_0, N_195_i_0 => N_195_i_0, N_194_i_0 => 
        N_194_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    masterstage_0 : COREAHBLITE_MASTERSTAGE_1_1_0_40_0
      port map(xhdl1221(3) => \xhdl1221[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0), 
        masterDataInProg(0) => \masterDataInProg[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        result_addr_net_0(3) => result_addr_net_0(3), 
        result_addr_net_0(2) => result_addr_net_0(2), 
        result_addr_net_0(1) => result_addr_net_0(1), 
        result_addr_net_0(0) => result_addr_net_0(0), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        masterDataInProg_0(0) => \masterDataInProg_0[0]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(31) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(31), 
        CoreAHBLite_0_AHBmslave3_HRDATA(30) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(30), 
        CoreAHBLite_0_AHBmslave3_HRDATA(29) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(29), 
        CoreAHBLite_0_AHBmslave3_HRDATA(28) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(28), 
        CoreAHBLite_0_AHBmslave3_HRDATA(27) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(27), 
        CoreAHBLite_0_AHBmslave3_HRDATA(26) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(26), 
        CoreAHBLite_0_AHBmslave3_HRDATA(25) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(25), 
        CoreAHBLite_0_AHBmslave3_HRDATA(24) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(24), 
        CoreAHBLite_0_AHBmslave3_HRDATA(23) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(23), 
        CoreAHBLite_0_AHBmslave3_HRDATA(22) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(22), 
        CoreAHBLite_0_AHBmslave3_HRDATA(21) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(21), 
        CoreAHBLite_0_AHBmslave3_HRDATA(20) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(20), 
        CoreAHBLite_0_AHBmslave3_HRDATA(19) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(19), 
        CoreAHBLite_0_AHBmslave3_HRDATA(18) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(18), 
        CoreAHBLite_0_AHBmslave3_HRDATA(17) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(17), 
        CoreAHBLite_0_AHBmslave3_HRDATA(16) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(16), 
        CoreAHBLite_0_AHBmslave3_HRDATA(15) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(15), 
        CoreAHBLite_0_AHBmslave3_HRDATA(14) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(14), 
        CoreAHBLite_0_AHBmslave3_HRDATA(13) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(13), 
        CoreAHBLite_0_AHBmslave3_HRDATA(12) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(12), 
        CoreAHBLite_0_AHBmslave3_HRDATA(11) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(11), 
        CoreAHBLite_0_AHBmslave3_HRDATA(10) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(10), 
        CoreAHBLite_0_AHBmslave3_HRDATA(9) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(9), 
        CoreAHBLite_0_AHBmslave3_HRDATA(8) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(8), 
        CoreAHBLite_0_AHBmslave3_HRDATA(7) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(7), 
        CoreAHBLite_0_AHBmslave3_HRDATA(6) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(6), 
        CoreAHBLite_0_AHBmslave3_HRDATA(5) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(5), 
        CoreAHBLite_0_AHBmslave3_HRDATA(4) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(4), 
        CoreAHBLite_0_AHBmslave3_HRDATA(3) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(3), 
        CoreAHBLite_0_AHBmslave3_HRDATA(2) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(2), 
        CoreAHBLite_0_AHBmslave3_HRDATA(1) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(1), 
        CoreAHBLite_0_AHBmslave3_HRDATA(0) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(0), line_7(2) => 
        line_7(2), line_7(1) => line_7(1), 
        arbRegSMCurrentState_ns_i_0(1) => 
        \arbRegSMCurrentState_ns_i_0[1]\, xhdl1222_0 => 
        xhdl1222_0, xhdl1222_2 => xhdl1222_2, SDATASELInt_0 => 
        SDATASELInt_0, SDATASELInt_1 => SDATASELInt_1, 
        SDATASELInt_2 => SDATASELInt_2, SDATASELInt_4 => 
        SDATASELInt_4, SDATASELInt_6 => SDATASELInt_6, 
        SDATASELInt_7 => SDATASELInt_7, SDATASELInt_8 => 
        SDATASELInt_8, SDATASELInt_9 => SDATASELInt_9, 
        SDATASELInt_10 => SDATASELInt_10, SDATASELInt_11 => 
        SDATASELInt_11, SDATASELInt_12 => SDATASELInt_12, 
        SDATASELInt_13 => SDATASELInt_13, regHADDR_11 => 
        \regHADDR[11]\, regHADDR_3 => \regHADDR[3]\, regHADDR_4
         => \regHADDR[4]\, regHADDR_5 => \regHADDR[5]\, 
        arbRegSMCurrentState_13 => \arbRegSMCurrentState_13\, 
        arbRegSMCurrentState_12 => \arbRegSMCurrentState[14]\, 
        arbRegSMCurrentState_8 => \arbRegSMCurrentState[10]\, 
        arbRegSMCurrentState_4 => \arbRegSMCurrentState[6]\, 
        arbRegSMCurrentState_0 => \arbRegSMCurrentState[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        line_13 => line_13, line_10 => line_10, line_21 => 
        line_21, line_24 => line_24, line_18 => line_18, line_23
         => line_23, line_16 => line_16, line_28 => line_28, 
        line_9 => line_9, line_3_d0 => line_3_d0, line_5_d0 => 
        line_5_d0, line_15 => line_15, line_26 => line_26, 
        line_14 => line_14, line_20 => line_20, line_2_d0 => 
        line_2_d0, line_25 => line_25, line_29 => line_29, 
        line_19 => line_19, line_27 => line_27, line_30 => 
        line_30, line_17 => line_17, line_8 => line_8, line_0_d0
         => line_0_d0, line_6_d0 => line_6_d0, line_1_d0 => 
        line_1_d0, line_0_10 => line_0_10, line_0_21 => line_0_21, 
        line_0_24 => line_0_24, line_0_18 => line_0_18, line_0_23
         => line_0_23, line_0_16 => line_0_16, line_0_28 => 
        line_0_28, line_0_9 => line_0_9, line_0_3 => line_0_3, 
        line_0_5 => line_0_5, line_0_15 => line_0_15, line_0_26
         => line_0_26, line_0_14 => line_0_14, line_0_20 => 
        line_0_20, line_0_2 => line_0_2, line_0_25 => line_0_25, 
        line_0_29 => line_0_29, line_0_19 => line_0_19, line_0_27
         => line_0_27, line_0_30 => line_0_30, line_0_17 => 
        line_0_17, line_0_8 => line_0_8, line_0_0 => line_0_0, 
        line_0_1 => line_0_1, line_0_6 => line_0_6, line_0_13 => 
        line_0_13, line_1_10 => line_1_10, line_1_21 => line_1_21, 
        line_1_24 => line_1_24, line_1_18 => line_1_18, line_1_23
         => line_1_23, line_1_16 => line_1_16, line_1_28 => 
        line_1_28, line_1_9 => line_1_9, line_1_3 => line_1_3, 
        line_1_5 => line_1_5, line_1_15 => line_1_15, line_1_26
         => line_1_26, line_1_14 => line_1_14, line_1_20 => 
        line_1_20, line_1_2 => line_1_2, line_1_25 => line_1_25, 
        line_1_29 => line_1_29, line_1_19 => line_1_19, line_1_27
         => line_1_27, line_1_30 => line_1_30, line_1_17 => 
        line_1_17, line_1_8 => line_1_8, line_1_0 => line_1_0, 
        line_1_1 => line_1_1, line_1_6 => line_1_6, line_1_13 => 
        line_1_13, line_2_19 => line_2_19, line_2_27 => line_2_27, 
        line_2_30 => line_2_30, line_2_17 => line_2_17, line_2_8
         => line_2_8, line_2_10 => line_2_10, line_2_15 => 
        line_2_15, line_2_26 => line_2_26, line_2_20 => line_2_20, 
        line_2_0 => line_2_0, line_2_1 => line_2_1, line_2_29 => 
        line_2_29, line_2_25 => line_2_25, line_2_2 => line_2_2, 
        line_2_6 => line_2_6, line_2_13 => line_2_13, line_2_14
         => line_2_14, line_2_5 => line_2_5, line_2_3 => line_2_3, 
        line_2_9 => line_2_9, line_2_28 => line_2_28, line_2_16
         => line_2_16, line_2_23 => line_2_23, line_2_18 => 
        line_2_18, line_2_24 => line_2_24, line_2_21 => line_2_21, 
        line_3_19 => line_3_19, line_3_17 => line_3_17, line_3_8
         => line_3_8, line_3_0 => line_3_0, line_3_1 => line_3_1, 
        line_3_29 => line_3_29, line_3_25 => line_3_25, line_3_2
         => line_3_2, line_3_20 => line_3_20, line_3_6 => 
        line_3_6, line_3_13 => line_3_13, line_3_14 => line_3_14, 
        line_3_26 => line_3_26, line_3_15 => line_3_15, line_3_5
         => line_3_5, line_3_3 => line_3_3, line_3_9 => line_3_9, 
        line_3_28 => line_3_28, line_3_16 => line_3_16, line_3_23
         => line_3_23, line_3_18 => line_3_18, line_3_24 => 
        line_3_24, line_3_21 => line_3_21, line_3_10 => line_3_10, 
        SHA256_Module_0_data_out_5 => SHA256_Module_0_data_out_5, 
        SHA256_Module_0_data_out_13 => 
        SHA256_Module_0_data_out_13, SHA256_Module_0_data_out_12
         => SHA256_Module_0_data_out_12, 
        SHA256_Module_0_data_out_8 => SHA256_Module_0_data_out_8, 
        SHA256_Module_0_data_out_23 => 
        SHA256_Module_0_data_out_23, SHA256_Module_0_data_out_0
         => SHA256_Module_0_data_out_0, line_4_19 => line_4_19, 
        line_4_17 => line_4_17, line_4_8 => line_4_8, line_4_0
         => line_4_0, line_4_1 => line_4_1, line_4_29 => 
        line_4_29, line_4_25 => line_4_25, line_4_2 => line_4_2, 
        line_4_20 => line_4_20, line_4_14 => line_4_14, line_4_26
         => line_4_26, line_4_15 => line_4_15, line_4_5 => 
        line_4_5, line_4_3 => line_4_3, line_4_9 => line_4_9, 
        line_4_28 => line_4_28, line_4_16 => line_4_16, line_4_23
         => line_4_23, line_4_18 => line_4_18, line_4_24 => 
        line_4_24, line_4_21 => line_4_21, line_4_10 => line_4_10, 
        line_4_6 => line_4_6, line_4_13 => line_4_13, line_5_19
         => line_5_19, line_5_17 => line_5_17, line_5_8 => 
        line_5_8, line_5_0 => line_5_0, line_5_1 => line_5_1, 
        line_5_29 => line_5_29, line_5_25 => line_5_25, line_5_2
         => line_5_2, line_5_20 => line_5_20, line_5_6 => 
        line_5_6, line_5_13 => line_5_13, line_5_14 => line_5_14, 
        line_5_26 => line_5_26, line_5_15 => line_5_15, line_5_5
         => line_5_5, line_5_3 => line_5_3, line_5_9 => line_5_9, 
        line_5_28 => line_5_28, line_5_16 => line_5_16, line_5_23
         => line_5_23, line_5_18 => line_5_18, line_5_24 => 
        line_5_24, line_5_21 => line_5_21, line_5_10 => line_5_10, 
        line_6_19 => line_6_19, line_6_17 => line_6_17, line_6_8
         => line_6_8, line_6_0 => line_6_0, line_6_1 => line_6_1, 
        line_6_29 => line_6_29, line_6_25 => line_6_25, line_6_2
         => line_6_2, line_6_20 => line_6_20, line_6_6 => 
        line_6_6, line_6_13 => line_6_13, line_6_14 => line_6_14, 
        line_6_26 => line_6_26, line_6_15 => line_6_15, line_6_5
         => line_6_5, line_6_3 => line_6_3, line_6_9 => line_6_9, 
        line_6_28 => line_6_28, line_6_16 => line_6_16, line_6_23
         => line_6_23, line_6_18 => line_6_18, line_6_24 => 
        line_6_24, line_6_21 => line_6_21, line_6_10 => line_6_10, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11, 
        MSS_READY => MSS_READY, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        masterRegAddrSel => masterRegAddrSel, N_138 => N_138, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, N_148 => N_148, 
        N_135 => N_135, 
        CertificationSystem_sb_0_AHBmslave5_HREADY => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, 
        hready_m_xhdl344_7 => hready_m_xhdl344_7, N_225 => 
        \N_225\, N_149 => N_149, N_276 => N_276, N_259 => N_259, 
        N_243 => N_243, N_236 => N_236, N_235 => N_235, N_277 => 
        N_277, N_255 => N_255, N_241 => N_241, N_242 => N_242, 
        N_244 => N_244, N_246 => N_246, N_247 => N_247, N_256 => 
        N_256, N_257 => N_257, N_258 => N_258, ren_pos => ren_pos, 
        hready_m_xhdl343_10 => hready_m_xhdl343_10, 
        hready_m_xhdl343_11 => hready_m_xhdl343_11, N_120 => 
        \N_120\, N_127 => N_127, N_216 => N_216, N_215 => N_215, 
        hready_m_xhdl345 => \hready_m_xhdl345\, un1_SDATASELInt_1
         => un1_SDATASELInt_1, N_335 => N_335, N_214 => N_214, 
        N_305 => N_305, N_206 => N_206, N_508 => N_508, N_478_i_0
         => N_478_i_0, N_507 => N_507, N_477_i_0 => N_477_i_0, 
        N_479_i_0 => N_479_i_0, N_480_i_0 => N_480_i_0, N_481_i_0
         => N_481_i_0, un8_hreadyin_i_0 => un8_hreadyin_i_0, 
        N_9_i_0 => N_9_i_0, N_226 => \N_226\, defSlaveSMNextState
         => defSlaveSMNextState);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLite is

    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE     : in    std_logic_vector(1 downto 0);
          arbRegSMCurrentState                                        : out   std_logic_vector(15 to 15);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS    : in    std_logic_vector(1 to 1);
          result_addr_net_0                                           : in    std_logic_vector(3 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP     : out   std_logic_vector(0 to 0);
          CoreAHBLite_0_AHBmslave3_HRDATA                             : in    std_logic_vector(31 downto 0);
          line_7                                                      : in    std_logic_vector(2 downto 1);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA    : in    std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave3_HADDR                              : out   std_logic_vector(11 to 11);
          xhdl1222_0                                                  : out   std_logic;
          xhdl1222_2                                                  : out   std_logic;
          SDATASELInt_0                                               : out   std_logic;
          SDATASELInt_1                                               : out   std_logic;
          SDATASELInt_2                                               : out   std_logic;
          SDATASELInt_4                                               : out   std_logic;
          SDATASELInt_6                                               : out   std_logic;
          SDATASELInt_7                                               : out   std_logic;
          SDATASELInt_8                                               : out   std_logic;
          SDATASELInt_9                                               : out   std_logic;
          SDATASELInt_10                                              : out   std_logic;
          SDATASELInt_11                                              : out   std_logic;
          SDATASELInt_12                                              : out   std_logic;
          SDATASELInt_13                                              : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31  : in    std_logic;
          line_13                                                     : in    std_logic;
          line_10                                                     : in    std_logic;
          line_21                                                     : in    std_logic;
          line_24                                                     : in    std_logic;
          line_18                                                     : in    std_logic;
          line_23                                                     : in    std_logic;
          line_16                                                     : in    std_logic;
          line_28                                                     : in    std_logic;
          line_9                                                      : in    std_logic;
          line_3_d0                                                   : in    std_logic;
          line_5_d0                                                   : in    std_logic;
          line_15                                                     : in    std_logic;
          line_26                                                     : in    std_logic;
          line_14                                                     : in    std_logic;
          line_20                                                     : in    std_logic;
          line_2_d0                                                   : in    std_logic;
          line_25                                                     : in    std_logic;
          line_29                                                     : in    std_logic;
          line_19                                                     : in    std_logic;
          line_27                                                     : in    std_logic;
          line_30                                                     : in    std_logic;
          line_17                                                     : in    std_logic;
          line_8                                                      : in    std_logic;
          line_0_d0                                                   : in    std_logic;
          line_6_d0                                                   : in    std_logic;
          line_1_d0                                                   : in    std_logic;
          line_0_10                                                   : in    std_logic;
          line_0_21                                                   : in    std_logic;
          line_0_24                                                   : in    std_logic;
          line_0_18                                                   : in    std_logic;
          line_0_23                                                   : in    std_logic;
          line_0_16                                                   : in    std_logic;
          line_0_28                                                   : in    std_logic;
          line_0_9                                                    : in    std_logic;
          line_0_3                                                    : in    std_logic;
          line_0_5                                                    : in    std_logic;
          line_0_15                                                   : in    std_logic;
          line_0_26                                                   : in    std_logic;
          line_0_14                                                   : in    std_logic;
          line_0_20                                                   : in    std_logic;
          line_0_2                                                    : in    std_logic;
          line_0_25                                                   : in    std_logic;
          line_0_29                                                   : in    std_logic;
          line_0_19                                                   : in    std_logic;
          line_0_27                                                   : in    std_logic;
          line_0_30                                                   : in    std_logic;
          line_0_17                                                   : in    std_logic;
          line_0_8                                                    : in    std_logic;
          line_0_0                                                    : in    std_logic;
          line_0_1                                                    : in    std_logic;
          line_0_6                                                    : in    std_logic;
          line_0_13                                                   : in    std_logic;
          line_1_10                                                   : in    std_logic;
          line_1_21                                                   : in    std_logic;
          line_1_24                                                   : in    std_logic;
          line_1_18                                                   : in    std_logic;
          line_1_23                                                   : in    std_logic;
          line_1_16                                                   : in    std_logic;
          line_1_28                                                   : in    std_logic;
          line_1_9                                                    : in    std_logic;
          line_1_3                                                    : in    std_logic;
          line_1_5                                                    : in    std_logic;
          line_1_15                                                   : in    std_logic;
          line_1_26                                                   : in    std_logic;
          line_1_14                                                   : in    std_logic;
          line_1_20                                                   : in    std_logic;
          line_1_2                                                    : in    std_logic;
          line_1_25                                                   : in    std_logic;
          line_1_29                                                   : in    std_logic;
          line_1_19                                                   : in    std_logic;
          line_1_27                                                   : in    std_logic;
          line_1_30                                                   : in    std_logic;
          line_1_17                                                   : in    std_logic;
          line_1_8                                                    : in    std_logic;
          line_1_0                                                    : in    std_logic;
          line_1_1                                                    : in    std_logic;
          line_1_6                                                    : in    std_logic;
          line_1_13                                                   : in    std_logic;
          line_2_19                                                   : in    std_logic;
          line_2_27                                                   : in    std_logic;
          line_2_30                                                   : in    std_logic;
          line_2_17                                                   : in    std_logic;
          line_2_8                                                    : in    std_logic;
          line_2_10                                                   : in    std_logic;
          line_2_15                                                   : in    std_logic;
          line_2_26                                                   : in    std_logic;
          line_2_20                                                   : in    std_logic;
          line_2_0                                                    : in    std_logic;
          line_2_1                                                    : in    std_logic;
          line_2_29                                                   : in    std_logic;
          line_2_25                                                   : in    std_logic;
          line_2_2                                                    : in    std_logic;
          line_2_6                                                    : in    std_logic;
          line_2_13                                                   : in    std_logic;
          line_2_14                                                   : in    std_logic;
          line_2_5                                                    : in    std_logic;
          line_2_3                                                    : in    std_logic;
          line_2_9                                                    : in    std_logic;
          line_2_28                                                   : in    std_logic;
          line_2_16                                                   : in    std_logic;
          line_2_23                                                   : in    std_logic;
          line_2_18                                                   : in    std_logic;
          line_2_24                                                   : in    std_logic;
          line_2_21                                                   : in    std_logic;
          line_3_19                                                   : in    std_logic;
          line_3_17                                                   : in    std_logic;
          line_3_8                                                    : in    std_logic;
          line_3_0                                                    : in    std_logic;
          line_3_1                                                    : in    std_logic;
          line_3_29                                                   : in    std_logic;
          line_3_25                                                   : in    std_logic;
          line_3_2                                                    : in    std_logic;
          line_3_20                                                   : in    std_logic;
          line_3_6                                                    : in    std_logic;
          line_3_13                                                   : in    std_logic;
          line_3_14                                                   : in    std_logic;
          line_3_26                                                   : in    std_logic;
          line_3_15                                                   : in    std_logic;
          line_3_5                                                    : in    std_logic;
          line_3_3                                                    : in    std_logic;
          line_3_9                                                    : in    std_logic;
          line_3_28                                                   : in    std_logic;
          line_3_16                                                   : in    std_logic;
          line_3_23                                                   : in    std_logic;
          line_3_18                                                   : in    std_logic;
          line_3_24                                                   : in    std_logic;
          line_3_21                                                   : in    std_logic;
          line_3_10                                                   : in    std_logic;
          SHA256_Module_0_data_out_5                                  : in    std_logic;
          SHA256_Module_0_data_out_13                                 : in    std_logic;
          SHA256_Module_0_data_out_12                                 : in    std_logic;
          SHA256_Module_0_data_out_8                                  : in    std_logic;
          SHA256_Module_0_data_out_23                                 : in    std_logic;
          SHA256_Module_0_data_out_0                                  : in    std_logic;
          line_4_19                                                   : in    std_logic;
          line_4_17                                                   : in    std_logic;
          line_4_8                                                    : in    std_logic;
          line_4_0                                                    : in    std_logic;
          line_4_1                                                    : in    std_logic;
          line_4_29                                                   : in    std_logic;
          line_4_25                                                   : in    std_logic;
          line_4_2                                                    : in    std_logic;
          line_4_20                                                   : in    std_logic;
          line_4_14                                                   : in    std_logic;
          line_4_26                                                   : in    std_logic;
          line_4_15                                                   : in    std_logic;
          line_4_5                                                    : in    std_logic;
          line_4_3                                                    : in    std_logic;
          line_4_9                                                    : in    std_logic;
          line_4_28                                                   : in    std_logic;
          line_4_16                                                   : in    std_logic;
          line_4_23                                                   : in    std_logic;
          line_4_18                                                   : in    std_logic;
          line_4_24                                                   : in    std_logic;
          line_4_21                                                   : in    std_logic;
          line_4_10                                                   : in    std_logic;
          line_4_6                                                    : in    std_logic;
          line_4_13                                                   : in    std_logic;
          line_5_19                                                   : in    std_logic;
          line_5_17                                                   : in    std_logic;
          line_5_8                                                    : in    std_logic;
          line_5_0                                                    : in    std_logic;
          line_5_1                                                    : in    std_logic;
          line_5_29                                                   : in    std_logic;
          line_5_25                                                   : in    std_logic;
          line_5_2                                                    : in    std_logic;
          line_5_20                                                   : in    std_logic;
          line_5_6                                                    : in    std_logic;
          line_5_13                                                   : in    std_logic;
          line_5_14                                                   : in    std_logic;
          line_5_26                                                   : in    std_logic;
          line_5_15                                                   : in    std_logic;
          line_5_5                                                    : in    std_logic;
          line_5_3                                                    : in    std_logic;
          line_5_9                                                    : in    std_logic;
          line_5_28                                                   : in    std_logic;
          line_5_16                                                   : in    std_logic;
          line_5_23                                                   : in    std_logic;
          line_5_18                                                   : in    std_logic;
          line_5_24                                                   : in    std_logic;
          line_5_21                                                   : in    std_logic;
          line_5_10                                                   : in    std_logic;
          line_6_19                                                   : in    std_logic;
          line_6_17                                                   : in    std_logic;
          line_6_8                                                    : in    std_logic;
          line_6_0                                                    : in    std_logic;
          line_6_1                                                    : in    std_logic;
          line_6_29                                                   : in    std_logic;
          line_6_25                                                   : in    std_logic;
          line_6_2                                                    : in    std_logic;
          line_6_20                                                   : in    std_logic;
          line_6_6                                                    : in    std_logic;
          line_6_13                                                   : in    std_logic;
          line_6_14                                                   : in    std_logic;
          line_6_26                                                   : in    std_logic;
          line_6_15                                                   : in    std_logic;
          line_6_5                                                    : in    std_logic;
          line_6_3                                                    : in    std_logic;
          line_6_9                                                    : in    std_logic;
          line_6_28                                                   : in    std_logic;
          line_6_16                                                   : in    std_logic;
          line_6_23                                                   : in    std_logic;
          line_6_18                                                   : in    std_logic;
          line_6_24                                                   : in    std_logic;
          line_6_21                                                   : in    std_logic;
          line_6_10                                                   : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11 : out   std_logic;
          MSS_READY                                                   : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                        : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE    : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                         : in    std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY                  : in    std_logic;
          hready_m_xhdl344_7                                          : out   std_logic;
          N_225                                                       : out   std_logic;
          N_276                                                       : out   std_logic;
          N_259                                                       : out   std_logic;
          N_243                                                       : out   std_logic;
          N_236                                                       : out   std_logic;
          N_235                                                       : out   std_logic;
          N_277                                                       : out   std_logic;
          N_255                                                       : out   std_logic;
          N_241                                                       : out   std_logic;
          N_242                                                       : out   std_logic;
          N_244                                                       : out   std_logic;
          N_246                                                       : out   std_logic;
          N_247                                                       : out   std_logic;
          N_256                                                       : out   std_logic;
          N_257                                                       : out   std_logic;
          N_258                                                       : out   std_logic;
          ren_pos                                                     : in    std_logic;
          hready_m_xhdl343_10                                         : out   std_logic;
          hready_m_xhdl343_11                                         : out   std_logic;
          N_120                                                       : out   std_logic;
          N_216                                                       : in    std_logic;
          N_215                                                       : in    std_logic;
          hready_m_xhdl345                                            : out   std_logic;
          N_335                                                       : in    std_logic;
          N_214                                                       : in    std_logic;
          N_305                                                       : in    std_logic;
          N_206                                                       : out   std_logic;
          N_508                                                       : in    std_logic;
          N_478_i_0                                                   : out   std_logic;
          N_507                                                       : in    std_logic;
          N_477_i_0                                                   : out   std_logic;
          N_479_i_0                                                   : out   std_logic;
          N_480_i_0                                                   : out   std_logic;
          N_481_i_0                                                   : out   std_logic;
          un8_hreadyin_i_0                                            : in    std_logic;
          N_9_i_0                                                     : out   std_logic;
          N_226                                                       : out   std_logic;
          defSlaveSMNextState                                         : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                     : in    std_logic;
          N_63_i_0                                                    : out   std_logic;
          N_62_i_0                                                    : out   std_logic;
          N_60_i_0                                                    : out   std_logic;
          N_98_i_0                                                    : out   std_logic;
          N_96_i_0                                                    : out   std_logic;
          N_94_i_0                                                    : out   std_logic;
          N_92_i_0                                                    : out   std_logic;
          N_90_i_0                                                    : out   std_logic;
          N_88_i_0                                                    : out   std_logic;
          N_86_i_0                                                    : out   std_logic;
          N_84_i_0                                                    : out   std_logic;
          N_82_i_0                                                    : out   std_logic;
          N_80_i_0                                                    : out   std_logic;
          N_78_i_0                                                    : out   std_logic;
          N_76_i_0                                                    : out   std_logic;
          N_74_i_0                                                    : out   std_logic;
          N_72_i_0                                                    : out   std_logic;
          N_70_i_0                                                    : out   std_logic;
          N_68_i_0                                                    : out   std_logic;
          N_66_i_0                                                    : out   std_logic;
          N_64_i_0                                                    : out   std_logic;
          N_58_i_0                                                    : out   std_logic;
          N_56_i_0                                                    : out   std_logic;
          N_54_i_0                                                    : out   std_logic;
          N_52_i_0                                                    : out   std_logic;
          N_50_i_0                                                    : out   std_logic;
          N_48_i_0                                                    : out   std_logic;
          N_46_i_0                                                    : out   std_logic;
          N_44_i_0                                                    : out   std_logic;
          N_42_i_0                                                    : out   std_logic;
          N_40_i_0                                                    : out   std_logic;
          N_38_i_0                                                    : out   std_logic;
          HTRANS_i_a2_0_0                                             : out   std_logic;
          N_271                                                       : in    std_logic;
          N_157_i_i_o2_0                                              : out   std_logic;
          N_157_i_i_o2_0_out                                          : out   std_logic;
          hsel2_i_4                                                   : out   std_logic;
          N_196_i_0                                                   : out   std_logic;
          N_195_i_0                                                   : out   std_logic;
          N_194_i_0                                                   : out   std_logic;
          N_65_i_0                                                    : out   std_logic;
          N_67_i_0                                                    : out   std_logic;
          N_110_i_0                                                   : out   std_logic;
          N_112_i_0                                                   : out   std_logic;
          N_114_i_0                                                   : out   std_logic;
          N_116_i_0                                                   : out   std_logic;
          N_69_i_0                                                    : out   std_logic;
          N_71_i_0                                                    : out   std_logic;
          N_73_i_0                                                    : out   std_logic;
          N_75_i_0                                                    : out   std_logic;
          N_77_i_0                                                    : out   std_logic;
          N_83_i_0                                                    : out   std_logic;
          N_85_i_0                                                    : out   std_logic;
          N_133_i_0                                                   : out   std_logic;
          N_87_i_0                                                    : out   std_logic;
          N_89_i_0                                                    : out   std_logic;
          N_140_i_0                                                   : out   std_logic;
          N_91_i_0                                                    : out   std_logic;
          N_93_i_0                                                    : out   std_logic;
          N_95_i_0                                                    : out   std_logic;
          N_97_i_0                                                    : out   std_logic;
          N_99_i_0                                                    : out   std_logic;
          N_152_i_0                                                   : out   std_logic;
          N_101_i_0                                                   : out   std_logic;
          N_156_i_0                                                   : out   std_logic;
          N_158_i_0                                                   : out   std_logic;
          N_103_i_0                                                   : out   std_logic;
          N_105_i_0                                                   : out   std_logic;
          N_107_i_0                                                   : out   std_logic;
          N_168_i_0                                                   : out   std_logic;
          N_109_i_0                                                   : out   std_logic;
          N_111_i_0                                                   : out   std_logic;
          N_218_i_0                                                   : out   std_logic;
          N_217_i_0                                                   : out   std_logic;
          N_203_i_0                                                   : out   std_logic
        );

end CoreAHBLite;

architecture DEF_ARCH of CoreAHBLite is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MATRIX4X16
    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE     : in    std_logic_vector(1 downto 0) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS    : in    std_logic_vector(1 to 1) := (others => 'U');
          result_addr_net_0                                           : in    std_logic_vector(3 downto 0) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP     : out   std_logic_vector(0 to 0);
          CoreAHBLite_0_AHBmslave3_HRDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          line_7                                                      : in    std_logic_vector(2 downto 1) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA    : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HADDR                              : out   std_logic_vector(11 to 11);
          xhdl1222_0                                                  : out   std_logic;
          xhdl1222_2                                                  : out   std_logic;
          SDATASELInt_0                                               : out   std_logic;
          SDATASELInt_1                                               : out   std_logic;
          SDATASELInt_2                                               : out   std_logic;
          SDATASELInt_4                                               : out   std_logic;
          SDATASELInt_6                                               : out   std_logic;
          SDATASELInt_7                                               : out   std_logic;
          SDATASELInt_8                                               : out   std_logic;
          SDATASELInt_9                                               : out   std_logic;
          SDATASELInt_10                                              : out   std_logic;
          SDATASELInt_11                                              : out   std_logic;
          SDATASELInt_12                                              : out   std_logic;
          SDATASELInt_13                                              : out   std_logic;
          arbRegSMCurrentState_13                                     : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31  : in    std_logic := 'U';
          line_13                                                     : in    std_logic := 'U';
          line_10                                                     : in    std_logic := 'U';
          line_21                                                     : in    std_logic := 'U';
          line_24                                                     : in    std_logic := 'U';
          line_18                                                     : in    std_logic := 'U';
          line_23                                                     : in    std_logic := 'U';
          line_16                                                     : in    std_logic := 'U';
          line_28                                                     : in    std_logic := 'U';
          line_9                                                      : in    std_logic := 'U';
          line_3_d0                                                   : in    std_logic := 'U';
          line_5_d0                                                   : in    std_logic := 'U';
          line_15                                                     : in    std_logic := 'U';
          line_26                                                     : in    std_logic := 'U';
          line_14                                                     : in    std_logic := 'U';
          line_20                                                     : in    std_logic := 'U';
          line_2_d0                                                   : in    std_logic := 'U';
          line_25                                                     : in    std_logic := 'U';
          line_29                                                     : in    std_logic := 'U';
          line_19                                                     : in    std_logic := 'U';
          line_27                                                     : in    std_logic := 'U';
          line_30                                                     : in    std_logic := 'U';
          line_17                                                     : in    std_logic := 'U';
          line_8                                                      : in    std_logic := 'U';
          line_0_d0                                                   : in    std_logic := 'U';
          line_6_d0                                                   : in    std_logic := 'U';
          line_1_d0                                                   : in    std_logic := 'U';
          line_0_10                                                   : in    std_logic := 'U';
          line_0_21                                                   : in    std_logic := 'U';
          line_0_24                                                   : in    std_logic := 'U';
          line_0_18                                                   : in    std_logic := 'U';
          line_0_23                                                   : in    std_logic := 'U';
          line_0_16                                                   : in    std_logic := 'U';
          line_0_28                                                   : in    std_logic := 'U';
          line_0_9                                                    : in    std_logic := 'U';
          line_0_3                                                    : in    std_logic := 'U';
          line_0_5                                                    : in    std_logic := 'U';
          line_0_15                                                   : in    std_logic := 'U';
          line_0_26                                                   : in    std_logic := 'U';
          line_0_14                                                   : in    std_logic := 'U';
          line_0_20                                                   : in    std_logic := 'U';
          line_0_2                                                    : in    std_logic := 'U';
          line_0_25                                                   : in    std_logic := 'U';
          line_0_29                                                   : in    std_logic := 'U';
          line_0_19                                                   : in    std_logic := 'U';
          line_0_27                                                   : in    std_logic := 'U';
          line_0_30                                                   : in    std_logic := 'U';
          line_0_17                                                   : in    std_logic := 'U';
          line_0_8                                                    : in    std_logic := 'U';
          line_0_0                                                    : in    std_logic := 'U';
          line_0_1                                                    : in    std_logic := 'U';
          line_0_6                                                    : in    std_logic := 'U';
          line_0_13                                                   : in    std_logic := 'U';
          line_1_10                                                   : in    std_logic := 'U';
          line_1_21                                                   : in    std_logic := 'U';
          line_1_24                                                   : in    std_logic := 'U';
          line_1_18                                                   : in    std_logic := 'U';
          line_1_23                                                   : in    std_logic := 'U';
          line_1_16                                                   : in    std_logic := 'U';
          line_1_28                                                   : in    std_logic := 'U';
          line_1_9                                                    : in    std_logic := 'U';
          line_1_3                                                    : in    std_logic := 'U';
          line_1_5                                                    : in    std_logic := 'U';
          line_1_15                                                   : in    std_logic := 'U';
          line_1_26                                                   : in    std_logic := 'U';
          line_1_14                                                   : in    std_logic := 'U';
          line_1_20                                                   : in    std_logic := 'U';
          line_1_2                                                    : in    std_logic := 'U';
          line_1_25                                                   : in    std_logic := 'U';
          line_1_29                                                   : in    std_logic := 'U';
          line_1_19                                                   : in    std_logic := 'U';
          line_1_27                                                   : in    std_logic := 'U';
          line_1_30                                                   : in    std_logic := 'U';
          line_1_17                                                   : in    std_logic := 'U';
          line_1_8                                                    : in    std_logic := 'U';
          line_1_0                                                    : in    std_logic := 'U';
          line_1_1                                                    : in    std_logic := 'U';
          line_1_6                                                    : in    std_logic := 'U';
          line_1_13                                                   : in    std_logic := 'U';
          line_2_19                                                   : in    std_logic := 'U';
          line_2_27                                                   : in    std_logic := 'U';
          line_2_30                                                   : in    std_logic := 'U';
          line_2_17                                                   : in    std_logic := 'U';
          line_2_8                                                    : in    std_logic := 'U';
          line_2_10                                                   : in    std_logic := 'U';
          line_2_15                                                   : in    std_logic := 'U';
          line_2_26                                                   : in    std_logic := 'U';
          line_2_20                                                   : in    std_logic := 'U';
          line_2_0                                                    : in    std_logic := 'U';
          line_2_1                                                    : in    std_logic := 'U';
          line_2_29                                                   : in    std_logic := 'U';
          line_2_25                                                   : in    std_logic := 'U';
          line_2_2                                                    : in    std_logic := 'U';
          line_2_6                                                    : in    std_logic := 'U';
          line_2_13                                                   : in    std_logic := 'U';
          line_2_14                                                   : in    std_logic := 'U';
          line_2_5                                                    : in    std_logic := 'U';
          line_2_3                                                    : in    std_logic := 'U';
          line_2_9                                                    : in    std_logic := 'U';
          line_2_28                                                   : in    std_logic := 'U';
          line_2_16                                                   : in    std_logic := 'U';
          line_2_23                                                   : in    std_logic := 'U';
          line_2_18                                                   : in    std_logic := 'U';
          line_2_24                                                   : in    std_logic := 'U';
          line_2_21                                                   : in    std_logic := 'U';
          line_3_19                                                   : in    std_logic := 'U';
          line_3_17                                                   : in    std_logic := 'U';
          line_3_8                                                    : in    std_logic := 'U';
          line_3_0                                                    : in    std_logic := 'U';
          line_3_1                                                    : in    std_logic := 'U';
          line_3_29                                                   : in    std_logic := 'U';
          line_3_25                                                   : in    std_logic := 'U';
          line_3_2                                                    : in    std_logic := 'U';
          line_3_20                                                   : in    std_logic := 'U';
          line_3_6                                                    : in    std_logic := 'U';
          line_3_13                                                   : in    std_logic := 'U';
          line_3_14                                                   : in    std_logic := 'U';
          line_3_26                                                   : in    std_logic := 'U';
          line_3_15                                                   : in    std_logic := 'U';
          line_3_5                                                    : in    std_logic := 'U';
          line_3_3                                                    : in    std_logic := 'U';
          line_3_9                                                    : in    std_logic := 'U';
          line_3_28                                                   : in    std_logic := 'U';
          line_3_16                                                   : in    std_logic := 'U';
          line_3_23                                                   : in    std_logic := 'U';
          line_3_18                                                   : in    std_logic := 'U';
          line_3_24                                                   : in    std_logic := 'U';
          line_3_21                                                   : in    std_logic := 'U';
          line_3_10                                                   : in    std_logic := 'U';
          SHA256_Module_0_data_out_5                                  : in    std_logic := 'U';
          SHA256_Module_0_data_out_13                                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_12                                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_8                                  : in    std_logic := 'U';
          SHA256_Module_0_data_out_23                                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_0                                  : in    std_logic := 'U';
          line_4_19                                                   : in    std_logic := 'U';
          line_4_17                                                   : in    std_logic := 'U';
          line_4_8                                                    : in    std_logic := 'U';
          line_4_0                                                    : in    std_logic := 'U';
          line_4_1                                                    : in    std_logic := 'U';
          line_4_29                                                   : in    std_logic := 'U';
          line_4_25                                                   : in    std_logic := 'U';
          line_4_2                                                    : in    std_logic := 'U';
          line_4_20                                                   : in    std_logic := 'U';
          line_4_14                                                   : in    std_logic := 'U';
          line_4_26                                                   : in    std_logic := 'U';
          line_4_15                                                   : in    std_logic := 'U';
          line_4_5                                                    : in    std_logic := 'U';
          line_4_3                                                    : in    std_logic := 'U';
          line_4_9                                                    : in    std_logic := 'U';
          line_4_28                                                   : in    std_logic := 'U';
          line_4_16                                                   : in    std_logic := 'U';
          line_4_23                                                   : in    std_logic := 'U';
          line_4_18                                                   : in    std_logic := 'U';
          line_4_24                                                   : in    std_logic := 'U';
          line_4_21                                                   : in    std_logic := 'U';
          line_4_10                                                   : in    std_logic := 'U';
          line_4_6                                                    : in    std_logic := 'U';
          line_4_13                                                   : in    std_logic := 'U';
          line_5_19                                                   : in    std_logic := 'U';
          line_5_17                                                   : in    std_logic := 'U';
          line_5_8                                                    : in    std_logic := 'U';
          line_5_0                                                    : in    std_logic := 'U';
          line_5_1                                                    : in    std_logic := 'U';
          line_5_29                                                   : in    std_logic := 'U';
          line_5_25                                                   : in    std_logic := 'U';
          line_5_2                                                    : in    std_logic := 'U';
          line_5_20                                                   : in    std_logic := 'U';
          line_5_6                                                    : in    std_logic := 'U';
          line_5_13                                                   : in    std_logic := 'U';
          line_5_14                                                   : in    std_logic := 'U';
          line_5_26                                                   : in    std_logic := 'U';
          line_5_15                                                   : in    std_logic := 'U';
          line_5_5                                                    : in    std_logic := 'U';
          line_5_3                                                    : in    std_logic := 'U';
          line_5_9                                                    : in    std_logic := 'U';
          line_5_28                                                   : in    std_logic := 'U';
          line_5_16                                                   : in    std_logic := 'U';
          line_5_23                                                   : in    std_logic := 'U';
          line_5_18                                                   : in    std_logic := 'U';
          line_5_24                                                   : in    std_logic := 'U';
          line_5_21                                                   : in    std_logic := 'U';
          line_5_10                                                   : in    std_logic := 'U';
          line_6_19                                                   : in    std_logic := 'U';
          line_6_17                                                   : in    std_logic := 'U';
          line_6_8                                                    : in    std_logic := 'U';
          line_6_0                                                    : in    std_logic := 'U';
          line_6_1                                                    : in    std_logic := 'U';
          line_6_29                                                   : in    std_logic := 'U';
          line_6_25                                                   : in    std_logic := 'U';
          line_6_2                                                    : in    std_logic := 'U';
          line_6_20                                                   : in    std_logic := 'U';
          line_6_6                                                    : in    std_logic := 'U';
          line_6_13                                                   : in    std_logic := 'U';
          line_6_14                                                   : in    std_logic := 'U';
          line_6_26                                                   : in    std_logic := 'U';
          line_6_15                                                   : in    std_logic := 'U';
          line_6_5                                                    : in    std_logic := 'U';
          line_6_3                                                    : in    std_logic := 'U';
          line_6_9                                                    : in    std_logic := 'U';
          line_6_28                                                   : in    std_logic := 'U';
          line_6_16                                                   : in    std_logic := 'U';
          line_6_23                                                   : in    std_logic := 'U';
          line_6_18                                                   : in    std_logic := 'U';
          line_6_24                                                   : in    std_logic := 'U';
          line_6_21                                                   : in    std_logic := 'U';
          line_6_10                                                   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11 : out   std_logic;
          MSS_READY                                                   : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                        : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE    : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                         : in    std_logic := 'U';
          CertificationSystem_sb_0_AHBmslave5_HREADY                  : in    std_logic := 'U';
          hready_m_xhdl344_7                                          : out   std_logic;
          N_225                                                       : out   std_logic;
          N_276                                                       : out   std_logic;
          N_259                                                       : out   std_logic;
          N_243                                                       : out   std_logic;
          N_236                                                       : out   std_logic;
          N_235                                                       : out   std_logic;
          N_277                                                       : out   std_logic;
          N_255                                                       : out   std_logic;
          N_241                                                       : out   std_logic;
          N_242                                                       : out   std_logic;
          N_244                                                       : out   std_logic;
          N_246                                                       : out   std_logic;
          N_247                                                       : out   std_logic;
          N_256                                                       : out   std_logic;
          N_257                                                       : out   std_logic;
          N_258                                                       : out   std_logic;
          ren_pos                                                     : in    std_logic := 'U';
          hready_m_xhdl343_10                                         : out   std_logic;
          hready_m_xhdl343_11                                         : out   std_logic;
          N_120                                                       : out   std_logic;
          N_216                                                       : in    std_logic := 'U';
          N_215                                                       : in    std_logic := 'U';
          hready_m_xhdl345                                            : out   std_logic;
          N_335                                                       : in    std_logic := 'U';
          N_214                                                       : in    std_logic := 'U';
          N_305                                                       : in    std_logic := 'U';
          N_206                                                       : out   std_logic;
          N_508                                                       : in    std_logic := 'U';
          N_478_i_0                                                   : out   std_logic;
          N_507                                                       : in    std_logic := 'U';
          N_477_i_0                                                   : out   std_logic;
          N_479_i_0                                                   : out   std_logic;
          N_480_i_0                                                   : out   std_logic;
          N_481_i_0                                                   : out   std_logic;
          un8_hreadyin_i_0                                            : in    std_logic := 'U';
          N_9_i_0                                                     : out   std_logic;
          N_226                                                       : out   std_logic;
          defSlaveSMNextState                                         : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                     : in    std_logic := 'U';
          N_63_i_0                                                    : out   std_logic;
          N_62_i_0                                                    : out   std_logic;
          N_60_i_0                                                    : out   std_logic;
          N_98_i_0                                                    : out   std_logic;
          N_96_i_0                                                    : out   std_logic;
          N_94_i_0                                                    : out   std_logic;
          N_92_i_0                                                    : out   std_logic;
          N_90_i_0                                                    : out   std_logic;
          N_88_i_0                                                    : out   std_logic;
          N_86_i_0                                                    : out   std_logic;
          N_84_i_0                                                    : out   std_logic;
          N_82_i_0                                                    : out   std_logic;
          N_80_i_0                                                    : out   std_logic;
          N_78_i_0                                                    : out   std_logic;
          N_76_i_0                                                    : out   std_logic;
          N_74_i_0                                                    : out   std_logic;
          N_72_i_0                                                    : out   std_logic;
          N_70_i_0                                                    : out   std_logic;
          N_68_i_0                                                    : out   std_logic;
          N_66_i_0                                                    : out   std_logic;
          N_64_i_0                                                    : out   std_logic;
          N_58_i_0                                                    : out   std_logic;
          N_56_i_0                                                    : out   std_logic;
          N_54_i_0                                                    : out   std_logic;
          N_52_i_0                                                    : out   std_logic;
          N_50_i_0                                                    : out   std_logic;
          N_48_i_0                                                    : out   std_logic;
          N_46_i_0                                                    : out   std_logic;
          N_44_i_0                                                    : out   std_logic;
          N_42_i_0                                                    : out   std_logic;
          N_40_i_0                                                    : out   std_logic;
          N_38_i_0                                                    : out   std_logic;
          HTRANS_i_a2_0_0                                             : out   std_logic;
          N_271                                                       : in    std_logic := 'U';
          N_157_i_i_o2_0                                              : out   std_logic;
          N_157_i_i_o2_0_out                                          : out   std_logic;
          hsel2_i_4                                                   : out   std_logic;
          N_196_i_0                                                   : out   std_logic;
          N_195_i_0                                                   : out   std_logic;
          N_194_i_0                                                   : out   std_logic;
          N_65_i_0                                                    : out   std_logic;
          N_67_i_0                                                    : out   std_logic;
          N_110_i_0                                                   : out   std_logic;
          N_112_i_0                                                   : out   std_logic;
          N_114_i_0                                                   : out   std_logic;
          N_116_i_0                                                   : out   std_logic;
          N_69_i_0                                                    : out   std_logic;
          N_71_i_0                                                    : out   std_logic;
          N_73_i_0                                                    : out   std_logic;
          N_75_i_0                                                    : out   std_logic;
          N_77_i_0                                                    : out   std_logic;
          N_83_i_0                                                    : out   std_logic;
          N_85_i_0                                                    : out   std_logic;
          N_133_i_0                                                   : out   std_logic;
          N_87_i_0                                                    : out   std_logic;
          N_89_i_0                                                    : out   std_logic;
          N_140_i_0                                                   : out   std_logic;
          N_91_i_0                                                    : out   std_logic;
          N_93_i_0                                                    : out   std_logic;
          N_95_i_0                                                    : out   std_logic;
          N_97_i_0                                                    : out   std_logic;
          N_99_i_0                                                    : out   std_logic;
          N_152_i_0                                                   : out   std_logic;
          N_101_i_0                                                   : out   std_logic;
          N_156_i_0                                                   : out   std_logic;
          N_158_i_0                                                   : out   std_logic;
          N_103_i_0                                                   : out   std_logic;
          N_105_i_0                                                   : out   std_logic;
          N_107_i_0                                                   : out   std_logic;
          N_168_i_0                                                   : out   std_logic;
          N_109_i_0                                                   : out   std_logic;
          N_111_i_0                                                   : out   std_logic;
          N_218_i_0                                                   : out   std_logic;
          N_217_i_0                                                   : out   std_logic;
          N_203_i_0                                                   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : COREAHBLITE_MATRIX4X16
	Use entity work.COREAHBLITE_MATRIX4X16(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    matrix4x16 : COREAHBLITE_MATRIX4X16
      port map(
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        result_addr_net_0(3) => result_addr_net_0(3), 
        result_addr_net_0(2) => result_addr_net_0(2), 
        result_addr_net_0(1) => result_addr_net_0(1), 
        result_addr_net_0(0) => result_addr_net_0(0), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        CoreAHBLite_0_AHBmslave3_HRDATA(31) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(31), 
        CoreAHBLite_0_AHBmslave3_HRDATA(30) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(30), 
        CoreAHBLite_0_AHBmslave3_HRDATA(29) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(29), 
        CoreAHBLite_0_AHBmslave3_HRDATA(28) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(28), 
        CoreAHBLite_0_AHBmslave3_HRDATA(27) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(27), 
        CoreAHBLite_0_AHBmslave3_HRDATA(26) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(26), 
        CoreAHBLite_0_AHBmslave3_HRDATA(25) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(25), 
        CoreAHBLite_0_AHBmslave3_HRDATA(24) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(24), 
        CoreAHBLite_0_AHBmslave3_HRDATA(23) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(23), 
        CoreAHBLite_0_AHBmslave3_HRDATA(22) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(22), 
        CoreAHBLite_0_AHBmslave3_HRDATA(21) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(21), 
        CoreAHBLite_0_AHBmslave3_HRDATA(20) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(20), 
        CoreAHBLite_0_AHBmslave3_HRDATA(19) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(19), 
        CoreAHBLite_0_AHBmslave3_HRDATA(18) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(18), 
        CoreAHBLite_0_AHBmslave3_HRDATA(17) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(17), 
        CoreAHBLite_0_AHBmslave3_HRDATA(16) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(16), 
        CoreAHBLite_0_AHBmslave3_HRDATA(15) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(15), 
        CoreAHBLite_0_AHBmslave3_HRDATA(14) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(14), 
        CoreAHBLite_0_AHBmslave3_HRDATA(13) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(13), 
        CoreAHBLite_0_AHBmslave3_HRDATA(12) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(12), 
        CoreAHBLite_0_AHBmslave3_HRDATA(11) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(11), 
        CoreAHBLite_0_AHBmslave3_HRDATA(10) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(10), 
        CoreAHBLite_0_AHBmslave3_HRDATA(9) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(9), 
        CoreAHBLite_0_AHBmslave3_HRDATA(8) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(8), 
        CoreAHBLite_0_AHBmslave3_HRDATA(7) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(7), 
        CoreAHBLite_0_AHBmslave3_HRDATA(6) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(6), 
        CoreAHBLite_0_AHBmslave3_HRDATA(5) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(5), 
        CoreAHBLite_0_AHBmslave3_HRDATA(4) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(4), 
        CoreAHBLite_0_AHBmslave3_HRDATA(3) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(3), 
        CoreAHBLite_0_AHBmslave3_HRDATA(2) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(2), 
        CoreAHBLite_0_AHBmslave3_HRDATA(1) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(1), 
        CoreAHBLite_0_AHBmslave3_HRDATA(0) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(0), line_7(2) => 
        line_7(2), line_7(1) => line_7(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        CoreAHBLite_0_AHBmslave3_HADDR(11) => 
        CoreAHBLite_0_AHBmslave3_HADDR(11), xhdl1222_0 => 
        xhdl1222_0, xhdl1222_2 => xhdl1222_2, SDATASELInt_0 => 
        SDATASELInt_0, SDATASELInt_1 => SDATASELInt_1, 
        SDATASELInt_2 => SDATASELInt_2, SDATASELInt_4 => 
        SDATASELInt_4, SDATASELInt_6 => SDATASELInt_6, 
        SDATASELInt_7 => SDATASELInt_7, SDATASELInt_8 => 
        SDATASELInt_8, SDATASELInt_9 => SDATASELInt_9, 
        SDATASELInt_10 => SDATASELInt_10, SDATASELInt_11 => 
        SDATASELInt_11, SDATASELInt_12 => SDATASELInt_12, 
        SDATASELInt_13 => SDATASELInt_13, arbRegSMCurrentState_13
         => arbRegSMCurrentState(15), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        line_13 => line_13, line_10 => line_10, line_21 => 
        line_21, line_24 => line_24, line_18 => line_18, line_23
         => line_23, line_16 => line_16, line_28 => line_28, 
        line_9 => line_9, line_3_d0 => line_3_d0, line_5_d0 => 
        line_5_d0, line_15 => line_15, line_26 => line_26, 
        line_14 => line_14, line_20 => line_20, line_2_d0 => 
        line_2_d0, line_25 => line_25, line_29 => line_29, 
        line_19 => line_19, line_27 => line_27, line_30 => 
        line_30, line_17 => line_17, line_8 => line_8, line_0_d0
         => line_0_d0, line_6_d0 => line_6_d0, line_1_d0 => 
        line_1_d0, line_0_10 => line_0_10, line_0_21 => line_0_21, 
        line_0_24 => line_0_24, line_0_18 => line_0_18, line_0_23
         => line_0_23, line_0_16 => line_0_16, line_0_28 => 
        line_0_28, line_0_9 => line_0_9, line_0_3 => line_0_3, 
        line_0_5 => line_0_5, line_0_15 => line_0_15, line_0_26
         => line_0_26, line_0_14 => line_0_14, line_0_20 => 
        line_0_20, line_0_2 => line_0_2, line_0_25 => line_0_25, 
        line_0_29 => line_0_29, line_0_19 => line_0_19, line_0_27
         => line_0_27, line_0_30 => line_0_30, line_0_17 => 
        line_0_17, line_0_8 => line_0_8, line_0_0 => line_0_0, 
        line_0_1 => line_0_1, line_0_6 => line_0_6, line_0_13 => 
        line_0_13, line_1_10 => line_1_10, line_1_21 => line_1_21, 
        line_1_24 => line_1_24, line_1_18 => line_1_18, line_1_23
         => line_1_23, line_1_16 => line_1_16, line_1_28 => 
        line_1_28, line_1_9 => line_1_9, line_1_3 => line_1_3, 
        line_1_5 => line_1_5, line_1_15 => line_1_15, line_1_26
         => line_1_26, line_1_14 => line_1_14, line_1_20 => 
        line_1_20, line_1_2 => line_1_2, line_1_25 => line_1_25, 
        line_1_29 => line_1_29, line_1_19 => line_1_19, line_1_27
         => line_1_27, line_1_30 => line_1_30, line_1_17 => 
        line_1_17, line_1_8 => line_1_8, line_1_0 => line_1_0, 
        line_1_1 => line_1_1, line_1_6 => line_1_6, line_1_13 => 
        line_1_13, line_2_19 => line_2_19, line_2_27 => line_2_27, 
        line_2_30 => line_2_30, line_2_17 => line_2_17, line_2_8
         => line_2_8, line_2_10 => line_2_10, line_2_15 => 
        line_2_15, line_2_26 => line_2_26, line_2_20 => line_2_20, 
        line_2_0 => line_2_0, line_2_1 => line_2_1, line_2_29 => 
        line_2_29, line_2_25 => line_2_25, line_2_2 => line_2_2, 
        line_2_6 => line_2_6, line_2_13 => line_2_13, line_2_14
         => line_2_14, line_2_5 => line_2_5, line_2_3 => line_2_3, 
        line_2_9 => line_2_9, line_2_28 => line_2_28, line_2_16
         => line_2_16, line_2_23 => line_2_23, line_2_18 => 
        line_2_18, line_2_24 => line_2_24, line_2_21 => line_2_21, 
        line_3_19 => line_3_19, line_3_17 => line_3_17, line_3_8
         => line_3_8, line_3_0 => line_3_0, line_3_1 => line_3_1, 
        line_3_29 => line_3_29, line_3_25 => line_3_25, line_3_2
         => line_3_2, line_3_20 => line_3_20, line_3_6 => 
        line_3_6, line_3_13 => line_3_13, line_3_14 => line_3_14, 
        line_3_26 => line_3_26, line_3_15 => line_3_15, line_3_5
         => line_3_5, line_3_3 => line_3_3, line_3_9 => line_3_9, 
        line_3_28 => line_3_28, line_3_16 => line_3_16, line_3_23
         => line_3_23, line_3_18 => line_3_18, line_3_24 => 
        line_3_24, line_3_21 => line_3_21, line_3_10 => line_3_10, 
        SHA256_Module_0_data_out_5 => SHA256_Module_0_data_out_5, 
        SHA256_Module_0_data_out_13 => 
        SHA256_Module_0_data_out_13, SHA256_Module_0_data_out_12
         => SHA256_Module_0_data_out_12, 
        SHA256_Module_0_data_out_8 => SHA256_Module_0_data_out_8, 
        SHA256_Module_0_data_out_23 => 
        SHA256_Module_0_data_out_23, SHA256_Module_0_data_out_0
         => SHA256_Module_0_data_out_0, line_4_19 => line_4_19, 
        line_4_17 => line_4_17, line_4_8 => line_4_8, line_4_0
         => line_4_0, line_4_1 => line_4_1, line_4_29 => 
        line_4_29, line_4_25 => line_4_25, line_4_2 => line_4_2, 
        line_4_20 => line_4_20, line_4_14 => line_4_14, line_4_26
         => line_4_26, line_4_15 => line_4_15, line_4_5 => 
        line_4_5, line_4_3 => line_4_3, line_4_9 => line_4_9, 
        line_4_28 => line_4_28, line_4_16 => line_4_16, line_4_23
         => line_4_23, line_4_18 => line_4_18, line_4_24 => 
        line_4_24, line_4_21 => line_4_21, line_4_10 => line_4_10, 
        line_4_6 => line_4_6, line_4_13 => line_4_13, line_5_19
         => line_5_19, line_5_17 => line_5_17, line_5_8 => 
        line_5_8, line_5_0 => line_5_0, line_5_1 => line_5_1, 
        line_5_29 => line_5_29, line_5_25 => line_5_25, line_5_2
         => line_5_2, line_5_20 => line_5_20, line_5_6 => 
        line_5_6, line_5_13 => line_5_13, line_5_14 => line_5_14, 
        line_5_26 => line_5_26, line_5_15 => line_5_15, line_5_5
         => line_5_5, line_5_3 => line_5_3, line_5_9 => line_5_9, 
        line_5_28 => line_5_28, line_5_16 => line_5_16, line_5_23
         => line_5_23, line_5_18 => line_5_18, line_5_24 => 
        line_5_24, line_5_21 => line_5_21, line_5_10 => line_5_10, 
        line_6_19 => line_6_19, line_6_17 => line_6_17, line_6_8
         => line_6_8, line_6_0 => line_6_0, line_6_1 => line_6_1, 
        line_6_29 => line_6_29, line_6_25 => line_6_25, line_6_2
         => line_6_2, line_6_20 => line_6_20, line_6_6 => 
        line_6_6, line_6_13 => line_6_13, line_6_14 => line_6_14, 
        line_6_26 => line_6_26, line_6_15 => line_6_15, line_6_5
         => line_6_5, line_6_3 => line_6_3, line_6_9 => line_6_9, 
        line_6_28 => line_6_28, line_6_16 => line_6_16, line_6_23
         => line_6_23, line_6_18 => line_6_18, line_6_24 => 
        line_6_24, line_6_21 => line_6_21, line_6_10 => line_6_10, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11, 
        MSS_READY => MSS_READY, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, 
        CertificationSystem_sb_0_AHBmslave5_HREADY => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, 
        hready_m_xhdl344_7 => hready_m_xhdl344_7, N_225 => N_225, 
        N_276 => N_276, N_259 => N_259, N_243 => N_243, N_236 => 
        N_236, N_235 => N_235, N_277 => N_277, N_255 => N_255, 
        N_241 => N_241, N_242 => N_242, N_244 => N_244, N_246 => 
        N_246, N_247 => N_247, N_256 => N_256, N_257 => N_257, 
        N_258 => N_258, ren_pos => ren_pos, hready_m_xhdl343_10
         => hready_m_xhdl343_10, hready_m_xhdl343_11 => 
        hready_m_xhdl343_11, N_120 => N_120, N_216 => N_216, 
        N_215 => N_215, hready_m_xhdl345 => hready_m_xhdl345, 
        N_335 => N_335, N_214 => N_214, N_305 => N_305, N_206 => 
        N_206, N_508 => N_508, N_478_i_0 => N_478_i_0, N_507 => 
        N_507, N_477_i_0 => N_477_i_0, N_479_i_0 => N_479_i_0, 
        N_480_i_0 => N_480_i_0, N_481_i_0 => N_481_i_0, 
        un8_hreadyin_i_0 => un8_hreadyin_i_0, N_9_i_0 => N_9_i_0, 
        N_226 => N_226, defSlaveSMNextState => 
        defSlaveSMNextState, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, N_63_i_0 => 
        N_63_i_0, N_62_i_0 => N_62_i_0, N_60_i_0 => N_60_i_0, 
        N_98_i_0 => N_98_i_0, N_96_i_0 => N_96_i_0, N_94_i_0 => 
        N_94_i_0, N_92_i_0 => N_92_i_0, N_90_i_0 => N_90_i_0, 
        N_88_i_0 => N_88_i_0, N_86_i_0 => N_86_i_0, N_84_i_0 => 
        N_84_i_0, N_82_i_0 => N_82_i_0, N_80_i_0 => N_80_i_0, 
        N_78_i_0 => N_78_i_0, N_76_i_0 => N_76_i_0, N_74_i_0 => 
        N_74_i_0, N_72_i_0 => N_72_i_0, N_70_i_0 => N_70_i_0, 
        N_68_i_0 => N_68_i_0, N_66_i_0 => N_66_i_0, N_64_i_0 => 
        N_64_i_0, N_58_i_0 => N_58_i_0, N_56_i_0 => N_56_i_0, 
        N_54_i_0 => N_54_i_0, N_52_i_0 => N_52_i_0, N_50_i_0 => 
        N_50_i_0, N_48_i_0 => N_48_i_0, N_46_i_0 => N_46_i_0, 
        N_44_i_0 => N_44_i_0, N_42_i_0 => N_42_i_0, N_40_i_0 => 
        N_40_i_0, N_38_i_0 => N_38_i_0, HTRANS_i_a2_0_0 => 
        HTRANS_i_a2_0_0, N_271 => N_271, N_157_i_i_o2_0 => 
        N_157_i_i_o2_0, N_157_i_i_o2_0_out => N_157_i_i_o2_0_out, 
        hsel2_i_4 => hsel2_i_4, N_196_i_0 => N_196_i_0, N_195_i_0
         => N_195_i_0, N_194_i_0 => N_194_i_0, N_65_i_0 => 
        N_65_i_0, N_67_i_0 => N_67_i_0, N_110_i_0 => N_110_i_0, 
        N_112_i_0 => N_112_i_0, N_114_i_0 => N_114_i_0, N_116_i_0
         => N_116_i_0, N_69_i_0 => N_69_i_0, N_71_i_0 => N_71_i_0, 
        N_73_i_0 => N_73_i_0, N_75_i_0 => N_75_i_0, N_77_i_0 => 
        N_77_i_0, N_83_i_0 => N_83_i_0, N_85_i_0 => N_85_i_0, 
        N_133_i_0 => N_133_i_0, N_87_i_0 => N_87_i_0, N_89_i_0
         => N_89_i_0, N_140_i_0 => N_140_i_0, N_91_i_0 => 
        N_91_i_0, N_93_i_0 => N_93_i_0, N_95_i_0 => N_95_i_0, 
        N_97_i_0 => N_97_i_0, N_99_i_0 => N_99_i_0, N_152_i_0 => 
        N_152_i_0, N_101_i_0 => N_101_i_0, N_156_i_0 => N_156_i_0, 
        N_158_i_0 => N_158_i_0, N_103_i_0 => N_103_i_0, N_105_i_0
         => N_105_i_0, N_107_i_0 => N_107_i_0, N_168_i_0 => 
        N_168_i_0, N_109_i_0 => N_109_i_0, N_111_i_0 => N_111_i_0, 
        N_218_i_0 => N_218_i_0, N_217_i_0 => N_217_i_0, N_203_i_0
         => N_203_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_MSS is

    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE     : out   std_logic_vector(1 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS    : out   std_logic_vector(1 to 1);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA    : out   std_logic_vector(31 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP     : in    std_logic_vector(0 to 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8  : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29 : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30 : in    std_logic;
          SPI_0_SS0                                                   : inout std_logic := 'Z';
          SPI_0_DO                                                    : out   std_logic;
          SPI_0_DI                                                    : in    std_logic;
          SPI_0_CLK                                                   : inout std_logic := 'Z';
          MMUART_1_TXD                                                : out   std_logic;
          MMUART_1_RXD                                                : in    std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N       : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE    : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F            : out   std_logic;
          CertificationSystem_sb_0_GPIO_1_M2F                         : out   std_logic;
          GPIO_0_M2F_c                                                : out   std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F                         : out   std_logic;
          N_481_i_0                                                   : in    std_logic;
          N_480_i_0                                                   : in    std_logic;
          N_479_i_0                                                   : in    std_logic;
          N_478_i_0                                                   : in    std_logic;
          N_477_i_0                                                   : in    std_logic;
          N_9_i_0                                                     : in    std_logic;
          FAB_CCC_LOCK                                                : in    std_logic;
          SHA256_Module_0_waiting_data                                : in    std_logic;
          SHA256_Module_0_data_available_lastbank_8                   : in    std_logic;
          SHA256_Module_0_di_req_o                                    : in    std_logic;
          SHA256_Module_0_do_valid_o                                  : in    std_logic;
          SHA256_Module_0_data_available                              : in    std_logic;
          SHA256_Module_0_error_o                                     : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                        : in    std_logic
        );

end CertificationSystem_sb_MSS;

architecture DEF_ARCH of CertificationSystem_sb_MSS is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component TRIBUFF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component MSS_075

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MGPIO0B_IN                              : in    std_logic := 'U';
          MGPIO10B_IN                             : in    std_logic := 'U';
          MGPIO1B_IN                              : in    std_logic := 'U';
          MGPIO25A_IN                             : in    std_logic := 'U';
          MGPIO26A_IN                             : in    std_logic := 'U';
          MGPIO27A_IN                             : in    std_logic := 'U';
          MGPIO28A_IN                             : in    std_logic := 'U';
          MGPIO29A_IN                             : in    std_logic := 'U';
          MGPIO2B_IN                              : in    std_logic := 'U';
          MGPIO30A_IN                             : in    std_logic := 'U';
          MGPIO31A_IN                             : in    std_logic := 'U';
          MGPIO3B_IN                              : in    std_logic := 'U';
          MGPIO4B_IN                              : in    std_logic := 'U';
          MGPIO5B_IN                              : in    std_logic := 'U';
          MGPIO6B_IN                              : in    std_logic := 'U';
          MGPIO7B_IN                              : in    std_logic := 'U';
          MGPIO8B_IN                              : in    std_logic := 'U';
          MGPIO9B_IN                              : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_CTS_MGPIO13B_IN                 : in    std_logic := 'U';
          MMUART1_DCD_MGPIO16B_IN                 : in    std_logic := 'U';
          MMUART1_DSR_MGPIO14B_IN                 : in    std_logic := 'U';
          MMUART1_DTR_MGPIO12B_IN                 : in    std_logic := 'U';
          MMUART1_RI_MGPIO15B_IN                  : in    std_logic := 'U';
          MMUART1_RTS_MGPIO11B_IN                 : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI0_SS4_MGPIO19A_IN                    : in    std_logic := 'U';
          SPI0_SS5_MGPIO20A_IN                    : in    std_logic := 'U';
          SPI0_SS6_MGPIO21A_IN                    : in    std_logic := 'U';
          SPI0_SS7_MGPIO22A_IN                    : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          USBD_DATA0_IN                           : in    std_logic := 'U';
          USBD_DATA1_IN                           : in    std_logic := 'U';
          USBD_DATA2_IN                           : in    std_logic := 'U';
          USBD_DATA3_IN                           : in    std_logic := 'U';
          USBD_DATA4_IN                           : in    std_logic := 'U';
          USBD_DATA5_IN                           : in    std_logic := 'U';
          USBD_DATA6_IN                           : in    std_logic := 'U';
          USBD_DATA7_MGPIO23B_IN                  : in    std_logic := 'U';
          USBD_DIR_IN                             : in    std_logic := 'U';
          USBD_NXT_IN                             : in    std_logic := 'U';
          USBD_STP_IN                             : in    std_logic := 'U';
          USBD_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MGPIO0B_OUT                             : out   std_logic;
          MGPIO10B_OUT                            : out   std_logic;
          MGPIO1B_OUT                             : out   std_logic;
          MGPIO25A_OUT                            : out   std_logic;
          MGPIO26A_OUT                            : out   std_logic;
          MGPIO27A_OUT                            : out   std_logic;
          MGPIO28A_OUT                            : out   std_logic;
          MGPIO29A_OUT                            : out   std_logic;
          MGPIO2B_OUT                             : out   std_logic;
          MGPIO30A_OUT                            : out   std_logic;
          MGPIO31A_OUT                            : out   std_logic;
          MGPIO3B_OUT                             : out   std_logic;
          MGPIO4B_OUT                             : out   std_logic;
          MGPIO5B_OUT                             : out   std_logic;
          MGPIO6B_OUT                             : out   std_logic;
          MGPIO7B_OUT                             : out   std_logic;
          MGPIO8B_OUT                             : out   std_logic;
          MGPIO9B_OUT                             : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_CTS_MGPIO13B_OUT                : out   std_logic;
          MMUART1_DCD_MGPIO16B_OUT                : out   std_logic;
          MMUART1_DSR_MGPIO14B_OUT                : out   std_logic;
          MMUART1_DTR_MGPIO12B_OUT                : out   std_logic;
          MMUART1_RI_MGPIO15B_OUT                 : out   std_logic;
          MMUART1_RTS_MGPIO11B_OUT                : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI0_SS4_MGPIO19A_OUT                   : out   std_logic;
          SPI0_SS5_MGPIO20A_OUT                   : out   std_logic;
          SPI0_SS6_MGPIO21A_OUT                   : out   std_logic;
          SPI0_SS7_MGPIO22A_OUT                   : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          USBD_DATA0_OUT                          : out   std_logic;
          USBD_DATA1_OUT                          : out   std_logic;
          USBD_DATA2_OUT                          : out   std_logic;
          USBD_DATA3_OUT                          : out   std_logic;
          USBD_DATA4_OUT                          : out   std_logic;
          USBD_DATA5_OUT                          : out   std_logic;
          USBD_DATA6_OUT                          : out   std_logic;
          USBD_DATA7_MGPIO23B_OUT                 : out   std_logic;
          USBD_DIR_OUT                            : out   std_logic;
          USBD_NXT_OUT                            : out   std_logic;
          USBD_STP_OUT                            : out   std_logic;
          USBD_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MGPIO0B_OE                              : out   std_logic;
          MGPIO10B_OE                             : out   std_logic;
          MGPIO1B_OE                              : out   std_logic;
          MGPIO25A_OE                             : out   std_logic;
          MGPIO26A_OE                             : out   std_logic;
          MGPIO27A_OE                             : out   std_logic;
          MGPIO28A_OE                             : out   std_logic;
          MGPIO29A_OE                             : out   std_logic;
          MGPIO2B_OE                              : out   std_logic;
          MGPIO30A_OE                             : out   std_logic;
          MGPIO31A_OE                             : out   std_logic;
          MGPIO3B_OE                              : out   std_logic;
          MGPIO4B_OE                              : out   std_logic;
          MGPIO5B_OE                              : out   std_logic;
          MGPIO6B_OE                              : out   std_logic;
          MGPIO7B_OE                              : out   std_logic;
          MGPIO8B_OE                              : out   std_logic;
          MGPIO9B_OE                              : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_CTS_MGPIO13B_OE                 : out   std_logic;
          MMUART1_DCD_MGPIO16B_OE                 : out   std_logic;
          MMUART1_DSR_MGPIO14B_OE                 : out   std_logic;
          MMUART1_DTR_MGPIO12B_OE                 : out   std_logic;
          MMUART1_RI_MGPIO15B_OE                  : out   std_logic;
          MMUART1_RTS_MGPIO11B_OE                 : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI0_SS4_MGPIO19A_OE                    : out   std_logic;
          SPI0_SS5_MGPIO20A_OE                    : out   std_logic;
          SPI0_SS6_MGPIO21A_OE                    : out   std_logic;
          SPI0_SS7_MGPIO22A_OE                    : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic;
          USBD_DATA0_OE                           : out   std_logic;
          USBD_DATA1_OE                           : out   std_logic;
          USBD_DATA2_OE                           : out   std_logic;
          USBD_DATA3_OE                           : out   std_logic;
          USBD_DATA4_OE                           : out   std_logic;
          USBD_DATA5_OE                           : out   std_logic;
          USBD_DATA6_OE                           : out   std_logic;
          USBD_DATA7_MGPIO23B_OE                  : out   std_logic;
          USBD_DIR_OE                             : out   std_logic;
          USBD_NXT_OE                             : out   std_logic;
          USBD_STP_OE                             : out   std_logic;
          USBD_XCLK_OE                            : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal SPI_0_SS0_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI_0_DI_PAD_Y, SPI_0_CLK_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        MMUART_1_RXD_PAD_Y, VCC_net_1, GND_net_1 : std_logic;
    signal nc228, nc203, nc265, nc216, nc194, nc151, nc23, nc175, 
        nc250, nc58, nc116, nc74, nc133, nc238, nc167, nc84, nc39, 
        nc72, nc256, nc212, nc205, nc82, nc145, nc181, nc160, 
        nc57, nc156, nc280, nc125, nc211, nc73, nc107, nc66, nc83, 
        nc9, nc252, nc171, nc54, nc286, nc307, nc135, nc41, nc100, 
        nc270, nc52, nc251, nc186, nc29, nc269, nc118, nc60, 
        nc141, nc311, nc276, nc193, nc214, nc298, nc282, nc240, 
        nc45, nc53, nc121, nc176, nc220, nc158, nc281, nc209, 
        nc246, nc162, nc11, nc272, nc131, nc254, nc267, nc96, 
        nc79, nc226, nc146, nc230, nc89, nc119, nc48, nc271, 
        nc213, nc300, nc126, nc195, nc188, nc242, nc15, nc308, 
        nc236, nc102, nc304, nc3, nc207, nc47, nc90, nc284, nc222, 
        nc159, nc136, nc241, nc253, nc178, nc306, nc215, nc59, 
        nc221, nc232, nc274, nc18, nc44, nc117, nc189, nc164, 
        nc148, nc42, nc231, nc191, nc255, nc283, nc317, nc290, 
        nc17, nc2, nc302, nc110, nc128, nc244, nc321, nc43, nc179, 
        nc157, nc36, nc224, nc296, nc273, nc61, nc104, nc138, 
        nc14, nc285, nc303, nc150, nc196, nc234, nc149, nc12, 
        nc219, nc30, nc243, nc187, nc65, nc7, nc292, nc129, nc275, 
        nc8, nc223, nc13, nc305, nc180, nc26, nc291, nc177, nc139, 
        nc310, nc259, nc245, nc233, nc163, nc318, nc268, nc112, 
        nc68, nc49, nc314, nc217, nc170, nc91, nc225, nc5, nc20, 
        nc198, nc147, nc316, nc67, nc289, nc294, nc152, nc127, 
        nc103, nc235, nc76, nc208, nc140, nc257, nc86, nc95, 
        nc120, nc165, nc279, nc137, nc64, nc19, nc312, nc70, 
        nc182, nc62, nc199, nc80, nc130, nc287, nc98, nc293, 
        nc249, nc114, nc56, nc105, nc63, nc313, nc309, nc172, 
        nc229, nc277, nc97, nc161, nc31, nc295, nc154, nc50, 
        nc260, nc239, nc142, nc320, nc315, nc247, nc94, nc197, 
        nc122, nc266, nc35, nc4, nc227, nc92, nc101, nc184, nc200, 
        nc190, nc166, nc132, nc21, nc237, nc93, nc262, nc69, 
        nc206, nc174, nc38, nc113, nc218, nc106, nc261, nc25, nc1, 
        nc299, nc37, nc202, nc144, nc153, nc46, nc258, nc71, 
        nc124, nc81, nc201, nc168, nc34, nc28, nc115, nc264, 
        nc192, nc319, nc134, nc32, nc40, nc297, nc99, nc75, nc183, 
        nc288, nc85, nc27, nc108, nc16, nc155, nc51, nc301, nc33, 
        nc204, nc173, nc278, nc169, nc78, nc263, nc24, nc88, 
        nc111, nc55, nc10, nc22, nc210, nc185, nc143, nc248, nc77, 
        nc6, nc109, nc87, nc123 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    SPI_0_DO_PAD : TRIBUFF
      port map(D => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        E => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, PAD => 
        SPI_0_DO);
    
    SPI_0_SS0_PAD : BIBUF
      port map(PAD => SPI_0_SS0, D => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, Y => 
        SPI_0_SS0_PAD_Y);
    
    SPI_0_DI_PAD : INBUF
      port map(PAD => SPI_0_DI, Y => SPI_0_DI_PAD_Y);
    
    MSS_ADLIB_INST : MSS_075

              generic map(INIT => "00" & x"0000000000000000000000000000036100080000000000000000000000000000000000000000000000000000000000001203610000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C35C00000000609300000003FFFFE4000000000000100000000F0E15C00000182DF34010842108421000001FE34001FF8000000400000000000451007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem", RTC_MAIN_XTL_FREQ => 0.0,
         DDR_CLK_FREQ => 50.0)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => OPEN, CAN_TX_EBL_MGPIO4A_H2F_A
         => OPEN, CAN_TX_EBL_MGPIO4A_H2F_B => OPEN, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => OPEN, CLK_CONFIG_APB => OPEN, COMMS_INT => OPEN, 
        CONFIG_PRESET_N => 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        EDAC_ERROR(7) => nc228, EDAC_ERROR(6) => nc203, 
        EDAC_ERROR(5) => nc265, EDAC_ERROR(4) => nc216, 
        EDAC_ERROR(3) => nc194, EDAC_ERROR(2) => nc151, 
        EDAC_ERROR(1) => nc23, EDAC_ERROR(0) => nc175, 
        F_FM0_RDATA(31) => nc250, F_FM0_RDATA(30) => nc58, 
        F_FM0_RDATA(29) => nc116, F_FM0_RDATA(28) => nc74, 
        F_FM0_RDATA(27) => nc133, F_FM0_RDATA(26) => nc238, 
        F_FM0_RDATA(25) => nc167, F_FM0_RDATA(24) => nc84, 
        F_FM0_RDATA(23) => nc39, F_FM0_RDATA(22) => nc72, 
        F_FM0_RDATA(21) => nc256, F_FM0_RDATA(20) => nc212, 
        F_FM0_RDATA(19) => nc205, F_FM0_RDATA(18) => nc82, 
        F_FM0_RDATA(17) => nc145, F_FM0_RDATA(16) => nc181, 
        F_FM0_RDATA(15) => nc160, F_FM0_RDATA(14) => nc57, 
        F_FM0_RDATA(13) => nc156, F_FM0_RDATA(12) => nc280, 
        F_FM0_RDATA(11) => nc125, F_FM0_RDATA(10) => nc211, 
        F_FM0_RDATA(9) => nc73, F_FM0_RDATA(8) => nc107, 
        F_FM0_RDATA(7) => nc66, F_FM0_RDATA(6) => nc83, 
        F_FM0_RDATA(5) => nc9, F_FM0_RDATA(4) => nc252, 
        F_FM0_RDATA(3) => nc171, F_FM0_RDATA(2) => nc54, 
        F_FM0_RDATA(1) => nc286, F_FM0_RDATA(0) => nc307, 
        F_FM0_READYOUT => OPEN, F_FM0_RESP => OPEN, 
        F_HM0_ADDR(31) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31, 
        F_HM0_ADDR(30) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30, 
        F_HM0_ADDR(29) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29, 
        F_HM0_ADDR(28) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28, 
        F_HM0_ADDR(27) => nc135, F_HM0_ADDR(26) => nc41, 
        F_HM0_ADDR(25) => nc100, F_HM0_ADDR(24) => nc270, 
        F_HM0_ADDR(23) => nc52, F_HM0_ADDR(22) => nc251, 
        F_HM0_ADDR(21) => nc186, F_HM0_ADDR(20) => nc29, 
        F_HM0_ADDR(19) => nc269, F_HM0_ADDR(18) => nc118, 
        F_HM0_ADDR(17) => nc60, F_HM0_ADDR(16) => nc141, 
        F_HM0_ADDR(15) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15, 
        F_HM0_ADDR(14) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14, 
        F_HM0_ADDR(13) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13, 
        F_HM0_ADDR(12) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12, 
        F_HM0_ADDR(11) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11, 
        F_HM0_ADDR(10) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10, 
        F_HM0_ADDR(9) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9, 
        F_HM0_ADDR(8) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8, 
        F_HM0_ADDR(7) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7, 
        F_HM0_ADDR(6) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6, 
        F_HM0_ADDR(5) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5, 
        F_HM0_ADDR(4) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4, 
        F_HM0_ADDR(3) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3, 
        F_HM0_ADDR(2) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2, 
        F_HM0_ADDR(1) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1, 
        F_HM0_ADDR(0) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0, 
        F_HM0_ENABLE => OPEN, F_HM0_SEL => OPEN, F_HM0_SIZE(1)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1), 
        F_HM0_SIZE(0) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0), 
        F_HM0_TRANS1 => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1), 
        F_HM0_WDATA(31) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31), 
        F_HM0_WDATA(30) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30), 
        F_HM0_WDATA(29) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29), 
        F_HM0_WDATA(28) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28), 
        F_HM0_WDATA(27) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27), 
        F_HM0_WDATA(26) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26), 
        F_HM0_WDATA(25) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25), 
        F_HM0_WDATA(24) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24), 
        F_HM0_WDATA(23) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23), 
        F_HM0_WDATA(22) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22), 
        F_HM0_WDATA(21) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21), 
        F_HM0_WDATA(20) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20), 
        F_HM0_WDATA(19) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19), 
        F_HM0_WDATA(18) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18), 
        F_HM0_WDATA(17) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17), 
        F_HM0_WDATA(16) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16), 
        F_HM0_WDATA(15) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15), 
        F_HM0_WDATA(14) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14), 
        F_HM0_WDATA(13) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13), 
        F_HM0_WDATA(12) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12), 
        F_HM0_WDATA(11) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11), 
        F_HM0_WDATA(10) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10), 
        F_HM0_WDATA(9) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9), 
        F_HM0_WDATA(8) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8), 
        F_HM0_WDATA(7) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7), 
        F_HM0_WDATA(6) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6), 
        F_HM0_WDATA(5) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5), 
        F_HM0_WDATA(4) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4), 
        F_HM0_WDATA(3) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3), 
        F_HM0_WDATA(2) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2), 
        F_HM0_WDATA(1) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1), 
        F_HM0_WDATA(0) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0), 
        F_HM0_WRITE => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        FAB_CHRGVBUS => OPEN, FAB_DISCHRGVBUS => OPEN, 
        FAB_DMPULLDOWN => OPEN, FAB_DPPULLDOWN => OPEN, 
        FAB_DRVVBUS => OPEN, FAB_IDPULLUP => OPEN, FAB_OPMODE(1)
         => nc311, FAB_OPMODE(0) => nc276, FAB_SUSPENDM => OPEN, 
        FAB_TERMSEL => OPEN, FAB_TXVALID => OPEN, FAB_VCONTROL(3)
         => nc193, FAB_VCONTROL(2) => nc214, FAB_VCONTROL(1) => 
        nc298, FAB_VCONTROL(0) => nc282, FAB_VCONTROLLOADM => 
        OPEN, FAB_XCVRSEL(1) => nc240, FAB_XCVRSEL(0) => nc45, 
        FAB_XDATAOUT(7) => nc53, FAB_XDATAOUT(6) => nc121, 
        FAB_XDATAOUT(5) => nc176, FAB_XDATAOUT(4) => nc220, 
        FAB_XDATAOUT(3) => nc158, FAB_XDATAOUT(2) => nc281, 
        FAB_XDATAOUT(1) => nc209, FAB_XDATAOUT(0) => nc246, 
        FACC_GLMUX_SEL => OPEN, FIC32_0_MASTER(1) => nc162, 
        FIC32_0_MASTER(0) => nc11, FIC32_1_MASTER(1) => nc272, 
        FIC32_1_MASTER(0) => nc131, FPGA_RESET_N => 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, GTX_CLK
         => OPEN, H2F_INTERRUPT(15) => nc254, H2F_INTERRUPT(14)
         => nc267, H2F_INTERRUPT(13) => nc96, H2F_INTERRUPT(12)
         => nc79, H2F_INTERRUPT(11) => nc226, H2F_INTERRUPT(10)
         => nc146, H2F_INTERRUPT(9) => nc230, H2F_INTERRUPT(8)
         => nc89, H2F_INTERRUPT(7) => nc119, H2F_INTERRUPT(6) => 
        nc48, H2F_INTERRUPT(5) => nc271, H2F_INTERRUPT(4) => 
        nc213, H2F_INTERRUPT(3) => nc300, H2F_INTERRUPT(2) => 
        nc126, H2F_INTERRUPT(1) => nc195, H2F_INTERRUPT(0) => 
        nc188, H2F_NMI => OPEN, H2FCALIB => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_A => OPEN, I2C0_SCL_MGPIO31B_H2F_B
         => OPEN, I2C0_SDA_MGPIO30B_H2F_A => OPEN, 
        I2C0_SDA_MGPIO30B_H2F_B => OPEN, I2C1_SCL_MGPIO1A_H2F_A
         => OPEN, I2C1_SCL_MGPIO1A_H2F_B => 
        CertificationSystem_sb_0_GPIO_1_M2F, 
        I2C1_SDA_MGPIO0A_H2F_A => OPEN, I2C1_SDA_MGPIO0A_H2F_B
         => GPIO_0_M2F_c, MDCF => OPEN, MDOENF => OPEN, MDOF => 
        OPEN, MMUART0_CTS_MGPIO19B_H2F_A => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => OPEN, MPLL_LOCK => OPEN, 
        PER2_FABRIC_PADDR(15) => nc242, PER2_FABRIC_PADDR(14) => 
        nc15, PER2_FABRIC_PADDR(13) => nc308, 
        PER2_FABRIC_PADDR(12) => nc236, PER2_FABRIC_PADDR(11) => 
        nc102, PER2_FABRIC_PADDR(10) => nc304, 
        PER2_FABRIC_PADDR(9) => nc3, PER2_FABRIC_PADDR(8) => 
        nc207, PER2_FABRIC_PADDR(7) => nc47, PER2_FABRIC_PADDR(6)
         => nc90, PER2_FABRIC_PADDR(5) => nc284, 
        PER2_FABRIC_PADDR(4) => nc222, PER2_FABRIC_PADDR(3) => 
        nc159, PER2_FABRIC_PADDR(2) => nc136, PER2_FABRIC_PENABLE
         => OPEN, PER2_FABRIC_PSEL => OPEN, 
        PER2_FABRIC_PWDATA(31) => nc241, PER2_FABRIC_PWDATA(30)
         => nc253, PER2_FABRIC_PWDATA(29) => nc178, 
        PER2_FABRIC_PWDATA(28) => nc306, PER2_FABRIC_PWDATA(27)
         => nc215, PER2_FABRIC_PWDATA(26) => nc59, 
        PER2_FABRIC_PWDATA(25) => nc221, PER2_FABRIC_PWDATA(24)
         => nc232, PER2_FABRIC_PWDATA(23) => nc274, 
        PER2_FABRIC_PWDATA(22) => nc18, PER2_FABRIC_PWDATA(21)
         => nc44, PER2_FABRIC_PWDATA(20) => nc117, 
        PER2_FABRIC_PWDATA(19) => nc189, PER2_FABRIC_PWDATA(18)
         => nc164, PER2_FABRIC_PWDATA(17) => nc148, 
        PER2_FABRIC_PWDATA(16) => nc42, PER2_FABRIC_PWDATA(15)
         => nc231, PER2_FABRIC_PWDATA(14) => nc191, 
        PER2_FABRIC_PWDATA(13) => nc255, PER2_FABRIC_PWDATA(12)
         => nc283, PER2_FABRIC_PWDATA(11) => nc317, 
        PER2_FABRIC_PWDATA(10) => nc290, PER2_FABRIC_PWDATA(9)
         => nc17, PER2_FABRIC_PWDATA(8) => nc2, 
        PER2_FABRIC_PWDATA(7) => nc302, PER2_FABRIC_PWDATA(6) => 
        nc110, PER2_FABRIC_PWDATA(5) => nc128, 
        PER2_FABRIC_PWDATA(4) => nc244, PER2_FABRIC_PWDATA(3) => 
        nc321, PER2_FABRIC_PWDATA(2) => nc43, 
        PER2_FABRIC_PWDATA(1) => nc179, PER2_FABRIC_PWDATA(0) => 
        nc157, PER2_FABRIC_PWRITE => OPEN, RTC_MATCH => OPEN, 
        SLEEPDEEP => OPEN, SLEEPHOLDACK => OPEN, SLEEPING => OPEN, 
        SMBALERT_NO0 => OPEN, SMBALERT_NO1 => OPEN, SMBSUS_NO0
         => OPEN, SMBSUS_NO1 => OPEN, SPI0_CLK_OUT => OPEN, 
        SPI0_SDI_MGPIO5A_H2F_A => OPEN, SPI0_SDI_MGPIO5A_H2F_B
         => OPEN, SPI0_SDO_MGPIO6A_H2F_A => OPEN, 
        SPI0_SDO_MGPIO6A_H2F_B => OPEN, SPI0_SS0_MGPIO7A_H2F_A
         => OPEN, SPI0_SS0_MGPIO7A_H2F_B => OPEN, 
        SPI0_SS1_MGPIO8A_H2F_A => OPEN, SPI0_SS1_MGPIO8A_H2F_B
         => OPEN, SPI0_SS2_MGPIO9A_H2F_A => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_B => 
        CertificationSystem_sb_0_GPIO_9_M2F, 
        SPI0_SS3_MGPIO10A_H2F_A => OPEN, SPI0_SS3_MGPIO10A_H2F_B
         => OPEN, SPI0_SS4_MGPIO19A_H2F_A => OPEN, 
        SPI0_SS5_MGPIO20A_H2F_A => OPEN, SPI0_SS6_MGPIO21A_H2F_A
         => OPEN, SPI0_SS7_MGPIO22A_H2F_A => OPEN, SPI1_CLK_OUT
         => OPEN, SPI1_SDI_MGPIO11A_H2F_A => OPEN, 
        SPI1_SDI_MGPIO11A_H2F_B => OPEN, SPI1_SDO_MGPIO12A_H2F_A
         => OPEN, SPI1_SDO_MGPIO12A_H2F_B => OPEN, 
        SPI1_SS0_MGPIO13A_H2F_A => OPEN, SPI1_SS0_MGPIO13A_H2F_B
         => OPEN, SPI1_SS1_MGPIO14A_H2F_A => OPEN, 
        SPI1_SS1_MGPIO14A_H2F_B => OPEN, SPI1_SS2_MGPIO15A_H2F_A
         => OPEN, SPI1_SS2_MGPIO15A_H2F_B => OPEN, 
        SPI1_SS3_MGPIO16A_H2F_A => OPEN, SPI1_SS3_MGPIO16A_H2F_B
         => OPEN, SPI1_SS4_MGPIO17A_H2F_A => OPEN, 
        SPI1_SS5_MGPIO18A_H2F_A => OPEN, SPI1_SS6_MGPIO23A_H2F_A
         => OPEN, SPI1_SS7_MGPIO24A_H2F_A => OPEN, TCGF(9) => 
        nc36, TCGF(8) => nc224, TCGF(7) => nc296, TCGF(6) => 
        nc273, TCGF(5) => nc61, TCGF(4) => nc104, TCGF(3) => 
        nc138, TCGF(2) => nc14, TCGF(1) => nc285, TCGF(0) => 
        nc303, TRACECLK => OPEN, TRACEDATA(3) => nc150, 
        TRACEDATA(2) => nc196, TRACEDATA(1) => nc234, 
        TRACEDATA(0) => nc149, TX_CLK => OPEN, TX_ENF => OPEN, 
        TX_ERRF => OPEN, TXCTL_EN_RIF => OPEN, TXD_RIF(3) => nc12, 
        TXD_RIF(2) => nc219, TXD_RIF(1) => nc30, TXD_RIF(0) => 
        nc243, TXDF(7) => nc187, TXDF(6) => nc65, TXDF(5) => nc7, 
        TXDF(4) => nc292, TXDF(3) => nc129, TXDF(2) => nc275, 
        TXDF(1) => nc8, TXDF(0) => nc223, TXEV => OPEN, 
        WDOGTIMEOUT => OPEN, F_ARREADY_HREADYOUT1 => OPEN, 
        F_AWREADY_HREADYOUT0 => OPEN, F_BID(3) => nc13, F_BID(2)
         => nc305, F_BID(1) => nc180, F_BID(0) => nc26, 
        F_BRESP_HRESP0(1) => nc291, F_BRESP_HRESP0(0) => nc177, 
        F_BVALID => OPEN, F_RDATA_HRDATA01(63) => nc139, 
        F_RDATA_HRDATA01(62) => nc310, F_RDATA_HRDATA01(61) => 
        nc259, F_RDATA_HRDATA01(60) => nc245, 
        F_RDATA_HRDATA01(59) => nc233, F_RDATA_HRDATA01(58) => 
        nc163, F_RDATA_HRDATA01(57) => nc318, 
        F_RDATA_HRDATA01(56) => nc268, F_RDATA_HRDATA01(55) => 
        nc112, F_RDATA_HRDATA01(54) => nc68, F_RDATA_HRDATA01(53)
         => nc49, F_RDATA_HRDATA01(52) => nc314, 
        F_RDATA_HRDATA01(51) => nc217, F_RDATA_HRDATA01(50) => 
        nc170, F_RDATA_HRDATA01(49) => nc91, F_RDATA_HRDATA01(48)
         => nc225, F_RDATA_HRDATA01(47) => nc5, 
        F_RDATA_HRDATA01(46) => nc20, F_RDATA_HRDATA01(45) => 
        nc198, F_RDATA_HRDATA01(44) => nc147, 
        F_RDATA_HRDATA01(43) => nc316, F_RDATA_HRDATA01(42) => 
        nc67, F_RDATA_HRDATA01(41) => nc289, F_RDATA_HRDATA01(40)
         => nc294, F_RDATA_HRDATA01(39) => nc152, 
        F_RDATA_HRDATA01(38) => nc127, F_RDATA_HRDATA01(37) => 
        nc103, F_RDATA_HRDATA01(36) => nc235, 
        F_RDATA_HRDATA01(35) => nc76, F_RDATA_HRDATA01(34) => 
        nc208, F_RDATA_HRDATA01(33) => nc140, 
        F_RDATA_HRDATA01(32) => nc257, F_RDATA_HRDATA01(31) => 
        nc86, F_RDATA_HRDATA01(30) => nc95, F_RDATA_HRDATA01(29)
         => nc120, F_RDATA_HRDATA01(28) => nc165, 
        F_RDATA_HRDATA01(27) => nc279, F_RDATA_HRDATA01(26) => 
        nc137, F_RDATA_HRDATA01(25) => nc64, F_RDATA_HRDATA01(24)
         => nc19, F_RDATA_HRDATA01(23) => nc312, 
        F_RDATA_HRDATA01(22) => nc70, F_RDATA_HRDATA01(21) => 
        nc182, F_RDATA_HRDATA01(20) => nc62, F_RDATA_HRDATA01(19)
         => nc199, F_RDATA_HRDATA01(18) => nc80, 
        F_RDATA_HRDATA01(17) => nc130, F_RDATA_HRDATA01(16) => 
        nc287, F_RDATA_HRDATA01(15) => nc98, F_RDATA_HRDATA01(14)
         => nc293, F_RDATA_HRDATA01(13) => nc249, 
        F_RDATA_HRDATA01(12) => nc114, F_RDATA_HRDATA01(11) => 
        nc56, F_RDATA_HRDATA01(10) => nc105, F_RDATA_HRDATA01(9)
         => nc63, F_RDATA_HRDATA01(8) => nc313, 
        F_RDATA_HRDATA01(7) => nc309, F_RDATA_HRDATA01(6) => 
        nc172, F_RDATA_HRDATA01(5) => nc229, F_RDATA_HRDATA01(4)
         => nc277, F_RDATA_HRDATA01(3) => nc97, 
        F_RDATA_HRDATA01(2) => nc161, F_RDATA_HRDATA01(1) => nc31, 
        F_RDATA_HRDATA01(0) => nc295, F_RID(3) => nc154, F_RID(2)
         => nc50, F_RID(1) => nc260, F_RID(0) => nc239, F_RLAST
         => OPEN, F_RRESP_HRESP1(1) => nc142, F_RRESP_HRESP1(0)
         => nc320, F_RVALID => OPEN, F_WREADY => OPEN, 
        MDDR_FABRIC_PRDATA(15) => nc315, MDDR_FABRIC_PRDATA(14)
         => nc247, MDDR_FABRIC_PRDATA(13) => nc94, 
        MDDR_FABRIC_PRDATA(12) => nc197, MDDR_FABRIC_PRDATA(11)
         => nc122, MDDR_FABRIC_PRDATA(10) => nc266, 
        MDDR_FABRIC_PRDATA(9) => nc35, MDDR_FABRIC_PRDATA(8) => 
        nc4, MDDR_FABRIC_PRDATA(7) => nc227, 
        MDDR_FABRIC_PRDATA(6) => nc92, MDDR_FABRIC_PRDATA(5) => 
        nc101, MDDR_FABRIC_PRDATA(4) => nc184, 
        MDDR_FABRIC_PRDATA(3) => nc200, MDDR_FABRIC_PRDATA(2) => 
        nc190, MDDR_FABRIC_PRDATA(1) => nc166, 
        MDDR_FABRIC_PRDATA(0) => nc132, MDDR_FABRIC_PREADY => 
        OPEN, MDDR_FABRIC_PSLVERR => OPEN, CAN_RXBUS_F2H_SCP => 
        VCC_net_1, CAN_TX_EBL_F2H_SCP => VCC_net_1, 
        CAN_TXBUS_F2H_SCP => VCC_net_1, COLF => VCC_net_1, CRSF
         => VCC_net_1, F2_DMAREADY(1) => VCC_net_1, 
        F2_DMAREADY(0) => VCC_net_1, F2H_INTERRUPT(15) => 
        GND_net_1, F2H_INTERRUPT(14) => GND_net_1, 
        F2H_INTERRUPT(13) => GND_net_1, F2H_INTERRUPT(12) => 
        GND_net_1, F2H_INTERRUPT(11) => GND_net_1, 
        F2H_INTERRUPT(10) => GND_net_1, F2H_INTERRUPT(9) => 
        GND_net_1, F2H_INTERRUPT(8) => GND_net_1, 
        F2H_INTERRUPT(7) => GND_net_1, F2H_INTERRUPT(6) => 
        GND_net_1, F2H_INTERRUPT(5) => GND_net_1, 
        F2H_INTERRUPT(4) => GND_net_1, F2H_INTERRUPT(3) => 
        GND_net_1, F2H_INTERRUPT(2) => GND_net_1, 
        F2H_INTERRUPT(1) => GND_net_1, F2H_INTERRUPT(0) => 
        GND_net_1, F2HCALIB => VCC_net_1, F_DMAREADY(1) => 
        VCC_net_1, F_DMAREADY(0) => VCC_net_1, F_FM0_ADDR(31) => 
        GND_net_1, F_FM0_ADDR(30) => GND_net_1, F_FM0_ADDR(29)
         => GND_net_1, F_FM0_ADDR(28) => GND_net_1, 
        F_FM0_ADDR(27) => GND_net_1, F_FM0_ADDR(26) => GND_net_1, 
        F_FM0_ADDR(25) => GND_net_1, F_FM0_ADDR(24) => GND_net_1, 
        F_FM0_ADDR(23) => GND_net_1, F_FM0_ADDR(22) => GND_net_1, 
        F_FM0_ADDR(21) => GND_net_1, F_FM0_ADDR(20) => GND_net_1, 
        F_FM0_ADDR(19) => GND_net_1, F_FM0_ADDR(18) => GND_net_1, 
        F_FM0_ADDR(17) => GND_net_1, F_FM0_ADDR(16) => GND_net_1, 
        F_FM0_ADDR(15) => GND_net_1, F_FM0_ADDR(14) => GND_net_1, 
        F_FM0_ADDR(13) => GND_net_1, F_FM0_ADDR(12) => GND_net_1, 
        F_FM0_ADDR(11) => GND_net_1, F_FM0_ADDR(10) => GND_net_1, 
        F_FM0_ADDR(9) => GND_net_1, F_FM0_ADDR(8) => GND_net_1, 
        F_FM0_ADDR(7) => GND_net_1, F_FM0_ADDR(6) => GND_net_1, 
        F_FM0_ADDR(5) => GND_net_1, F_FM0_ADDR(4) => GND_net_1, 
        F_FM0_ADDR(3) => GND_net_1, F_FM0_ADDR(2) => GND_net_1, 
        F_FM0_ADDR(1) => GND_net_1, F_FM0_ADDR(0) => GND_net_1, 
        F_FM0_ENABLE => GND_net_1, F_FM0_MASTLOCK => GND_net_1, 
        F_FM0_READY => VCC_net_1, F_FM0_SEL => GND_net_1, 
        F_FM0_SIZE(1) => GND_net_1, F_FM0_SIZE(0) => GND_net_1, 
        F_FM0_TRANS1 => GND_net_1, F_FM0_WDATA(31) => GND_net_1, 
        F_FM0_WDATA(30) => GND_net_1, F_FM0_WDATA(29) => 
        GND_net_1, F_FM0_WDATA(28) => GND_net_1, F_FM0_WDATA(27)
         => GND_net_1, F_FM0_WDATA(26) => GND_net_1, 
        F_FM0_WDATA(25) => GND_net_1, F_FM0_WDATA(24) => 
        GND_net_1, F_FM0_WDATA(23) => GND_net_1, F_FM0_WDATA(22)
         => GND_net_1, F_FM0_WDATA(21) => GND_net_1, 
        F_FM0_WDATA(20) => GND_net_1, F_FM0_WDATA(19) => 
        GND_net_1, F_FM0_WDATA(18) => GND_net_1, F_FM0_WDATA(17)
         => GND_net_1, F_FM0_WDATA(16) => GND_net_1, 
        F_FM0_WDATA(15) => GND_net_1, F_FM0_WDATA(14) => 
        GND_net_1, F_FM0_WDATA(13) => GND_net_1, F_FM0_WDATA(12)
         => GND_net_1, F_FM0_WDATA(11) => GND_net_1, 
        F_FM0_WDATA(10) => GND_net_1, F_FM0_WDATA(9) => GND_net_1, 
        F_FM0_WDATA(8) => GND_net_1, F_FM0_WDATA(7) => GND_net_1, 
        F_FM0_WDATA(6) => GND_net_1, F_FM0_WDATA(5) => GND_net_1, 
        F_FM0_WDATA(4) => GND_net_1, F_FM0_WDATA(3) => GND_net_1, 
        F_FM0_WDATA(2) => GND_net_1, F_FM0_WDATA(1) => GND_net_1, 
        F_FM0_WDATA(0) => GND_net_1, F_FM0_WRITE => GND_net_1, 
        F_HM0_RDATA(31) => N_477_i_0, F_HM0_RDATA(30) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30, 
        F_HM0_RDATA(29) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29, 
        F_HM0_RDATA(28) => N_478_i_0, F_HM0_RDATA(27) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27, 
        F_HM0_RDATA(26) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26, 
        F_HM0_RDATA(25) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25, 
        F_HM0_RDATA(24) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24, 
        F_HM0_RDATA(23) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23, 
        F_HM0_RDATA(22) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22, 
        F_HM0_RDATA(21) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21, 
        F_HM0_RDATA(20) => N_479_i_0, F_HM0_RDATA(19) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19, 
        F_HM0_RDATA(18) => N_480_i_0, F_HM0_RDATA(17) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17, 
        F_HM0_RDATA(16) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16, 
        F_HM0_RDATA(15) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15, 
        F_HM0_RDATA(14) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14, 
        F_HM0_RDATA(13) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13, 
        F_HM0_RDATA(12) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12, 
        F_HM0_RDATA(11) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11, 
        F_HM0_RDATA(10) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10, 
        F_HM0_RDATA(9) => N_481_i_0, F_HM0_RDATA(8) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8, 
        F_HM0_RDATA(7) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7, 
        F_HM0_RDATA(6) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6, 
        F_HM0_RDATA(5) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5, 
        F_HM0_RDATA(4) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4, 
        F_HM0_RDATA(3) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3, 
        F_HM0_RDATA(2) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2, 
        F_HM0_RDATA(1) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1, 
        F_HM0_RDATA(0) => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0, 
        F_HM0_READY => N_9_i_0, F_HM0_RESP => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        FAB_AVALID => VCC_net_1, FAB_HOSTDISCON => VCC_net_1, 
        FAB_IDDIG => VCC_net_1, FAB_LINESTATE(1) => VCC_net_1, 
        FAB_LINESTATE(0) => VCC_net_1, FAB_M3_RESET_N => 
        VCC_net_1, FAB_PLL_LOCK => FAB_CCC_LOCK, FAB_RXACTIVE => 
        VCC_net_1, FAB_RXERROR => VCC_net_1, FAB_RXVALID => 
        VCC_net_1, FAB_RXVALIDH => GND_net_1, FAB_SESSEND => 
        VCC_net_1, FAB_TXREADY => VCC_net_1, FAB_VBUSVALID => 
        VCC_net_1, FAB_VSTATUS(7) => VCC_net_1, FAB_VSTATUS(6)
         => VCC_net_1, FAB_VSTATUS(5) => VCC_net_1, 
        FAB_VSTATUS(4) => VCC_net_1, FAB_VSTATUS(3) => VCC_net_1, 
        FAB_VSTATUS(2) => VCC_net_1, FAB_VSTATUS(1) => VCC_net_1, 
        FAB_VSTATUS(0) => VCC_net_1, FAB_XDATAIN(7) => VCC_net_1, 
        FAB_XDATAIN(6) => VCC_net_1, FAB_XDATAIN(5) => VCC_net_1, 
        FAB_XDATAIN(4) => VCC_net_1, FAB_XDATAIN(3) => VCC_net_1, 
        FAB_XDATAIN(2) => VCC_net_1, FAB_XDATAIN(1) => VCC_net_1, 
        FAB_XDATAIN(0) => VCC_net_1, GTX_CLKPF => VCC_net_1, 
        I2C0_BCLK => VCC_net_1, I2C0_SCL_F2H_SCP => VCC_net_1, 
        I2C0_SDA_F2H_SCP => VCC_net_1, I2C1_BCLK => VCC_net_1, 
        I2C1_SCL_F2H_SCP => VCC_net_1, I2C1_SDA_F2H_SCP => 
        VCC_net_1, MDIF => VCC_net_1, MGPIO0A_F2H_GPIN => 
        VCC_net_1, MGPIO10A_F2H_GPIN => VCC_net_1, 
        MGPIO11A_F2H_GPIN => VCC_net_1, MGPIO11B_F2H_GPIN => 
        VCC_net_1, MGPIO12A_F2H_GPIN => VCC_net_1, 
        MGPIO13A_F2H_GPIN => VCC_net_1, MGPIO14A_F2H_GPIN => 
        VCC_net_1, MGPIO15A_F2H_GPIN => VCC_net_1, 
        MGPIO16A_F2H_GPIN => VCC_net_1, MGPIO17B_F2H_GPIN => 
        VCC_net_1, MGPIO18B_F2H_GPIN => VCC_net_1, 
        MGPIO19B_F2H_GPIN => VCC_net_1, MGPIO1A_F2H_GPIN => 
        VCC_net_1, MGPIO20B_F2H_GPIN => VCC_net_1, 
        MGPIO21B_F2H_GPIN => VCC_net_1, MGPIO22B_F2H_GPIN => 
        VCC_net_1, MGPIO24B_F2H_GPIN => VCC_net_1, 
        MGPIO25B_F2H_GPIN => VCC_net_1, MGPIO26B_F2H_GPIN => 
        VCC_net_1, MGPIO27B_F2H_GPIN => VCC_net_1, 
        MGPIO28B_F2H_GPIN => VCC_net_1, MGPIO29B_F2H_GPIN => 
        VCC_net_1, MGPIO2A_F2H_GPIN => 
        SHA256_Module_0_waiting_data, MGPIO30B_F2H_GPIN => 
        VCC_net_1, MGPIO31B_F2H_GPIN => VCC_net_1, 
        MGPIO3A_F2H_GPIN => 
        SHA256_Module_0_data_available_lastbank_8, 
        MGPIO4A_F2H_GPIN => SHA256_Module_0_di_req_o, 
        MGPIO5A_F2H_GPIN => GND_net_1, MGPIO6A_F2H_GPIN => 
        SHA256_Module_0_do_valid_o, MGPIO7A_F2H_GPIN => 
        SHA256_Module_0_data_available, MGPIO8A_F2H_GPIN => 
        SHA256_Module_0_error_o, MGPIO9A_F2H_GPIN => VCC_net_1, 
        MMUART0_CTS_F2H_SCP => VCC_net_1, MMUART0_DCD_F2H_SCP => 
        VCC_net_1, MMUART0_DSR_F2H_SCP => VCC_net_1, 
        MMUART0_DTR_F2H_SCP => VCC_net_1, MMUART0_RI_F2H_SCP => 
        VCC_net_1, MMUART0_RTS_F2H_SCP => VCC_net_1, 
        MMUART0_RXD_F2H_SCP => VCC_net_1, MMUART0_SCK_F2H_SCP => 
        VCC_net_1, MMUART0_TXD_F2H_SCP => VCC_net_1, 
        MMUART1_CTS_F2H_SCP => VCC_net_1, MMUART1_DCD_F2H_SCP => 
        VCC_net_1, MMUART1_DSR_F2H_SCP => VCC_net_1, 
        MMUART1_RI_F2H_SCP => VCC_net_1, MMUART1_RTS_F2H_SCP => 
        VCC_net_1, MMUART1_RXD_F2H_SCP => VCC_net_1, 
        MMUART1_SCK_F2H_SCP => VCC_net_1, MMUART1_TXD_F2H_SCP => 
        VCC_net_1, PER2_FABRIC_PRDATA(31) => GND_net_1, 
        PER2_FABRIC_PRDATA(30) => GND_net_1, 
        PER2_FABRIC_PRDATA(29) => GND_net_1, 
        PER2_FABRIC_PRDATA(28) => GND_net_1, 
        PER2_FABRIC_PRDATA(27) => GND_net_1, 
        PER2_FABRIC_PRDATA(26) => GND_net_1, 
        PER2_FABRIC_PRDATA(25) => GND_net_1, 
        PER2_FABRIC_PRDATA(24) => GND_net_1, 
        PER2_FABRIC_PRDATA(23) => GND_net_1, 
        PER2_FABRIC_PRDATA(22) => GND_net_1, 
        PER2_FABRIC_PRDATA(21) => GND_net_1, 
        PER2_FABRIC_PRDATA(20) => GND_net_1, 
        PER2_FABRIC_PRDATA(19) => GND_net_1, 
        PER2_FABRIC_PRDATA(18) => GND_net_1, 
        PER2_FABRIC_PRDATA(17) => GND_net_1, 
        PER2_FABRIC_PRDATA(16) => GND_net_1, 
        PER2_FABRIC_PRDATA(15) => GND_net_1, 
        PER2_FABRIC_PRDATA(14) => GND_net_1, 
        PER2_FABRIC_PRDATA(13) => GND_net_1, 
        PER2_FABRIC_PRDATA(12) => GND_net_1, 
        PER2_FABRIC_PRDATA(11) => GND_net_1, 
        PER2_FABRIC_PRDATA(10) => GND_net_1, 
        PER2_FABRIC_PRDATA(9) => GND_net_1, PER2_FABRIC_PRDATA(8)
         => GND_net_1, PER2_FABRIC_PRDATA(7) => GND_net_1, 
        PER2_FABRIC_PRDATA(6) => GND_net_1, PER2_FABRIC_PRDATA(5)
         => GND_net_1, PER2_FABRIC_PRDATA(4) => GND_net_1, 
        PER2_FABRIC_PRDATA(3) => GND_net_1, PER2_FABRIC_PRDATA(2)
         => GND_net_1, PER2_FABRIC_PRDATA(1) => GND_net_1, 
        PER2_FABRIC_PRDATA(0) => GND_net_1, PER2_FABRIC_PREADY
         => VCC_net_1, PER2_FABRIC_PSLVERR => GND_net_1, RCGF(9)
         => VCC_net_1, RCGF(8) => VCC_net_1, RCGF(7) => VCC_net_1, 
        RCGF(6) => VCC_net_1, RCGF(5) => VCC_net_1, RCGF(4) => 
        VCC_net_1, RCGF(3) => VCC_net_1, RCGF(2) => VCC_net_1, 
        RCGF(1) => VCC_net_1, RCGF(0) => VCC_net_1, RX_CLKPF => 
        VCC_net_1, RX_DVF => VCC_net_1, RX_ERRF => VCC_net_1, 
        RX_EV => VCC_net_1, RXDF(7) => VCC_net_1, RXDF(6) => 
        VCC_net_1, RXDF(5) => VCC_net_1, RXDF(4) => VCC_net_1, 
        RXDF(3) => VCC_net_1, RXDF(2) => VCC_net_1, RXDF(1) => 
        VCC_net_1, RXDF(0) => VCC_net_1, SLEEPHOLDREQ => 
        GND_net_1, SMBALERT_NI0 => VCC_net_1, SMBALERT_NI1 => 
        VCC_net_1, SMBSUS_NI0 => VCC_net_1, SMBSUS_NI1 => 
        VCC_net_1, SPI0_CLK_IN => VCC_net_1, SPI0_SDI_F2H_SCP => 
        VCC_net_1, SPI0_SDO_F2H_SCP => VCC_net_1, 
        SPI0_SS0_F2H_SCP => VCC_net_1, SPI0_SS1_F2H_SCP => 
        VCC_net_1, SPI0_SS2_F2H_SCP => VCC_net_1, 
        SPI0_SS3_F2H_SCP => VCC_net_1, SPI1_CLK_IN => VCC_net_1, 
        SPI1_SDI_F2H_SCP => VCC_net_1, SPI1_SDO_F2H_SCP => 
        VCC_net_1, SPI1_SS0_F2H_SCP => VCC_net_1, 
        SPI1_SS1_F2H_SCP => VCC_net_1, SPI1_SS2_F2H_SCP => 
        VCC_net_1, SPI1_SS3_F2H_SCP => VCC_net_1, TX_CLKPF => 
        VCC_net_1, USER_MSS_GPIO_RESET_N => VCC_net_1, 
        USER_MSS_RESET_N => VCC_net_1, XCLK_FAB => VCC_net_1, 
        CLK_BASE => CertificationSystem_sb_0_FAB_CCC_GL0, 
        CLK_MDDR_APB => VCC_net_1, F_ARADDR_HADDR1(31) => 
        VCC_net_1, F_ARADDR_HADDR1(30) => VCC_net_1, 
        F_ARADDR_HADDR1(29) => VCC_net_1, F_ARADDR_HADDR1(28) => 
        VCC_net_1, F_ARADDR_HADDR1(27) => VCC_net_1, 
        F_ARADDR_HADDR1(26) => VCC_net_1, F_ARADDR_HADDR1(25) => 
        VCC_net_1, F_ARADDR_HADDR1(24) => VCC_net_1, 
        F_ARADDR_HADDR1(23) => VCC_net_1, F_ARADDR_HADDR1(22) => 
        VCC_net_1, F_ARADDR_HADDR1(21) => VCC_net_1, 
        F_ARADDR_HADDR1(20) => VCC_net_1, F_ARADDR_HADDR1(19) => 
        VCC_net_1, F_ARADDR_HADDR1(18) => VCC_net_1, 
        F_ARADDR_HADDR1(17) => VCC_net_1, F_ARADDR_HADDR1(16) => 
        VCC_net_1, F_ARADDR_HADDR1(15) => VCC_net_1, 
        F_ARADDR_HADDR1(14) => VCC_net_1, F_ARADDR_HADDR1(13) => 
        VCC_net_1, F_ARADDR_HADDR1(12) => VCC_net_1, 
        F_ARADDR_HADDR1(11) => VCC_net_1, F_ARADDR_HADDR1(10) => 
        VCC_net_1, F_ARADDR_HADDR1(9) => VCC_net_1, 
        F_ARADDR_HADDR1(8) => VCC_net_1, F_ARADDR_HADDR1(7) => 
        VCC_net_1, F_ARADDR_HADDR1(6) => VCC_net_1, 
        F_ARADDR_HADDR1(5) => VCC_net_1, F_ARADDR_HADDR1(4) => 
        VCC_net_1, F_ARADDR_HADDR1(3) => VCC_net_1, 
        F_ARADDR_HADDR1(2) => VCC_net_1, F_ARADDR_HADDR1(1) => 
        VCC_net_1, F_ARADDR_HADDR1(0) => VCC_net_1, 
        F_ARBURST_HTRANS1(1) => GND_net_1, F_ARBURST_HTRANS1(0)
         => GND_net_1, F_ARID_HSEL1(3) => GND_net_1, 
        F_ARID_HSEL1(2) => GND_net_1, F_ARID_HSEL1(1) => 
        GND_net_1, F_ARID_HSEL1(0) => GND_net_1, 
        F_ARLEN_HBURST1(3) => GND_net_1, F_ARLEN_HBURST1(2) => 
        GND_net_1, F_ARLEN_HBURST1(1) => GND_net_1, 
        F_ARLEN_HBURST1(0) => GND_net_1, F_ARLOCK_HMASTLOCK1(1)
         => GND_net_1, F_ARLOCK_HMASTLOCK1(0) => GND_net_1, 
        F_ARSIZE_HSIZE1(1) => GND_net_1, F_ARSIZE_HSIZE1(0) => 
        GND_net_1, F_ARVALID_HWRITE1 => GND_net_1, 
        F_AWADDR_HADDR0(31) => VCC_net_1, F_AWADDR_HADDR0(30) => 
        VCC_net_1, F_AWADDR_HADDR0(29) => VCC_net_1, 
        F_AWADDR_HADDR0(28) => VCC_net_1, F_AWADDR_HADDR0(27) => 
        VCC_net_1, F_AWADDR_HADDR0(26) => VCC_net_1, 
        F_AWADDR_HADDR0(25) => VCC_net_1, F_AWADDR_HADDR0(24) => 
        VCC_net_1, F_AWADDR_HADDR0(23) => VCC_net_1, 
        F_AWADDR_HADDR0(22) => VCC_net_1, F_AWADDR_HADDR0(21) => 
        VCC_net_1, F_AWADDR_HADDR0(20) => VCC_net_1, 
        F_AWADDR_HADDR0(19) => VCC_net_1, F_AWADDR_HADDR0(18) => 
        VCC_net_1, F_AWADDR_HADDR0(17) => VCC_net_1, 
        F_AWADDR_HADDR0(16) => VCC_net_1, F_AWADDR_HADDR0(15) => 
        VCC_net_1, F_AWADDR_HADDR0(14) => VCC_net_1, 
        F_AWADDR_HADDR0(13) => VCC_net_1, F_AWADDR_HADDR0(12) => 
        VCC_net_1, F_AWADDR_HADDR0(11) => VCC_net_1, 
        F_AWADDR_HADDR0(10) => VCC_net_1, F_AWADDR_HADDR0(9) => 
        VCC_net_1, F_AWADDR_HADDR0(8) => VCC_net_1, 
        F_AWADDR_HADDR0(7) => VCC_net_1, F_AWADDR_HADDR0(6) => 
        VCC_net_1, F_AWADDR_HADDR0(5) => VCC_net_1, 
        F_AWADDR_HADDR0(4) => VCC_net_1, F_AWADDR_HADDR0(3) => 
        VCC_net_1, F_AWADDR_HADDR0(2) => VCC_net_1, 
        F_AWADDR_HADDR0(1) => VCC_net_1, F_AWADDR_HADDR0(0) => 
        VCC_net_1, F_AWBURST_HTRANS0(1) => GND_net_1, 
        F_AWBURST_HTRANS0(0) => GND_net_1, F_AWID_HSEL0(3) => 
        GND_net_1, F_AWID_HSEL0(2) => GND_net_1, F_AWID_HSEL0(1)
         => GND_net_1, F_AWID_HSEL0(0) => GND_net_1, 
        F_AWLEN_HBURST0(3) => GND_net_1, F_AWLEN_HBURST0(2) => 
        GND_net_1, F_AWLEN_HBURST0(1) => GND_net_1, 
        F_AWLEN_HBURST0(0) => GND_net_1, F_AWLOCK_HMASTLOCK0(1)
         => GND_net_1, F_AWLOCK_HMASTLOCK0(0) => GND_net_1, 
        F_AWSIZE_HSIZE0(1) => GND_net_1, F_AWSIZE_HSIZE0(0) => 
        GND_net_1, F_AWVALID_HWRITE0 => GND_net_1, F_BREADY => 
        GND_net_1, F_RMW_AXI => GND_net_1, F_RREADY => GND_net_1, 
        F_WDATA_HWDATA01(63) => VCC_net_1, F_WDATA_HWDATA01(62)
         => VCC_net_1, F_WDATA_HWDATA01(61) => VCC_net_1, 
        F_WDATA_HWDATA01(60) => VCC_net_1, F_WDATA_HWDATA01(59)
         => VCC_net_1, F_WDATA_HWDATA01(58) => VCC_net_1, 
        F_WDATA_HWDATA01(57) => VCC_net_1, F_WDATA_HWDATA01(56)
         => VCC_net_1, F_WDATA_HWDATA01(55) => VCC_net_1, 
        F_WDATA_HWDATA01(54) => VCC_net_1, F_WDATA_HWDATA01(53)
         => VCC_net_1, F_WDATA_HWDATA01(52) => VCC_net_1, 
        F_WDATA_HWDATA01(51) => VCC_net_1, F_WDATA_HWDATA01(50)
         => VCC_net_1, F_WDATA_HWDATA01(49) => VCC_net_1, 
        F_WDATA_HWDATA01(48) => VCC_net_1, F_WDATA_HWDATA01(47)
         => VCC_net_1, F_WDATA_HWDATA01(46) => VCC_net_1, 
        F_WDATA_HWDATA01(45) => VCC_net_1, F_WDATA_HWDATA01(44)
         => VCC_net_1, F_WDATA_HWDATA01(43) => VCC_net_1, 
        F_WDATA_HWDATA01(42) => VCC_net_1, F_WDATA_HWDATA01(41)
         => VCC_net_1, F_WDATA_HWDATA01(40) => VCC_net_1, 
        F_WDATA_HWDATA01(39) => VCC_net_1, F_WDATA_HWDATA01(38)
         => VCC_net_1, F_WDATA_HWDATA01(37) => VCC_net_1, 
        F_WDATA_HWDATA01(36) => VCC_net_1, F_WDATA_HWDATA01(35)
         => VCC_net_1, F_WDATA_HWDATA01(34) => VCC_net_1, 
        F_WDATA_HWDATA01(33) => VCC_net_1, F_WDATA_HWDATA01(32)
         => VCC_net_1, F_WDATA_HWDATA01(31) => VCC_net_1, 
        F_WDATA_HWDATA01(30) => VCC_net_1, F_WDATA_HWDATA01(29)
         => VCC_net_1, F_WDATA_HWDATA01(28) => VCC_net_1, 
        F_WDATA_HWDATA01(27) => VCC_net_1, F_WDATA_HWDATA01(26)
         => VCC_net_1, F_WDATA_HWDATA01(25) => VCC_net_1, 
        F_WDATA_HWDATA01(24) => VCC_net_1, F_WDATA_HWDATA01(23)
         => VCC_net_1, F_WDATA_HWDATA01(22) => VCC_net_1, 
        F_WDATA_HWDATA01(21) => VCC_net_1, F_WDATA_HWDATA01(20)
         => VCC_net_1, F_WDATA_HWDATA01(19) => VCC_net_1, 
        F_WDATA_HWDATA01(18) => VCC_net_1, F_WDATA_HWDATA01(17)
         => VCC_net_1, F_WDATA_HWDATA01(16) => VCC_net_1, 
        F_WDATA_HWDATA01(15) => VCC_net_1, F_WDATA_HWDATA01(14)
         => VCC_net_1, F_WDATA_HWDATA01(13) => VCC_net_1, 
        F_WDATA_HWDATA01(12) => VCC_net_1, F_WDATA_HWDATA01(11)
         => VCC_net_1, F_WDATA_HWDATA01(10) => VCC_net_1, 
        F_WDATA_HWDATA01(9) => VCC_net_1, F_WDATA_HWDATA01(8) => 
        VCC_net_1, F_WDATA_HWDATA01(7) => VCC_net_1, 
        F_WDATA_HWDATA01(6) => VCC_net_1, F_WDATA_HWDATA01(5) => 
        VCC_net_1, F_WDATA_HWDATA01(4) => VCC_net_1, 
        F_WDATA_HWDATA01(3) => VCC_net_1, F_WDATA_HWDATA01(2) => 
        VCC_net_1, F_WDATA_HWDATA01(1) => VCC_net_1, 
        F_WDATA_HWDATA01(0) => VCC_net_1, F_WID_HREADY01(3) => 
        GND_net_1, F_WID_HREADY01(2) => GND_net_1, 
        F_WID_HREADY01(1) => GND_net_1, F_WID_HREADY01(0) => 
        GND_net_1, F_WLAST => GND_net_1, F_WSTRB(7) => GND_net_1, 
        F_WSTRB(6) => GND_net_1, F_WSTRB(5) => GND_net_1, 
        F_WSTRB(4) => GND_net_1, F_WSTRB(3) => GND_net_1, 
        F_WSTRB(2) => GND_net_1, F_WSTRB(1) => GND_net_1, 
        F_WSTRB(0) => GND_net_1, F_WVALID => GND_net_1, 
        FPGA_MDDR_ARESET_N => VCC_net_1, MDDR_FABRIC_PADDR(10)
         => VCC_net_1, MDDR_FABRIC_PADDR(9) => VCC_net_1, 
        MDDR_FABRIC_PADDR(8) => VCC_net_1, MDDR_FABRIC_PADDR(7)
         => VCC_net_1, MDDR_FABRIC_PADDR(6) => VCC_net_1, 
        MDDR_FABRIC_PADDR(5) => VCC_net_1, MDDR_FABRIC_PADDR(4)
         => VCC_net_1, MDDR_FABRIC_PADDR(3) => VCC_net_1, 
        MDDR_FABRIC_PADDR(2) => VCC_net_1, MDDR_FABRIC_PENABLE
         => VCC_net_1, MDDR_FABRIC_PSEL => VCC_net_1, 
        MDDR_FABRIC_PWDATA(15) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(14) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(13) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(12) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(11) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(10) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(9) => VCC_net_1, MDDR_FABRIC_PWDATA(8)
         => VCC_net_1, MDDR_FABRIC_PWDATA(7) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(6) => VCC_net_1, MDDR_FABRIC_PWDATA(5)
         => VCC_net_1, MDDR_FABRIC_PWDATA(4) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(3) => VCC_net_1, MDDR_FABRIC_PWDATA(2)
         => VCC_net_1, MDDR_FABRIC_PWDATA(1) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(0) => VCC_net_1, MDDR_FABRIC_PWRITE
         => VCC_net_1, PRESET_N => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => GND_net_1, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => GND_net_1, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => GND_net_1, DM_IN(2)
         => GND_net_1, DM_IN(1) => GND_net_1, DM_IN(0) => 
        GND_net_1, DRAM_DQ_IN(17) => GND_net_1, DRAM_DQ_IN(16)
         => GND_net_1, DRAM_DQ_IN(15) => GND_net_1, 
        DRAM_DQ_IN(14) => GND_net_1, DRAM_DQ_IN(13) => GND_net_1, 
        DRAM_DQ_IN(12) => GND_net_1, DRAM_DQ_IN(11) => GND_net_1, 
        DRAM_DQ_IN(10) => GND_net_1, DRAM_DQ_IN(9) => GND_net_1, 
        DRAM_DQ_IN(8) => GND_net_1, DRAM_DQ_IN(7) => GND_net_1, 
        DRAM_DQ_IN(6) => GND_net_1, DRAM_DQ_IN(5) => GND_net_1, 
        DRAM_DQ_IN(4) => GND_net_1, DRAM_DQ_IN(3) => GND_net_1, 
        DRAM_DQ_IN(2) => GND_net_1, DRAM_DQ_IN(1) => GND_net_1, 
        DRAM_DQ_IN(0) => GND_net_1, DRAM_DQS_IN(2) => GND_net_1, 
        DRAM_DQS_IN(1) => GND_net_1, DRAM_DQS_IN(0) => GND_net_1, 
        DRAM_FIFO_WE_IN(1) => GND_net_1, DRAM_FIFO_WE_IN(0) => 
        GND_net_1, I2C0_SCL_USBC_DATA1_MGPIO31B_IN => GND_net_1, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => GND_net_1, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => GND_net_1, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => GND_net_1, MGPIO0B_IN
         => GND_net_1, MGPIO10B_IN => GND_net_1, MGPIO1B_IN => 
        GND_net_1, MGPIO25A_IN => GND_net_1, MGPIO26A_IN => 
        GND_net_1, MGPIO27A_IN => GND_net_1, MGPIO28A_IN => 
        GND_net_1, MGPIO29A_IN => GND_net_1, MGPIO2B_IN => 
        GND_net_1, MGPIO30A_IN => GND_net_1, MGPIO31A_IN => 
        GND_net_1, MGPIO3B_IN => GND_net_1, MGPIO4B_IN => 
        GND_net_1, MGPIO5B_IN => GND_net_1, MGPIO6B_IN => 
        GND_net_1, MGPIO7B_IN => GND_net_1, MGPIO8B_IN => 
        GND_net_1, MGPIO9B_IN => GND_net_1, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => GND_net_1, 
        MMUART0_DCD_MGPIO22B_IN => GND_net_1, 
        MMUART0_DSR_MGPIO20B_IN => GND_net_1, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => GND_net_1, 
        MMUART0_RI_MGPIO21B_IN => GND_net_1, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => GND_net_1, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => GND_net_1, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => GND_net_1, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => GND_net_1, 
        MMUART1_CTS_MGPIO13B_IN => GND_net_1, 
        MMUART1_DCD_MGPIO16B_IN => GND_net_1, 
        MMUART1_DSR_MGPIO14B_IN => GND_net_1, 
        MMUART1_DTR_MGPIO12B_IN => GND_net_1, 
        MMUART1_RI_MGPIO15B_IN => GND_net_1, 
        MMUART1_RTS_MGPIO11B_IN => GND_net_1, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => MMUART_1_RXD_PAD_Y, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => GND_net_1, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => GND_net_1, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => GND_net_1, 
        RGMII_MDC_RMII_MDC_IN => GND_net_1, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => GND_net_1, 
        RGMII_RX_CLK_IN => GND_net_1, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => GND_net_1, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => GND_net_1, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => GND_net_1, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => GND_net_1, 
        RGMII_RXD3_USBB_DATA4_IN => GND_net_1, RGMII_TX_CLK_IN
         => GND_net_1, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => 
        GND_net_1, RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => GND_net_1, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => GND_net_1, 
        RGMII_TXD2_USBB_DATA5_IN => GND_net_1, 
        RGMII_TXD3_USBB_DATA6_IN => GND_net_1, 
        SPI0_SCK_USBA_XCLK_IN => SPI_0_CLK_PAD_Y, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => SPI_0_DI_PAD_Y, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => GND_net_1, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => SPI_0_SS0_PAD_Y, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => GND_net_1, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => GND_net_1, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => GND_net_1, 
        SPI0_SS4_MGPIO19A_IN => GND_net_1, SPI0_SS5_MGPIO20A_IN
         => GND_net_1, SPI0_SS6_MGPIO21A_IN => GND_net_1, 
        SPI0_SS7_MGPIO22A_IN => GND_net_1, SPI1_SCK_IN => 
        GND_net_1, SPI1_SDI_MGPIO11A_IN => GND_net_1, 
        SPI1_SDO_MGPIO12A_IN => GND_net_1, SPI1_SS0_MGPIO13A_IN
         => GND_net_1, SPI1_SS1_MGPIO14A_IN => GND_net_1, 
        SPI1_SS2_MGPIO15A_IN => GND_net_1, SPI1_SS3_MGPIO16A_IN
         => GND_net_1, SPI1_SS4_MGPIO17A_IN => GND_net_1, 
        SPI1_SS5_MGPIO18A_IN => GND_net_1, SPI1_SS6_MGPIO23A_IN
         => GND_net_1, SPI1_SS7_MGPIO24A_IN => GND_net_1, 
        USBC_XCLK_IN => GND_net_1, USBD_DATA0_IN => GND_net_1, 
        USBD_DATA1_IN => GND_net_1, USBD_DATA2_IN => GND_net_1, 
        USBD_DATA3_IN => GND_net_1, USBD_DATA4_IN => GND_net_1, 
        USBD_DATA5_IN => GND_net_1, USBD_DATA6_IN => GND_net_1, 
        USBD_DATA7_MGPIO23B_IN => GND_net_1, USBD_DIR_IN => 
        GND_net_1, USBD_NXT_IN => GND_net_1, USBD_STP_IN => 
        GND_net_1, USBD_XCLK_IN => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => OPEN, DRAM_ADDR(15)
         => nc21, DRAM_ADDR(14) => nc237, DRAM_ADDR(13) => nc93, 
        DRAM_ADDR(12) => nc262, DRAM_ADDR(11) => nc69, 
        DRAM_ADDR(10) => nc206, DRAM_ADDR(9) => nc174, 
        DRAM_ADDR(8) => nc38, DRAM_ADDR(7) => nc113, DRAM_ADDR(6)
         => nc218, DRAM_ADDR(5) => nc106, DRAM_ADDR(4) => nc261, 
        DRAM_ADDR(3) => nc25, DRAM_ADDR(2) => nc1, DRAM_ADDR(1)
         => nc299, DRAM_ADDR(0) => nc37, DRAM_BA(2) => nc202, 
        DRAM_BA(1) => nc144, DRAM_BA(0) => nc153, DRAM_CASN => 
        OPEN, DRAM_CKE => OPEN, DRAM_CLK => OPEN, DRAM_CSN => 
        OPEN, DRAM_DM_RDQS_OUT(2) => nc46, DRAM_DM_RDQS_OUT(1)
         => nc258, DRAM_DM_RDQS_OUT(0) => nc71, DRAM_DQ_OUT(17)
         => nc124, DRAM_DQ_OUT(16) => nc81, DRAM_DQ_OUT(15) => 
        nc201, DRAM_DQ_OUT(14) => nc168, DRAM_DQ_OUT(13) => nc34, 
        DRAM_DQ_OUT(12) => nc28, DRAM_DQ_OUT(11) => nc115, 
        DRAM_DQ_OUT(10) => nc264, DRAM_DQ_OUT(9) => nc192, 
        DRAM_DQ_OUT(8) => nc319, DRAM_DQ_OUT(7) => nc134, 
        DRAM_DQ_OUT(6) => nc32, DRAM_DQ_OUT(5) => nc40, 
        DRAM_DQ_OUT(4) => nc297, DRAM_DQ_OUT(3) => nc99, 
        DRAM_DQ_OUT(2) => nc75, DRAM_DQ_OUT(1) => nc183, 
        DRAM_DQ_OUT(0) => nc288, DRAM_DQS_OUT(2) => nc85, 
        DRAM_DQS_OUT(1) => nc27, DRAM_DQS_OUT(0) => nc108, 
        DRAM_FIFO_WE_OUT(1) => nc16, DRAM_FIFO_WE_OUT(0) => nc155, 
        DRAM_ODT => OPEN, DRAM_RASN => OPEN, DRAM_RSTN => OPEN, 
        DRAM_WEN => OPEN, I2C0_SCL_USBC_DATA1_MGPIO31B_OUT => 
        OPEN, I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => OPEN, MGPIO0B_OUT => 
        OPEN, MGPIO10B_OUT => OPEN, MGPIO1B_OUT => OPEN, 
        MGPIO25A_OUT => OPEN, MGPIO26A_OUT => OPEN, MGPIO27A_OUT
         => OPEN, MGPIO28A_OUT => OPEN, MGPIO29A_OUT => OPEN, 
        MGPIO2B_OUT => OPEN, MGPIO30A_OUT => OPEN, MGPIO31A_OUT
         => OPEN, MGPIO3B_OUT => OPEN, MGPIO4B_OUT => OPEN, 
        MGPIO5B_OUT => OPEN, MGPIO6B_OUT => OPEN, MGPIO7B_OUT => 
        OPEN, MGPIO8B_OUT => OPEN, MGPIO9B_OUT => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT => OPEN, 
        MMUART0_DCD_MGPIO22B_OUT => OPEN, 
        MMUART0_DSR_MGPIO20B_OUT => OPEN, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => OPEN, 
        MMUART1_CTS_MGPIO13B_OUT => OPEN, 
        MMUART1_DCD_MGPIO16B_OUT => OPEN, 
        MMUART1_DSR_MGPIO14B_OUT => OPEN, 
        MMUART1_DTR_MGPIO12B_OUT => OPEN, MMUART1_RI_MGPIO15B_OUT
         => OPEN, MMUART1_RTS_MGPIO11B_OUT => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => OPEN, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => OPEN, 
        RGMII_RXD3_USBB_DATA4_OUT => OPEN, RGMII_TX_CLK_OUT => 
        OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => OPEN, 
        RGMII_TXD2_USBB_DATA5_OUT => OPEN, 
        RGMII_TXD3_USBB_DATA6_OUT => OPEN, SPI0_SCK_USBA_XCLK_OUT
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => OPEN, 
        SPI0_SS4_MGPIO19A_OUT => OPEN, SPI0_SS5_MGPIO20A_OUT => 
        OPEN, SPI0_SS6_MGPIO21A_OUT => OPEN, 
        SPI0_SS7_MGPIO22A_OUT => OPEN, SPI1_SCK_OUT => OPEN, 
        SPI1_SDI_MGPIO11A_OUT => OPEN, SPI1_SDO_MGPIO12A_OUT => 
        OPEN, SPI1_SS0_MGPIO13A_OUT => OPEN, 
        SPI1_SS1_MGPIO14A_OUT => OPEN, SPI1_SS2_MGPIO15A_OUT => 
        OPEN, SPI1_SS3_MGPIO16A_OUT => OPEN, 
        SPI1_SS4_MGPIO17A_OUT => OPEN, SPI1_SS5_MGPIO18A_OUT => 
        OPEN, SPI1_SS6_MGPIO23A_OUT => OPEN, 
        SPI1_SS7_MGPIO24A_OUT => OPEN, USBC_XCLK_OUT => OPEN, 
        USBD_DATA0_OUT => OPEN, USBD_DATA1_OUT => OPEN, 
        USBD_DATA2_OUT => OPEN, USBD_DATA3_OUT => OPEN, 
        USBD_DATA4_OUT => OPEN, USBD_DATA5_OUT => OPEN, 
        USBD_DATA6_OUT => OPEN, USBD_DATA7_MGPIO23B_OUT => OPEN, 
        USBD_DIR_OUT => OPEN, USBD_NXT_OUT => OPEN, USBD_STP_OUT
         => OPEN, USBD_XCLK_OUT => OPEN, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => OPEN, DM_OE(2) => nc51, 
        DM_OE(1) => nc301, DM_OE(0) => nc33, DRAM_DQ_OE(17) => 
        nc204, DRAM_DQ_OE(16) => nc173, DRAM_DQ_OE(15) => nc278, 
        DRAM_DQ_OE(14) => nc169, DRAM_DQ_OE(13) => nc78, 
        DRAM_DQ_OE(12) => nc263, DRAM_DQ_OE(11) => nc24, 
        DRAM_DQ_OE(10) => nc88, DRAM_DQ_OE(9) => nc111, 
        DRAM_DQ_OE(8) => nc55, DRAM_DQ_OE(7) => nc10, 
        DRAM_DQ_OE(6) => nc22, DRAM_DQ_OE(5) => nc210, 
        DRAM_DQ_OE(4) => nc185, DRAM_DQ_OE(3) => nc143, 
        DRAM_DQ_OE(2) => nc248, DRAM_DQ_OE(1) => nc77, 
        DRAM_DQ_OE(0) => nc6, DRAM_DQS_OE(2) => nc109, 
        DRAM_DQS_OE(1) => nc87, DRAM_DQS_OE(0) => nc123, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => OPEN, MGPIO0B_OE => 
        OPEN, MGPIO10B_OE => OPEN, MGPIO1B_OE => OPEN, 
        MGPIO25A_OE => OPEN, MGPIO26A_OE => OPEN, MGPIO27A_OE => 
        OPEN, MGPIO28A_OE => OPEN, MGPIO29A_OE => OPEN, 
        MGPIO2B_OE => OPEN, MGPIO30A_OE => OPEN, MGPIO31A_OE => 
        OPEN, MGPIO3B_OE => OPEN, MGPIO4B_OE => OPEN, MGPIO5B_OE
         => OPEN, MGPIO6B_OE => OPEN, MGPIO7B_OE => OPEN, 
        MGPIO8B_OE => OPEN, MGPIO9B_OE => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => OPEN, 
        MMUART0_DCD_MGPIO22B_OE => OPEN, MMUART0_DSR_MGPIO20B_OE
         => OPEN, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => OPEN, 
        MMUART1_CTS_MGPIO13B_OE => OPEN, MMUART1_DCD_MGPIO16B_OE
         => OPEN, MMUART1_DSR_MGPIO14B_OE => OPEN, 
        MMUART1_DTR_MGPIO12B_OE => OPEN, MMUART1_RI_MGPIO15B_OE
         => OPEN, MMUART1_RTS_MGPIO11B_OE => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => OPEN, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => OPEN, 
        RGMII_RXD3_USBB_DATA4_OE => OPEN, RGMII_TX_CLK_OE => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => OPEN, 
        RGMII_TXD2_USBB_DATA5_OE => OPEN, 
        RGMII_TXD3_USBB_DATA6_OE => OPEN, SPI0_SCK_USBA_XCLK_OE
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => OPEN, 
        SPI0_SS4_MGPIO19A_OE => OPEN, SPI0_SS5_MGPIO20A_OE => 
        OPEN, SPI0_SS6_MGPIO21A_OE => OPEN, SPI0_SS7_MGPIO22A_OE
         => OPEN, SPI1_SCK_OE => OPEN, SPI1_SDI_MGPIO11A_OE => 
        OPEN, SPI1_SDO_MGPIO12A_OE => OPEN, SPI1_SS0_MGPIO13A_OE
         => OPEN, SPI1_SS1_MGPIO14A_OE => OPEN, 
        SPI1_SS2_MGPIO15A_OE => OPEN, SPI1_SS3_MGPIO16A_OE => 
        OPEN, SPI1_SS4_MGPIO17A_OE => OPEN, SPI1_SS5_MGPIO18A_OE
         => OPEN, SPI1_SS6_MGPIO23A_OE => OPEN, 
        SPI1_SS7_MGPIO24A_OE => OPEN, USBC_XCLK_OE => OPEN, 
        USBD_DATA0_OE => OPEN, USBD_DATA1_OE => OPEN, 
        USBD_DATA2_OE => OPEN, USBD_DATA3_OE => OPEN, 
        USBD_DATA4_OE => OPEN, USBD_DATA5_OE => OPEN, 
        USBD_DATA6_OE => OPEN, USBD_DATA7_MGPIO23B_OE => OPEN, 
        USBD_DIR_OE => OPEN, USBD_NXT_OE => OPEN, USBD_STP_OE => 
        OPEN, USBD_XCLK_OE => OPEN);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    SPI_0_CLK_PAD : BIBUF
      port map(PAD => SPI_0_CLK, D => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, E => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, Y => 
        SPI_0_CLK_PAD_Y);
    
    MMUART_1_TXD_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, PAD
         => MMUART_1_TXD);
    
    MMUART_1_RXD_PAD : INBUF
      port map(PAD => MMUART_1_RXD, Y => MMUART_1_RXD_PAD_Y);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_CCC_0_FCCC is

    port( CertificationSystem_sb_0_FAB_CCC_GL0               : out   std_logic;
          FAB_CCC_LOCK                                       : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic
        );

end CertificationSystem_sb_CCC_0_FCCC;

architecture DEF_ARCH of CertificationSystem_sb_CCC_0_FCCC is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => 
        CertificationSystem_sb_0_FAB_CCC_GL0);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007FB8000045174000318C6318C1F18C61EC0404040400101",
         VCOFREQUENCY => 800.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => FAB_CCC_LOCK, 
        BUSY => OPEN, CLK0 => VCC_net_1, CLK1 => VCC_net_1, CLK2
         => VCC_net_1, CLK3 => VCC_net_1, NGMUX0_SEL => GND_net_1, 
        NGMUX1_SEL => GND_net_1, NGMUX2_SEL => GND_net_1, 
        NGMUX3_SEL => GND_net_1, NGMUX0_HOLD_N => VCC_net_1, 
        NGMUX1_HOLD_N => VCC_net_1, NGMUX2_HOLD_N => VCC_net_1, 
        NGMUX3_HOLD_N => VCC_net_1, NGMUX0_ARST_N => VCC_net_1, 
        NGMUX1_ARST_N => VCC_net_1, NGMUX2_ARST_N => VCC_net_1, 
        NGMUX3_ARST_N => VCC_net_1, PLL_BYPASS_N => VCC_net_1, 
        PLL_ARST_N => VCC_net_1, PLL_POWERDOWN_N => VCC_net_1, 
        GPD0_ARST_N => VCC_net_1, GPD1_ARST_N => VCC_net_1, 
        GPD2_ARST_N => VCC_net_1, GPD3_ARST_N => VCC_net_1, 
        PRESET_N => GND_net_1, PCLK => VCC_net_1, PSEL => 
        VCC_net_1, PENABLE => VCC_net_1, PWRITE => VCC_net_1, 
        PADDR(7) => VCC_net_1, PADDR(6) => VCC_net_1, PADDR(5)
         => VCC_net_1, PADDR(4) => VCC_net_1, PADDR(3) => 
        VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7) => VCC_net_1, 
        PWDATA(6) => VCC_net_1, PWDATA(5) => VCC_net_1, PWDATA(4)
         => VCC_net_1, PWDATA(3) => VCC_net_1, PWDATA(2) => 
        VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0) => VCC_net_1, 
        CLK0_PAD => GND_net_1, CLK1_PAD => GND_net_1, CLK2_PAD
         => GND_net_1, CLK3_PAD => GND_net_1, GL0 => GL0_net, GL1
         => OPEN, GL2 => OPEN, GL3 => OPEN, RCOSC_25_50MHZ => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        RCOSC_1MHZ => GND_net_1, XTLOSC => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity 
        CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8 is

    port( ram_rdata                            : out   std_logic_vector(31 downto 0);
          sram_wen_mem_m3                      : in    std_logic_vector(3 downto 2);
          sram_wen_mem                         : in    std_logic_vector(1 downto 0);
          ahbsram_addr                         : in    std_logic_vector(15 downto 2);
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          MSS_READY                            : in    std_logic;
          N_375_i_0                            : in    std_logic;
          N_38_i_0                             : in    std_logic;
          N_40_i_0                             : in    std_logic;
          N_42_i_0                             : in    std_logic;
          N_44_i_0                             : in    std_logic;
          N_46_i_0                             : in    std_logic;
          N_48_i_0                             : in    std_logic;
          N_50_i_0                             : in    std_logic;
          N_52_i_0                             : in    std_logic;
          N_54_i_0                             : in    std_logic;
          N_56_i_0                             : in    std_logic;
          N_58_i_0                             : in    std_logic;
          N_64_i_0                             : in    std_logic;
          N_66_i_0                             : in    std_logic;
          N_68_i_0                             : in    std_logic;
          N_70_i_0                             : in    std_logic;
          N_72_i_0                             : in    std_logic;
          N_74_i_0                             : in    std_logic;
          N_76_i_0                             : in    std_logic;
          N_78_i_0                             : in    std_logic;
          N_80_i_0                             : in    std_logic;
          N_82_i_0                             : in    std_logic;
          N_84_i_0                             : in    std_logic;
          N_86_i_0                             : in    std_logic;
          N_88_i_0                             : in    std_logic;
          N_90_i_0                             : in    std_logic;
          N_92_i_0                             : in    std_logic;
          N_94_i_0                             : in    std_logic;
          N_96_i_0                             : in    std_logic;
          N_98_i_0                             : in    std_logic;
          N_60_i_0                             : in    std_logic;
          N_62_i_0                             : in    std_logic;
          N_63_i_0                             : in    std_logic
        );

end CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8;

architecture DEF_ARCH of 
        CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal N_497, \readData_31_am_1_1[31]_net_1\, N_401, 
        \readData_31_am[31]_net_1\, N_273, N_177, N_977, 
        \readData_31_bm_1_1[31]_net_1\, N_881, 
        \readData_31_bm[31]_net_1\, N_753, N_657, N_496, 
        \readData_31_am_1_1[30]_net_1\, N_400, 
        \readData_31_am[30]_net_1\, N_272, N_176, N_976, 
        \readData_31_bm_1_1[30]_net_1\, N_880, 
        \readData_31_bm[30]_net_1\, N_752, N_656, N_495, 
        \readData_31_am_1_1[29]_net_1\, N_399, 
        \readData_31_am[29]_net_1\, N_271, N_175, N_975, 
        \readData_31_bm_1_1[29]_net_1\, N_879, 
        \readData_31_bm[29]_net_1\, N_751, N_655, N_494, 
        \readData_31_am_1_1[28]_net_1\, N_398, 
        \readData_31_am[28]_net_1\, N_270, N_174, N_974, 
        \readData_31_bm_1_1[28]_net_1\, N_878, 
        \readData_31_bm[28]_net_1\, N_750, N_654, N_493, 
        \readData_31_am_1_1[27]_net_1\, N_397, 
        \readData_31_am[27]_net_1\, N_269, N_173, N_973, 
        \readData_31_bm_1_1[27]_net_1\, N_877, 
        \readData_31_bm[27]_net_1\, N_749, N_653, N_492, 
        \readData_31_am_1_1[26]_net_1\, N_396, 
        \readData_31_am[26]_net_1\, N_268, N_172, N_972, 
        \readData_31_bm_1_1[26]_net_1\, N_876, 
        \readData_31_bm[26]_net_1\, N_748, N_652, N_491, 
        \readData_31_am_1_1[25]_net_1\, N_395, 
        \readData_31_am[25]_net_1\, N_267, N_171, N_971, 
        \readData_31_bm_1_1[25]_net_1\, N_875, 
        \readData_31_bm[25]_net_1\, N_747, N_651, N_490, 
        \readData_31_am_1_1[24]_net_1\, N_394, 
        \readData_31_am[24]_net_1\, N_266, N_170, N_970, 
        \readData_31_bm_1_1[24]_net_1\, N_874, 
        \readData_31_bm[24]_net_1\, N_746, N_650, N_489, 
        \readData_31_am_1_1[23]_net_1\, N_393, 
        \readData_31_am[23]_net_1\, N_265, N_169, N_969, 
        \readData_31_bm_1_1[23]_net_1\, N_873, 
        \readData_31_bm[23]_net_1\, N_745, N_649, N_488, 
        \readData_31_am_1_1[22]_net_1\, N_392, 
        \readData_31_am[22]_net_1\, N_264, N_168, N_968, 
        \readData_31_bm_1_1[22]_net_1\, N_872, 
        \readData_31_bm[22]_net_1\, N_744, N_648, N_487, 
        \readData_31_am_1_1[21]_net_1\, N_391, 
        \readData_31_am[21]_net_1\, N_263, N_167, N_967, 
        \readData_31_bm_1_1[21]_net_1\, N_871, 
        \readData_31_bm[21]_net_1\, N_743, N_647, N_486, 
        \readData_31_am_1_1[20]_net_1\, N_390, 
        \readData_31_am[20]_net_1\, N_262, N_166, N_966, 
        \readData_31_bm_1_1[20]_net_1\, N_870, 
        \readData_31_bm[20]_net_1\, N_742, N_646, N_485, 
        \readData_31_am_1_1[19]_net_1\, N_389, 
        \readData_31_am[19]_net_1\, N_261, N_165, N_965, 
        \readData_31_bm_1_1[19]_net_1\, N_869, 
        \readData_31_bm[19]_net_1\, N_741, N_645, N_484, 
        \readData_31_am_1_1[18]_net_1\, N_388, 
        \readData_31_am[18]_net_1\, N_260, N_164, N_964, 
        \readData_31_bm_1_1[18]_net_1\, N_868, 
        \readData_31_bm[18]_net_1\, N_740, N_644, N_483, 
        \readData_31_am_1_1[17]_net_1\, N_387, 
        \readData_31_am[17]_net_1\, N_259, N_163, N_963, 
        \readData_31_bm_1_1[17]_net_1\, N_867, 
        \readData_31_bm[17]_net_1\, N_739, N_643, N_482, 
        \readData_31_am_1_1[16]_net_1\, N_386, 
        \readData_31_am[16]_net_1\, N_258, N_162, N_962, 
        \readData_31_bm_1_1[16]_net_1\, N_866, 
        \readData_31_bm[16]_net_1\, N_738, N_642, N_481, 
        \readData_31_am_1_1[15]_net_1\, N_385, 
        \readData_31_am[15]_net_1\, N_257, N_161, N_961, 
        \readData_31_bm_1_1[15]_net_1\, N_865, 
        \readData_31_bm[15]_net_1\, N_737, N_641, N_480, 
        \readData_31_am_1_1[14]_net_1\, N_384, 
        \readData_31_am[14]_net_1\, N_256, N_160, N_960, 
        \readData_31_bm_1_1[14]_net_1\, N_864, 
        \readData_31_bm[14]_net_1\, N_736, N_640, N_479, 
        \readData_31_am_1_1[13]_net_1\, N_383, 
        \readData_31_am[13]_net_1\, N_255, N_159, N_959, 
        \readData_31_bm_1_1[13]_net_1\, N_863, 
        \readData_31_bm[13]_net_1\, N_735, N_639, N_478, 
        \readData_31_am_1_1[12]_net_1\, N_382, 
        \readData_31_am[12]_net_1\, N_254, N_158, N_958, 
        \readData_31_bm_1_1[12]_net_1\, N_862, 
        \readData_31_bm[12]_net_1\, N_734, N_638, N_477, 
        \readData_31_am_1_1[11]_net_1\, N_381, 
        \readData_31_am[11]_net_1\, N_253, N_157, N_957, 
        \readData_31_bm_1_1[11]_net_1\, N_861, 
        \readData_31_bm[11]_net_1\, N_733, N_637, N_476, 
        \readData_31_am_1_1[10]_net_1\, N_380, 
        \readData_31_am[10]_net_1\, N_252, N_156, N_956, 
        \readData_31_bm_1_1[10]_net_1\, N_860, 
        \readData_31_bm[10]_net_1\, N_732, N_636, N_475, 
        \readData_31_am_1_1[9]_net_1\, N_379, 
        \readData_31_am[9]_net_1\, N_251, N_155, N_955, 
        \readData_31_bm_1_1[9]_net_1\, N_859, 
        \readData_31_bm[9]_net_1\, N_731, N_635, N_474, 
        \readData_31_am_1_1[8]_net_1\, N_378, 
        \readData_31_am[8]_net_1\, N_250, N_154, N_954, 
        \readData_31_bm_1_1[8]_net_1\, N_858, 
        \readData_31_bm[8]_net_1\, N_730, N_634, N_473, 
        \readData_31_am_1_1[7]_net_1\, N_377, 
        \readData_31_am[7]_net_1\, N_249, N_153, N_953, 
        \readData_31_bm_1_1[7]_net_1\, N_857, 
        \readData_31_bm[7]_net_1\, N_729, N_633, N_472, 
        \readData_31_am_1_1[6]_net_1\, N_376, 
        \readData_31_am[6]_net_1\, N_248, N_152, N_952, 
        \readData_31_bm_1_1[6]_net_1\, N_856, 
        \readData_31_bm[6]_net_1\, N_728, N_632, N_471, 
        \readData_31_am_1_1[5]_net_1\, N_375, 
        \readData_31_am[5]_net_1\, N_247, N_151, N_951, 
        \readData_31_bm_1_1[5]_net_1\, N_855, 
        \readData_31_bm[5]_net_1\, N_727, N_631, N_470, 
        \readData_31_am_1_1[4]_net_1\, N_374, 
        \readData_31_am[4]_net_1\, N_246, N_150, N_950, 
        \readData_31_bm_1_1[4]_net_1\, N_854, 
        \readData_31_bm[4]_net_1\, N_726, N_630, N_469, 
        \readData_31_am_1_1[3]_net_1\, N_373, 
        \readData_31_am[3]_net_1\, N_245, N_149, N_949, 
        \readData_31_bm_1_1[3]_net_1\, N_853, 
        \readData_31_bm[3]_net_1\, N_725, N_629, N_468, 
        \readData_31_am_1_1[2]_net_1\, N_372, 
        \readData_31_am[2]_net_1\, N_244, N_148, N_948, 
        \readData_31_bm_1_1[2]_net_1\, N_852, 
        \readData_31_bm[2]_net_1\, N_724, N_628, N_467, 
        \readData_31_am_1_1[1]_net_1\, N_371, 
        \readData_31_am[1]_net_1\, N_243, N_147, N_947, 
        \readData_31_bm_1_1[1]_net_1\, N_851, 
        \readData_31_bm[1]_net_1\, N_723, N_627, N_466, 
        \readData_31_am_1_1[0]_net_1\, N_370, 
        \readData_31_am[0]_net_1\, N_242, N_146, N_946, 
        \readData_31_bm_1_1[0]_net_1\, N_850, 
        \readData_31_bm[0]_net_1\, N_722, N_626, \readData31[29]\, 
        \readData_28_1_1[26]\, \readData15[29]\, \readData23[29]\, 
        \readData7[29]\, \readData31[24]\, \readData_28_1_1[22]\, 
        \readData15[24]\, \readData23[24]\, \readData7[24]\, 
        \readData27[7]\, \readData_25_1_1[7]\, \readData11[7]\, 
        \readData19[7]\, \readData3[7]\, \readData31[25]\, 
        \readData_28_1_1[23]\, \readData15[25]\, \readData23[25]\, 
        \readData7[25]\, \readData31[30]\, \readData_28_1_1[27]\, 
        \readData15[30]\, \readData23[30]\, \readData7[30]\, 
        \readData31[19]\, \readData_28_1_1[17]\, \readData15[19]\, 
        \readData23[19]\, \readData7[19]\, \readData31[27]\, 
        \readData_28_1_1[24]\, \readData15[27]\, \readData23[27]\, 
        \readData7[27]\, \readData31[21]\, \readData_28_1_1[19]\, 
        \readData15[21]\, \readData23[21]\, \readData7[21]\, 
        \readData31[32]\, \readData_28_1_1[29]\, \readData15[32]\, 
        \readData23[32]\, \readData7[32]\, \readData27[2]\, 
        \readData_25_1_1[2]\, \readData11[2]\, \readData19[2]\, 
        \readData3[2]\, \readData31[6]\, \readData_28_1_1[6]\, 
        \readData15[6]\, \readData23[6]\, \readData7[6]\, 
        \readData27[1]\, \readData_25_1_1[1]\, \readData11[1]\, 
        \readData19[1]\, \readData3[1]\, \readData31[31]\, 
        \readData_28_1_1[28]\, \readData15[31]\, \readData23[31]\, 
        \readData7[31]\, \readData29[13]\, \readData_21_1_1[12]\, 
        \readData13[13]\, \readData21[13]\, \readData5[13]\, 
        \readData27[0]\, \readData_25_1_1[0]\, \readData11[0]\, 
        \readData19[0]\, \readData3[0]\, \readData27[5]\, 
        \readData_25_1_1[5]\, \readData11[5]\, \readData19[5]\, 
        \readData3[5]\, \readData30[20]\, \readData_13_1_1[18]\, 
        \readData14[20]\, \readData22[20]\, \readData6[20]\, 
        \readData27[6]\, \readData_25_1_1[6]\, \readData11[6]\, 
        \readData19[6]\, \readData3[6]\, \readData31[13]\, 
        \readData_28_1_1[12]\, \readData15[13]\, \readData23[13]\, 
        \readData7[13]\, \readData30[16]\, \readData_13_1_1[15]\, 
        \readData14[16]\, \readData22[16]\, \readData6[16]\, 
        \readData31[20]\, \readData_28_1_1[18]\, \readData15[20]\, 
        \readData23[20]\, \readData7[20]\, \readData30[13]\, 
        \readData_13_1_1[12]\, \readData14[13]\, \readData22[13]\, 
        \readData6[13]\, \readData31[16]\, \readData_28_1_1[15]\, 
        \readData15[16]\, \readData23[16]\, \readData7[16]\, 
        \readData29[2]\, \readData_21_1_1[2]\, \readData13[2]\, 
        \readData21[2]\, \readData5[2]\, \readData31[14]\, 
        \readData_28_1_1[13]\, \readData15[14]\, \readData23[14]\, 
        \readData7[14]\, \readData29[10]\, \readData_21_1_1[9]\, 
        \readData13[10]\, \readData21[10]\, \readData5[10]\, 
        \readData30[11]\, \readData_13_1_1[10]\, \readData14[11]\, 
        \readData22[11]\, \readData6[11]\, \readData30[19]\, 
        \readData_13_1_1[17]\, \readData14[19]\, \readData22[19]\, 
        \readData6[19]\, \readData30[18]\, \readData_13_1_1[16]\, 
        \readData14[18]\, \readData22[18]\, \readData6[18]\, 
        \readData31[9]\, \readData_28_1_1[8]\, \readData15[9]\, 
        \readData23[9]\, \readData7[9]\, \readData31[7]\, 
        \readData_28_1_1[7]\, \readData15[7]\, \readData23[7]\, 
        \readData7[7]\, \readData31[5]\, \readData_28_1_1[5]\, 
        \readData15[5]\, \readData23[5]\, \readData7[5]\, 
        \readData30[1]\, \readData_13_1_1[1]\, \readData14[1]\, 
        \readData22[1]\, \readData6[1]\, \readData31[3]\, 
        \readData_28_1_1[3]\, \readData15[3]\, \readData23[3]\, 
        \readData7[3]\, \readData31[2]\, \readData_28_1_1[2]\, 
        \readData15[2]\, \readData23[2]\, \readData7[2]\, 
        \readData31[1]\, \readData_28_1_1[1]\, \readData15[1]\, 
        \readData23[1]\, \readData7[1]\, \readData29[9]\, 
        \readData_21_1_1[8]\, \readData13[9]\, \readData21[9]\, 
        \readData5[9]\, \readData29[6]\, \readData_21_1_1[6]\, 
        \readData13[6]\, \readData21[6]\, \readData5[6]\, 
        \readData27[11]\, \readData_25_1_1[10]\, \readData11[11]\, 
        \readData19[11]\, \readData3[11]\, \readData27[10]\, 
        \readData_25_1_1[9]\, \readData11[10]\, \readData19[10]\, 
        \readData3[10]\, \readData28[12]\, \readData_6_1_1[11]\, 
        \readData12[12]\, \readData20[12]\, \readData4[12]\, 
        \readData29[14]\, \readData_21_1_1[13]\, \readData13[14]\, 
        \readData21[14]\, \readData5[14]\, \readData31[34]\, 
        \readData_28_1_1[31]\, \readData15[34]\, \readData23[34]\, 
        \readData7[34]\, \readData31[33]\, \readData_28_1_1[30]\, 
        \readData15[33]\, \readData23[33]\, \readData7[33]\, 
        \readData29[7]\, \readData_21_1_1[7]\, \readData13[7]\, 
        \readData21[7]\, \readData5[7]\, \readData29[1]\, 
        \readData_21_1_1[1]\, \readData13[1]\, \readData21[1]\, 
        \readData5[1]\, \readData29[0]\, \readData_21_1_1[0]\, 
        \readData13[0]\, \readData21[0]\, \readData5[0]\, 
        \readData30[12]\, \readData_13_1_1[11]\, \readData14[12]\, 
        \readData22[12]\, \readData6[12]\, \readData31[15]\, 
        \readData_28_1_1[14]\, \readData15[15]\, \readData23[15]\, 
        \readData7[15]\, \readData28[2]\, \readData_6_1_1[2]\, 
        \readData12[2]\, \readData20[2]\, \readData4[2]\, 
        \readData31[10]\, \readData_28_1_1[9]\, \readData15[10]\, 
        \readData23[10]\, \readData7[10]\, \readData25[5]\, 
        \readData_18_1_1[5]\, \readData9[5]\, \readData17[5]\, 
        \readData1[5]\, \readData30[3]\, \readData_13_1_1[3]\, 
        \readData14[3]\, \readData22[3]\, \readData6[3]\, 
        \readData27[24]\, \readData_25_1_1[22]\, \readData11[24]\, 
        \readData19[24]\, \readData3[24]\, \readData27[23]\, 
        \readData_25_1_1[21]\, \readData11[23]\, \readData19[23]\, 
        \readData3[23]\, \readData31[4]\, \readData_28_1_1[4]\, 
        \readData15[4]\, \readData23[4]\, \readData7[4]\, 
        \readData28[19]\, \readData_6_1_1[17]\, \readData12[19]\, 
        \readData20[19]\, \readData4[19]\, \readData28[18]\, 
        \readData_6_1_1[16]\, \readData12[18]\, \readData20[18]\, 
        \readData4[18]\, \readData28[16]\, \readData_6_1_1[15]\, 
        \readData12[16]\, \readData20[16]\, \readData4[16]\, 
        \readData27[15]\, \readData_25_1_1[14]\, \readData11[15]\, 
        \readData19[15]\, \readData3[15]\, \readData28[13]\, 
        \readData_6_1_1[12]\, \readData12[13]\, \readData20[13]\, 
        \readData4[13]\, \readData30[34]\, \readData_13_1_1[31]\, 
        \readData14[34]\, \readData22[34]\, \readData6[34]\, 
        \readData28[10]\, \readData_6_1_1[9]\, \readData12[10]\, 
        \readData20[10]\, \readData4[10]\, \readData28[9]\, 
        \readData_6_1_1[8]\, \readData12[9]\, \readData20[9]\, 
        \readData4[9]\, \readData30[30]\, \readData_13_1_1[27]\, 
        \readData14[30]\, \readData22[30]\, \readData6[30]\, 
        \readData30[29]\, \readData_13_1_1[26]\, \readData14[29]\, 
        \readData22[29]\, \readData6[29]\, \readData28[5]\, 
        \readData_6_1_1[5]\, \readData12[5]\, \readData20[5]\, 
        \readData4[5]\, \readData28[4]\, \readData_6_1_1[4]\, 
        \readData12[4]\, \readData20[4]\, \readData4[4]\, 
        \readData28[3]\, \readData_6_1_1[3]\, \readData12[3]\, 
        \readData20[3]\, \readData4[3]\, \readData31[28]\, 
        \readData_28_1_1[25]\, \readData15[28]\, \readData23[28]\, 
        \readData7[28]\, \readData28[0]\, \readData_6_1_1[0]\, 
        \readData12[0]\, \readData20[0]\, \readData4[0]\, 
        \readData31[23]\, \readData_28_1_1[21]\, \readData15[23]\, 
        \readData23[23]\, \readData7[23]\, \readData31[22]\, 
        \readData_28_1_1[20]\, \readData15[22]\, \readData23[22]\, 
        \readData7[22]\, \readData30[14]\, \readData_13_1_1[13]\, 
        \readData14[14]\, \readData22[14]\, \readData6[14]\, 
        \readData30[9]\, \readData_13_1_1[8]\, \readData14[9]\, 
        \readData22[9]\, \readData6[9]\, \readData31[12]\, 
        \readData_28_1_1[11]\, \readData15[12]\, \readData23[12]\, 
        \readData7[12]\, \readData30[4]\, \readData_13_1_1[4]\, 
        \readData14[4]\, \readData22[4]\, \readData6[4]\, 
        \readData27[27]\, \readData_25_1_1[24]\, \readData11[27]\, 
        \readData19[27]\, \readData3[27]\, \readData25[4]\, 
        \readData_18_1_1[4]\, \readData9[4]\, \readData17[4]\, 
        \readData1[4]\, \readData30[2]\, \readData_13_1_1[2]\, 
        \readData14[2]\, \readData22[2]\, \readData6[2]\, 
        \readData25[1]\, \readData_18_1_1[1]\, \readData9[1]\, 
        \readData17[1]\, \readData1[1]\, \readData25[0]\, 
        \readData_18_1_1[0]\, \readData9[0]\, \readData17[0]\, 
        \readData1[0]\, \readData31[0]\, \readData_28_1_1[0]\, 
        \readData15[0]\, \readData23[0]\, \readData7[0]\, 
        \readData29[24]\, \readData_21_1_1[22]\, \readData13[24]\, 
        \readData21[24]\, \readData5[24]\, \readData29[23]\, 
        \readData_21_1_1[21]\, \readData13[23]\, \readData21[23]\, 
        \readData5[23]\, \readData29[21]\, \readData_21_1_1[19]\, 
        \readData13[21]\, \readData21[21]\, \readData5[21]\, 
        \readData30[33]\, \readData_13_1_1[30]\, \readData14[33]\, 
        \readData22[33]\, \readData6[33]\, \readData30[32]\, 
        \readData_13_1_1[29]\, \readData14[32]\, \readData22[32]\, 
        \readData6[32]\, \readData27[9]\, \readData_25_1_1[8]\, 
        \readData11[9]\, \readData19[9]\, \readData3[9]\, 
        \readData29[16]\, \readData_21_1_1[15]\, \readData13[16]\, 
        \readData21[16]\, \readData5[16]\, \readData29[15]\, 
        \readData_21_1_1[14]\, \readData13[15]\, \readData21[15]\, 
        \readData5[15]\, \readData27[4]\, \readData_25_1_1[4]\, 
        \readData11[4]\, \readData19[4]\, \readData3[4]\, 
        \readData27[3]\, \readData_25_1_1[3]\, \readData11[3]\, 
        \readData19[3]\, \readData3[3]\, \readData30[24]\, 
        \readData_13_1_1[22]\, \readData14[24]\, \readData22[24]\, 
        \readData6[24]\, \readData30[23]\, \readData_13_1_1[21]\, 
        \readData14[23]\, \readData22[23]\, \readData6[23]\, 
        \readData29[5]\, \readData_21_1_1[5]\, \readData13[5]\, 
        \readData21[5]\, \readData5[5]\, \readData30[15]\, 
        \readData_13_1_1[14]\, \readData14[15]\, \readData22[15]\, 
        \readData6[15]\, \readData25[11]\, \readData_18_1_1[10]\, 
        \readData9[11]\, \readData17[11]\, \readData1[11]\, 
        \readData30[7]\, \readData_13_1_1[7]\, \readData14[7]\, 
        \readData22[7]\, \readData6[7]\, \readData31[11]\, 
        \readData_28_1_1[10]\, \readData15[11]\, \readData23[11]\, 
        \readData7[11]\, \readData30[5]\, \readData_13_1_1[5]\, 
        \readData14[5]\, \readData22[5]\, \readData6[5]\, 
        \readData29[34]\, \readData_21_1_1[31]\, \readData13[34]\, 
        \readData21[34]\, \readData5[34]\, \readData29[33]\, 
        \readData_21_1_1[30]\, \readData13[33]\, \readData21[33]\, 
        \readData5[33]\, \readData29[32]\, \readData_21_1_1[29]\, 
        \readData13[32]\, \readData21[32]\, \readData5[32]\, 
        \readData27[20]\, \readData_25_1_1[18]\, \readData11[20]\, 
        \readData19[20]\, \readData3[20]\, \readData28[20]\, 
        \readData_6_1_1[18]\, \readData12[20]\, \readData20[20]\, 
        \readData4[20]\, \readData27[18]\, \readData_25_1_1[16]\, 
        \readData11[18]\, \readData19[18]\, \readData3[18]\, 
        \readData27[16]\, \readData_25_1_1[15]\, \readData11[16]\, 
        \readData19[16]\, \readData3[16]\, \readData27[12]\, 
        \readData_25_1_1[11]\, \readData11[12]\, \readData19[12]\, 
        \readData3[12]\, \readData29[20]\, \readData_21_1_1[18]\, 
        \readData13[20]\, \readData21[20]\, \readData5[20]\, 
        \readData29[18]\, \readData_21_1_1[16]\, \readData13[18]\, 
        \readData21[18]\, \readData5[18]\, \readData25[33]\, 
        \readData_18_1_1[30]\, \readData9[33]\, \readData17[33]\, 
        \readData1[33]\, \readData30[28]\, \readData_13_1_1[25]\, 
        \readData14[28]\, \readData22[28]\, \readData6[28]\, 
        \readData26[0]\, \readData_10_1_1[0]\, \readData10[0]\, 
        \readData18[0]\, \readData2[0]\, \readData29[12]\, 
        \readData_21_1_1[11]\, \readData13[12]\, \readData21[12]\, 
        \readData5[12]\, \readData29[11]\, \readData_21_1_1[10]\, 
        \readData13[11]\, \readData21[11]\, \readData5[11]\, 
        \readData30[22]\, \readData_13_1_1[20]\, \readData14[22]\, 
        \readData22[22]\, \readData6[22]\, \readData29[4]\, 
        \readData_21_1_1[4]\, \readData13[4]\, \readData21[4]\, 
        \readData5[4]\, \readData31[18]\, \readData_28_1_1[16]\, 
        \readData15[18]\, \readData23[18]\, \readData7[18]\, 
        \readData30[10]\, \readData_13_1_1[9]\, \readData14[10]\, 
        \readData22[10]\, \readData6[10]\, \readData27[32]\, 
        \readData_25_1_1[29]\, \readData11[32]\, \readData19[32]\, 
        \readData3[32]\, \readData25[10]\, \readData_18_1_1[9]\, 
        \readData9[10]\, \readData17[10]\, \readData1[10]\, 
        \readData25[6]\, \readData_18_1_1[6]\, \readData9[6]\, 
        \readData17[6]\, \readData1[6]\, \readData28[29]\, 
        \readData_6_1_1[26]\, \readData12[29]\, \readData20[29]\, 
        \readData4[29]\, \readData29[31]\, \readData_21_1_1[28]\, 
        \readData13[31]\, \readData21[31]\, \readData5[31]\, 
        \readData29[30]\, \readData_21_1_1[27]\, \readData13[30]\, 
        \readData21[30]\, \readData5[30]\, \readData29[28]\, 
        \readData_21_1_1[25]\, \readData13[28]\, \readData21[28]\, 
        \readData5[28]\, \readData28[15]\, \readData_6_1_1[14]\, 
        \readData12[15]\, \readData20[15]\, \readData4[15]\, 
        \readData24[31]\, \readData_3_1_1[28]\, \readData8[31]\, 
        \readData16[31]\, \readData0[31]\, \readData28[11]\, 
        \readData_6_1_1[10]\, \readData12[11]\, \readData20[11]\, 
        \readData4[11]\, \readData26[1]\, \readData_10_1_1[1]\, 
        \readData10[1]\, \readData18[1]\, \readData2[1]\, 
        \readData28[7]\, \readData_6_1_1[7]\, \readData12[7]\, 
        \readData20[7]\, \readData4[7]\, \readData25[29]\, 
        \readData_18_1_1[26]\, \readData9[29]\, \readData17[29]\, 
        \readData1[29]\, \readData30[27]\, \readData_13_1_1[24]\, 
        \readData14[27]\, \readData22[27]\, \readData6[27]\, 
        \readData30[21]\, \readData_13_1_1[19]\, \readData14[21]\, 
        \readData22[21]\, \readData6[21]\, \readData25[24]\, 
        \readData_18_1_1[22]\, \readData9[24]\, \readData17[24]\, 
        \readData1[24]\, \readData25[22]\, \readData_18_1_1[20]\, 
        \readData9[22]\, \readData17[22]\, \readData1[22]\, 
        \readData25[15]\, \readData_18_1_1[14]\, \readData9[15]\, 
        \readData17[15]\, \readData1[15]\, \readData25[7]\, 
        \readData_18_1_1[7]\, \readData9[7]\, \readData17[7]\, 
        \readData1[7]\, \readData30[6]\, \readData_13_1_1[6]\, 
        \readData14[6]\, \readData22[6]\, \readData6[6]\, 
        \readData27[28]\, \readData_25_1_1[25]\, \readData11[28]\, 
        \readData19[28]\, \readData3[28]\, \readData28[30]\, 
        \readData_6_1_1[27]\, \readData12[30]\, \readData20[30]\, 
        \readData4[30]\, \readData28[28]\, \readData_6_1_1[25]\, 
        \readData12[28]\, \readData20[28]\, \readData4[28]\, 
        \readData30[0]\, \readData_13_1_1[0]\, \readData14[0]\, 
        \readData22[0]\, \readData6[0]\, \readData28[23]\, 
        \readData_6_1_1[21]\, \readData12[23]\, \readData20[23]\, 
        \readData4[23]\, \readData29[27]\, \readData_21_1_1[24]\, 
        \readData13[27]\, \readData21[27]\, \readData5[27]\, 
        \readData24[33]\, \readData_3_1_1[30]\, \readData8[33]\, 
        \readData16[33]\, \readData0[33]\, \readData28[14]\, 
        \readData_6_1_1[13]\, \readData12[14]\, \readData20[14]\, 
        \readData4[14]\, \readData25[34]\, \readData_18_1_1[31]\, 
        \readData9[34]\, \readData17[34]\, \readData1[34]\, 
        \readData25[32]\, \readData_18_1_1[29]\, \readData9[32]\, 
        \readData17[32]\, \readData1[32]\, \readData24[25]\, 
        \readData_3_1_1[23]\, \readData8[25]\, \readData16[25]\, 
        \readData0[25]\, \readData28[6]\, \readData_6_1_1[6]\, 
        \readData12[6]\, \readData20[6]\, \readData4[6]\, 
        \readData24[23]\, \readData_3_1_1[21]\, \readData8[23]\, 
        \readData16[23]\, \readData0[23]\, \readData30[25]\, 
        \readData_13_1_1[23]\, \readData14[25]\, \readData22[25]\, 
        \readData6[25]\, \readData28[1]\, \readData_6_1_1[1]\, 
        \readData12[1]\, \readData20[1]\, \readData4[1]\, 
        \readData25[23]\, \readData_18_1_1[21]\, \readData9[23]\, 
        \readData17[23]\, \readData1[23]\, \readData29[3]\, 
        \readData_21_1_1[3]\, \readData13[3]\, \readData21[3]\, 
        \readData5[3]\, \readData25[20]\, \readData_18_1_1[18]\, 
        \readData9[20]\, \readData17[20]\, \readData1[20]\, 
        \readData24[10]\, \readData_3_1_1[9]\, \readData8[10]\, 
        \readData16[10]\, \readData0[10]\, \readData25[12]\, 
        \readData_18_1_1[11]\, \readData9[12]\, \readData17[12]\, 
        \readData1[12]\, \readData28[34]\, \readData_6_1_1[31]\, 
        \readData12[34]\, \readData20[34]\, \readData4[34]\, 
        \readData28[33]\, \readData_6_1_1[30]\, \readData12[33]\, 
        \readData20[33]\, \readData4[33]\, \readData25[9]\, 
        \readData_18_1_1[8]\, \readData9[9]\, \readData17[9]\, 
        \readData1[9]\, \readData27[30]\, \readData_25_1_1[27]\, 
        \readData11[30]\, \readData19[30]\, \readData3[30]\, 
        \readData24[1]\, \readData_3_1_1[1]\, \readData8[1]\, 
        \readData16[1]\, \readData0[1]\, \readData28[27]\, 
        \readData_6_1_1[24]\, \readData12[27]\, \readData20[27]\, 
        \readData4[27]\, \readData25[2]\, \readData_18_1_1[2]\, 
        \readData9[2]\, \readData17[2]\, \readData1[2]\, 
        \readData28[22]\, \readData_6_1_1[20]\, \readData12[22]\, 
        \readData20[22]\, \readData4[22]\, \readData27[19]\, 
        \readData_25_1_1[17]\, \readData11[19]\, \readData19[19]\, 
        \readData3[19]\, \readData29[25]\, \readData_21_1_1[23]\, 
        \readData13[25]\, \readData21[25]\, \readData5[25]\, 
        \readData27[14]\, \readData_25_1_1[13]\, \readData11[14]\, 
        \readData19[14]\, \readData3[14]\, \readData27[13]\, 
        \readData_25_1_1[12]\, \readData11[13]\, \readData19[13]\, 
        \readData3[13]\, \readData24[28]\, \readData_3_1_1[25]\, 
        \readData8[28]\, \readData16[28]\, \readData0[28]\, 
        \readData30[31]\, \readData_13_1_1[28]\, \readData14[31]\, 
        \readData22[31]\, \readData6[31]\, \readData25[30]\, 
        \readData_18_1_1[27]\, \readData9[30]\, \readData17[30]\, 
        \readData1[30]\, \readData25[28]\, \readData_18_1_1[25]\, 
        \readData9[28]\, \readData17[28]\, \readData1[28]\, 
        \readData24[20]\, \readData_3_1_1[18]\, \readData8[20]\, 
        \readData16[20]\, \readData0[20]\, \readData24[19]\, 
        \readData_3_1_1[17]\, \readData8[19]\, \readData16[19]\, 
        \readData0[19]\, \readData24[16]\, \readData_3_1_1[15]\, 
        \readData8[16]\, \readData16[16]\, \readData0[16]\, 
        \readData25[19]\, \readData_18_1_1[17]\, \readData9[19]\, 
        \readData17[19]\, \readData1[19]\, \readData25[16]\, 
        \readData_18_1_1[15]\, \readData9[16]\, \readData17[16]\, 
        \readData1[16]\, \readData24[11]\, \readData_3_1_1[10]\, 
        \readData8[11]\, \readData16[11]\, \readData0[11]\, 
        \readData26[32]\, \readData_10_1_1[29]\, \readData10[32]\, 
        \readData18[32]\, \readData2[32]\, \readData26[31]\, 
        \readData_10_1_1[28]\, \readData10[31]\, \readData18[31]\, 
        \readData2[31]\, \readData27[33]\, \readData_25_1_1[30]\, 
        \readData11[33]\, \readData19[33]\, \readData3[33]\, 
        \readData24[6]\, \readData_3_1_1[6]\, \readData8[6]\, 
        \readData16[6]\, \readData0[6]\, \readData28[32]\, 
        \readData_6_1_1[29]\, \readData12[32]\, \readData20[32]\, 
        \readData4[32]\, \readData27[29]\, \readData_25_1_1[26]\, 
        \readData11[29]\, \readData19[29]\, \readData3[29]\, 
        \readData26[25]\, \readData_10_1_1[23]\, \readData10[25]\, 
        \readData18[25]\, \readData2[25]\, \readData24[2]\, 
        \readData_3_1_1[2]\, \readData8[2]\, \readData16[2]\, 
        \readData0[2]\, \readData24[0]\, \readData_3_1_1[0]\, 
        \readData8[0]\, \readData16[0]\, \readData0[0]\, 
        \readData25[3]\, \readData_18_1_1[3]\, \readData9[3]\, 
        \readData17[3]\, \readData1[3]\, \readData28[21]\, 
        \readData_6_1_1[19]\, \readData12[21]\, \readData20[21]\, 
        \readData4[21]\, \readData29[29]\, \readData_21_1_1[26]\, 
        \readData13[29]\, \readData21[29]\, \readData5[29]\, 
        \readData26[14]\, \readData_10_1_1[13]\, \readData10[14]\, 
        \readData18[14]\, \readData2[14]\, \readData26[13]\, 
        \readData_10_1_1[12]\, \readData10[13]\, \readData18[13]\, 
        \readData2[13]\, \readData24[32]\, \readData_3_1_1[29]\, 
        \readData8[32]\, \readData16[32]\, \readData0[32]\, 
        \readData26[7]\, \readData_10_1_1[7]\, \readData10[7]\, 
        \readData18[7]\, \readData2[7]\, \readData24[24]\, 
        \readData_3_1_1[22]\, \readData8[24]\, \readData16[24]\, 
        \readData0[24]\, \readData24[15]\, \readData_3_1_1[14]\, 
        \readData8[15]\, \readData16[15]\, \readData0[15]\, 
        \readData24[14]\, \readData_3_1_1[13]\, \readData8[14]\, 
        \readData16[14]\, \readData0[14]\, \readData25[18]\, 
        \readData_18_1_1[16]\, \readData9[18]\, \readData17[18]\, 
        \readData1[18]\, \readData24[9]\, \readData_3_1_1[8]\, 
        \readData8[9]\, \readData16[9]\, \readData0[9]\, 
        \readData27[34]\, \readData_25_1_1[31]\, \readData11[34]\, 
        \readData19[34]\, \readData3[34]\, \readData24[5]\, 
        \readData_3_1_1[5]\, \readData8[5]\, \readData16[5]\, 
        \readData0[5]\, \readData26[22]\, \readData_10_1_1[20]\, 
        \readData10[22]\, \readData18[22]\, \readData2[22]\, 
        \readData27[25]\, \readData_25_1_1[23]\, \readData11[25]\, 
        \readData19[25]\, \readData3[25]\, \readData26[19]\, 
        \readData_10_1_1[17]\, \readData10[19]\, \readData18[19]\, 
        \readData2[19]\, \readData27[22]\, \readData_25_1_1[20]\, 
        \readData11[22]\, \readData19[22]\, \readData3[22]\, 
        \readData27[21]\, \readData_25_1_1[19]\, \readData11[21]\, 
        \readData19[21]\, \readData3[21]\, \readData28[24]\, 
        \readData_6_1_1[22]\, \readData12[24]\, \readData20[24]\, 
        \readData4[24]\, \readData26[11]\, \readData_10_1_1[10]\, 
        \readData10[11]\, \readData18[11]\, \readData2[11]\, 
        \readData26[10]\, \readData_10_1_1[9]\, \readData10[10]\, 
        \readData18[10]\, \readData2[10]\, \readData29[22]\, 
        \readData_21_1_1[20]\, \readData13[22]\, \readData21[22]\, 
        \readData5[22]\, \readData26[6]\, \readData_10_1_1[6]\, 
        \readData10[6]\, \readData18[6]\, \readData2[6]\, 
        \readData24[29]\, \readData_3_1_1[26]\, \readData8[29]\, 
        \readData16[29]\, \readData0[29]\, \readData26[4]\, 
        \readData_10_1_1[4]\, \readData10[4]\, \readData18[4]\, 
        \readData2[4]\, \readData26[3]\, \readData_10_1_1[3]\, 
        \readData10[3]\, \readData18[3]\, \readData2[3]\, 
        \readData25[27]\, \readData_18_1_1[24]\, \readData9[27]\, 
        \readData17[27]\, \readData1[27]\, \readData25[25]\, 
        \readData_18_1_1[23]\, \readData9[25]\, \readData17[25]\, 
        \readData1[25]\, \readData26[34]\, \readData_10_1_1[31]\, 
        \readData10[34]\, \readData18[34]\, \readData2[34]\, 
        \readData26[18]\, \readData_10_1_1[16]\, \readData10[18]\, 
        \readData18[18]\, \readData2[18]\, \readData24[13]\, 
        \readData_3_1_1[12]\, \readData8[13]\, \readData16[13]\, 
        \readData0[13]\, \readData27[31]\, \readData_25_1_1[28]\, 
        \readData11[31]\, \readData19[31]\, \readData3[31]\, 
        \readData24[7]\, \readData_3_1_1[7]\, \readData8[7]\, 
        \readData16[7]\, \readData0[7]\, \readData26[29]\, 
        \readData_10_1_1[26]\, \readData10[29]\, \readData18[29]\, 
        \readData2[29]\, \readData28[31]\, \readData_6_1_1[28]\, 
        \readData12[31]\, \readData20[31]\, \readData4[31]\, 
        \readData26[21]\, \readData_10_1_1[19]\, \readData10[21]\, 
        \readData18[21]\, \readData2[21]\, \readData26[20]\, 
        \readData_10_1_1[18]\, \readData10[20]\, \readData18[20]\, 
        \readData2[20]\, \readData24[34]\, \readData_3_1_1[31]\, 
        \readData8[34]\, \readData16[34]\, \readData0[34]\, 
        \readData29[19]\, \readData_21_1_1[17]\, \readData13[19]\, 
        \readData21[19]\, \readData5[19]\, \readData24[30]\, 
        \readData_3_1_1[27]\, \readData8[30]\, \readData16[30]\, 
        \readData0[30]\, \readData26[2]\, \readData_10_1_1[2]\, 
        \readData10[2]\, \readData18[2]\, \readData2[2]\, 
        \readData24[22]\, \readData_3_1_1[20]\, \readData8[22]\, 
        \readData16[22]\, \readData0[22]\, \readData24[21]\, 
        \readData_3_1_1[19]\, \readData8[21]\, \readData16[21]\, 
        \readData0[21]\, \readData24[18]\, \readData_3_1_1[16]\, 
        \readData8[18]\, \readData16[18]\, \readData0[18]\, 
        \readData25[21]\, \readData_18_1_1[19]\, \readData9[21]\, 
        \readData17[21]\, \readData1[21]\, \readData26[16]\, 
        \readData_10_1_1[15]\, \readData10[16]\, \readData18[16]\, 
        \readData2[16]\, \readData24[12]\, \readData_3_1_1[11]\, 
        \readData8[12]\, \readData16[12]\, \readData0[12]\, 
        \readData25[14]\, \readData_18_1_1[13]\, \readData9[14]\, 
        \readData17[14]\, \readData1[14]\, \readData26[30]\, 
        \readData_10_1_1[27]\, \readData10[30]\, \readData18[30]\, 
        \readData2[30]\, \readData26[28]\, \readData_10_1_1[25]\, 
        \readData10[28]\, \readData18[28]\, \readData2[28]\, 
        \readData24[4]\, \readData_3_1_1[4]\, \readData8[4]\, 
        \readData16[4]\, \readData0[4]\, \readData26[27]\, 
        \readData_10_1_1[24]\, \readData10[27]\, \readData18[27]\, 
        \readData2[27]\, \readData26[23]\, \readData_10_1_1[21]\, 
        \readData10[23]\, \readData18[23]\, \readData2[23]\, 
        \readData25[31]\, \readData_18_1_1[28]\, \readData9[31]\, 
        \readData17[31]\, \readData1[31]\, \readData26[33]\, 
        \readData_10_1_1[30]\, \readData10[33]\, \readData18[33]\, 
        \readData2[33]\, \readData25[13]\, \readData_18_1_1[12]\, 
        \readData9[13]\, \readData17[13]\, \readData1[13]\, 
        \readData26[15]\, \readData_10_1_1[14]\, \readData10[15]\, 
        \readData18[15]\, \readData2[15]\, \readData24[3]\, 
        \readData_3_1_1[3]\, \readData8[3]\, \readData16[3]\, 
        \readData0[3]\, \readData28[25]\, \readData_6_1_1[23]\, 
        \readData12[25]\, \readData20[25]\, \readData4[25]\, 
        \readData26[12]\, \readData_10_1_1[11]\, \readData10[12]\, 
        \readData18[12]\, \readData2[12]\, \readData26[24]\, 
        \readData_10_1_1[22]\, \readData10[24]\, \readData18[24]\, 
        \readData2[24]\, \readData26[5]\, \readData_10_1_1[5]\, 
        \readData10[5]\, \readData18[5]\, \readData2[5]\, 
        \readData24[27]\, \readData_3_1_1[24]\, \readData8[27]\, 
        \readData16[27]\, \readData0[27]\, \readData26[9]\, 
        \readData_10_1_1[8]\, \readData10[9]\, \readData18[9]\, 
        \readData2[9]\, readdata_xhdl1401_1, readdata_xhdl1414_1, 
        readdata_xhdl1403_0, readdata_xhdl1419_0_a2_0, N_1150, 
        N_1149, N_1147, N_1143, N_1168, N_1148, N_1144, 
        \wen_b12_1[0]\, \wen_b12_1[1]\, \wen_b13_1[0]\, 
        \wen_b13_1[1]\, \wen_b16_1[0]\, \wen_b16_1[1]\, 
        \wen_b17_1[0]\, \wen_b17_1[1]\, \wen_b19_1[0]\, 
        \wen_b19_1[1]\, \wen_b20_1[0]\, \wen_b20_1[1]\, 
        \wen_b2_1[0]\, \wen_b2_1[1]\, \wen_b4_1[0]\, 
        \wen_b4_1[1]\, \wen_b5_1[0]\, \wen_b5_1[1]\, 
        \wen_a12_1[0]\, \wen_a12_1[1]\, \wen_a13_1[0]\, 
        \wen_a13_1[1]\, \wen_a16_1[0]\, \wen_a16_1[1]\, 
        \wen_a17_1[0]\, \wen_a17_1[1]\, \wen_a19_1[0]\, 
        \wen_a19_1[1]\, \wen_a20_1[0]\, \wen_a20_1[1]\, 
        \wen_a31_1[0]\, \wen_a31_1[1]\, \wen_b31_1[0]\, 
        \wen_b31_1[1]\, \wen_a2_1[0]\, \wen_a2_1[1]\, 
        \wen_a4_1[0]\, \wen_a5_1[0]\, \wen_a5_1[1]\, 
        \wen_b18_1[0]\, \wen_b18_1[1]\, \wen_b0_1[0]\, 
        \wen_b0_1[1]\, \wen_b1_1[0]\, \wen_b1_1[1]\, 
        \wen_b3_1[0]\, \wen_b3_1[1]\, \wen_a18_1[0]\, 
        \wen_a18_1[1]\, \wen_a0_1[0]\, \wen_a0_1[1]\, 
        \wen_a1_1[0]\, \wen_a1_1[1]\, \wen_a3_1[0]\, 
        \wen_a3_1[1]\, \wen_a4_1[1]\, \wen_b_m[0]\, \wen_b_m[1]\, 
        \wen_b22_1[0]\, \wen_b22_1[1]\, \wen_b23_1[0]\, 
        \wen_b23_1[1]\, \wen_b24_1[0]\, \wen_b24_1[1]\, 
        \wen_b25_1[0]\, \wen_b25_1[1]\, \wen_b26_1[0]\, 
        \wen_b26_1[1]\, \wen_b27_1[0]\, \wen_b27_1[1]\, 
        \wen_b28_1[0]\, \wen_b28_1[1]\, \wen_b29_1[0]\, 
        \wen_b29_1[1]\, \wen_b30_1[0]\, \wen_b30_1[1]\, 
        \wen_b6_1[0]\, \wen_b6_1[1]\, \wen_b7_1[0]\, 
        \wen_b7_1[1]\, \wen_b8_1[0]\, \wen_b8_1[1]\, 
        \wen_b9_1[0]\, \wen_b9_1[1]\, \wen_b10_1[0]\, 
        \wen_b10_1[1]\, \wen_b11_1[0]\, \wen_b11_1[1]\, 
        \wen_b14_1[0]\, \wen_b14_1[1]\, \wen_b15_1[0]\, 
        \wen_b15_1[1]\, \wen_a_m[0]\, \wen_a_m[1]\, 
        \wen_a23_1[0]\, \wen_a23_1[1]\, \wen_a24_1[0]\, 
        \wen_a24_1[1]\, \wen_a25_1[0]\, \wen_a25_1[1]\, 
        \wen_a26_1[0]\, \wen_a26_1[1]\, \wen_a27_1[0]\, 
        \wen_a27_1[1]\, \wen_a28_1[0]\, \wen_a28_1[1]\, 
        \wen_a29_1[0]\, \wen_a29_1[1]\, \wen_a30_1[0]\, 
        \wen_a30_1[1]\, \wen_a7_1[0]\, \wen_a7_1[1]\, 
        \wen_a8_1[0]\, \wen_a8_1[1]\, \wen_a9_1[0]\, 
        \wen_a9_1[1]\, \wen_a10_1[0]\, \wen_a10_1[1]\, 
        \wen_a11_1[0]\, \wen_a11_1[1]\, \wen_a14_1[0]\, 
        \wen_a14_1[1]\, \wen_a15_1[0]\, \wen_a15_1[1]\, 
        \wen_a21_1[0]\, \wen_a21_1[1]\, \wen_a6_1[0]\, 
        \wen_a6_1[1]\, VCC_net_1, GND_net_1 : std_logic;
    signal nc123, nc121, nc47, nc113, nc111, nc34, nc98, nc89, 
        nc70, nc60, nc105, nc74, nc120, nc119, nc64, nc110, nc9, 
        nc92, nc91, nc13, nc23, nc55, nc80, nc33, nc84, nc16, 
        nc26, nc45, nc73, nc58, nc63, nc27, nc17, nc127, nc99, 
        nc126, nc117, nc36, nc116, nc48, nc37, nc5, nc103, nc101, 
        nc52, nc76, nc51, nc66, nc77, nc67, nc4, nc124, nc109, 
        nc42, nc114, nc100, nc83, nc41, nc90, nc94, nc122, nc112, 
        nc86, nc59, nc25, nc15, nc87, nc35, nc49, nc28, nc18, 
        nc128, nc107, nc118, nc106, nc75, nc65, nc38, nc93, nc1, 
        nc2, nc50, nc22, nc12, nc21, nc11, nc78, nc54, nc68, nc3, 
        nc32, nc104, nc40, nc31, nc96, nc44, nc7, nc97, nc85, 
        nc72, nc6, nc71, nc62, nc61, nc125, nc115, nc102, nc19, 
        nc29, nc88, nc53, nc39, nc8, nc82, nc108, nc81, nc79, 
        nc43, nc69, nc56, nc20, nc10, nc57, nc95, nc24, nc14, 
        nc46, nc30 : std_logic;

begin 


    block2_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem_m3(3), Y => \wen_b2_1[1]\);
    
    \readData_31_am_RNO_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[22]\, D => \readData6[22]\, Y => 
        \readData_13_1_1[20]\);
    
    \readData_31_am_RNO_0[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[10]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[9]\, D => \readData10[10]\, Y => 
        N_379);
    
    \readData_31_am_RNO_0[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[18]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[16]\, D => \readData10[18]\, Y => 
        N_386);
    
    \readData_31_am_1_1_RNO_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[22]\, D => \readData4[22]\, Y => 
        \readData_6_1_1[20]\);
    
    block28_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem_m3(3), Y => \wen_b28_1[1]\);
    
    \readData_31_bm[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_970, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[24]_net_1\, D => N_874, Y => 
        \readData_31_bm[24]_net_1\);
    
    \readData_31_am_RNO_0[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[3]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[3]\, D => \readData10[3]\, Y => N_373);
    
    \readData_31_am_1_1_RNO_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[1]\, D => \readData4[1]\, Y => 
        \readData_6_1_1[1]\);
    
    block19_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem_m3(2), Y => \wen_b19_1[0]\);
    
    \readData_31_am_RNO[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[22]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[20]\, D => \readData14[22]\, Y => 
        N_486);
    
    \readData_31_am_1_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_243, D => N_147, Y => \readData_31_am_1_1[1]_net_1\);
    
    \readData_31_am_RNO[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[0]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[0]\, D => \readData14[0]\, Y => N_466);
    
    \readData_31_bm_RNO_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[3]\, D => \readData7[3]\, Y => 
        \readData_28_1_1[3]\);
    
    \readData_31_am_1_1_RNO_2[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[5]\, D => \readData0[5]\, Y => 
        \readData_3_1_1[5]\);
    
    \readData_31_am[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_487, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[21]_net_1\, D => N_391, Y => 
        \readData_31_am[21]_net_1\);
    
    block28_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(0), Y => \wen_a28_1[0]\);
    
    \readData_31_am[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_489, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[23]_net_1\, D => N_393, Y => 
        \readData_31_am[23]_net_1\);
    
    block31_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(0), Y => \wen_a31_1[0]\);
    
    \readData_31_bm[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_972, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[26]_net_1\, D => N_876, Y => 
        \readData_31_bm[26]_net_1\);
    
    \readData_31_am_1_1_RNO_2[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[27]\, D => \readData0[27]\, Y => 
        \readData_3_1_1[24]\);
    
    \readData_31_bm_RNO_2[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[0]\, D => \readData3[0]\, Y => 
        \readData_25_1_1[0]\);
    
    block7_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem_m3(2), Y => \wen_b7_1[0]\);
    
    \readData_31_am_RNO_0[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[21]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[19]\, D => \readData10[21]\, Y => 
        N_389);
    
    block6_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(1), Y => \wen_a6_1[1]\);
    
    \readData_31_am_1_1_RNO[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[9]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[8]\, D => \readData12[9]\, Y => N_250);
    
    \readData_31_bm_RNO_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[0]\, D => \readData7[0]\, Y => 
        \readData_28_1_1[0]\);
    
    \readData_31_am_1_1_RNO_2[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[28]\, D => \readData0[28]\, Y => 
        \readData_3_1_1[25]\);
    
    \readData_31_am_RNO_2[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[29]\, D => \readData2[29]\, Y => 
        \readData_10_1_1[26]\);
    
    \readData_31_am_RNO_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[7]\, D => \readData6[7]\, Y => 
        \readData_13_1_1[7]\);
    
    \readData_31_am_RNO_0[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[15]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[14]\, D => \readData10[15]\, Y => 
        N_384);
    
    \readData_31_ns[22]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[22]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[22]_net_1\, Y => 
        ram_rdata(22));
    
    block2_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(0), Y => \wen_a2_1[0]\);
    
    block10_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem_m3(3), Y => \wen_b10_1[1]\);
    
    \readData_31_bm_RNO[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[19]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[17]\, D => \readData15[19]\, Y => 
        N_963);
    
    \readData_31_bm_1_1_RNO_2[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[14]\, D => \readData1[14]\, Y => 
        \readData_18_1_1[13]\);
    
    block1_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem(0), Y => 
        \wen_a1_1[0]\);
    
    \readData_31_am_RNO[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[12]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[11]\, D => \readData14[12]\, Y => 
        N_477);
    
    block15_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem_m3(3), Y => \wen_b15_1[1]\);
    
    \readData_31_bm_1_1_RNO_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[14]\, D => \readData5[14]\, Y => 
        \readData_21_1_1[13]\);
    
    \readData_31_bm_1_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_731, D => N_635, Y => \readData_31_bm_1_1[9]_net_1\);
    
    block16_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem_m3(2), Y => 
        \wen_b16_1[0]\);
    
    \readData_31_bm_RNO[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[10]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[9]\, D => \readData15[10]\, Y => 
        N_955);
    
    \readData_31_am_RNO_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[25]\, D => \readData6[25]\, Y => 
        \readData_13_1_1[23]\);
    
    block26_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem_m3(3), Y => \wen_b26_1[1]\);
    
    block26_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(0), Y => \wen_a26_1[0]\);
    
    block23_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem_m3(3), Y => \wen_b23_1[1]\);
    
    \readData_31_bm_1_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_747, D => N_651, Y => 
        \readData_31_bm_1_1[25]_net_1\);
    
    \readData_31_bm_RNO[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[20]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[18]\, D => \readData15[20]\, Y => 
        N_964);
    
    \readData_31_am_RNO_2[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[32]\, D => \readData2[32]\, Y => 
        \readData_10_1_1[29]\);
    
    block8_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem_m3(2), Y => \wen_b8_1[0]\);
    
    \readData_31_am[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_471, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[5]_net_1\, D => N_375, Y => 
        \readData_31_am[5]_net_1\);
    
    block11_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(0), Y => \wen_a11_1[0]\);
    
    \readData_31_am_RNO_2[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[27]\, D => \readData2[27]\, Y => 
        \readData_10_1_1[24]\);
    
    \readData_31_am_1_1_RNO_2[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[21]\, D => \readData0[21]\, Y => 
        \readData_3_1_1[19]\);
    
    block10 : RAM1K18
      port map(A_DOUT(17) => nc123, A_DOUT(16) => 
        \readData10[16]\, A_DOUT(15) => \readData10[15]\, 
        A_DOUT(14) => \readData10[14]\, A_DOUT(13) => 
        \readData10[13]\, A_DOUT(12) => \readData10[12]\, 
        A_DOUT(11) => \readData10[11]\, A_DOUT(10) => 
        \readData10[10]\, A_DOUT(9) => \readData10[9]\, A_DOUT(8)
         => nc121, A_DOUT(7) => \readData10[7]\, A_DOUT(6) => 
        \readData10[6]\, A_DOUT(5) => \readData10[5]\, A_DOUT(4)
         => \readData10[4]\, A_DOUT(3) => \readData10[3]\, 
        A_DOUT(2) => \readData10[2]\, A_DOUT(1) => 
        \readData10[1]\, A_DOUT(0) => \readData10[0]\, B_DOUT(17)
         => nc47, B_DOUT(16) => \readData10[34]\, B_DOUT(15) => 
        \readData10[33]\, B_DOUT(14) => \readData10[32]\, 
        B_DOUT(13) => \readData10[31]\, B_DOUT(12) => 
        \readData10[30]\, B_DOUT(11) => \readData10[29]\, 
        B_DOUT(10) => \readData10[28]\, B_DOUT(9) => 
        \readData10[27]\, B_DOUT(8) => nc113, B_DOUT(7) => 
        \readData10[25]\, B_DOUT(6) => \readData10[24]\, 
        B_DOUT(5) => \readData10[23]\, B_DOUT(4) => 
        \readData10[22]\, B_DOUT(3) => \readData10[21]\, 
        B_DOUT(2) => \readData10[20]\, B_DOUT(1) => 
        \readData10[19]\, B_DOUT(0) => \readData10[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a10_1[1]\, A_WEN(0) => \wen_a10_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b10_1[1]\, 
        B_WEN(0) => \wen_b10_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_1_1_RNO[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[11]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[10]\, D => \readData12[11]\, Y => 
        N_252);
    
    \readData_31_am_RNO_0[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[0]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[0]\, D => \readData10[0]\, Y => N_370);
    
    block23_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(1), Y => \wen_a23_1[1]\);
    
    \readData_31_am_RNO_0[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[28]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[25]\, D => \readData10[28]\, Y => 
        N_395);
    
    \readData_31_am_1_1_RNO_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[21]\, D => \readData4[21]\, Y => 
        \readData_6_1_1[19]\);
    
    \readData_31_bm_1_1_RNO_2[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[21]\, D => \readData1[21]\, Y => 
        \readData_18_1_1[19]\);
    
    \readData_31_bm_1_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_741, D => N_645, Y => 
        \readData_31_bm_1_1[19]_net_1\);
    
    \readData_31_am_1_1_RNO_0[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[19]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[17]\, D => \readData8[19]\, Y => 
        N_163);
    
    \readData_31_bm_RNO_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[27]\, D => \readData7[27]\, Y => 
        \readData_28_1_1[24]\);
    
    \readData_31_bm_RNO[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[9]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[8]\, D => \readData15[9]\, Y => N_954);
    
    \readData_31_bm_RNO_2[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[1]\, D => \readData3[1]\, Y => 
        \readData_25_1_1[1]\);
    
    \readData_31_bm_1_1_RNO_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[21]\, D => \readData5[21]\, Y => 
        \readData_21_1_1[19]\);
    
    \readData_31_am_1_1_RNO_0[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[3]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[3]\, D => \readData8[3]\, Y => N_149);
    
    \readData_31_bm_RNO_0[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[18]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[16]\, D => \readData11[18]\, Y => 
        N_866);
    
    \readData_31_bm_1_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_733, D => N_637, Y => 
        \readData_31_bm_1_1[11]_net_1\);
    
    block21 : RAM1K18
      port map(A_DOUT(17) => nc111, A_DOUT(16) => 
        \readData21[16]\, A_DOUT(15) => \readData21[15]\, 
        A_DOUT(14) => \readData21[14]\, A_DOUT(13) => 
        \readData21[13]\, A_DOUT(12) => \readData21[12]\, 
        A_DOUT(11) => \readData21[11]\, A_DOUT(10) => 
        \readData21[10]\, A_DOUT(9) => \readData21[9]\, A_DOUT(8)
         => nc34, A_DOUT(7) => \readData21[7]\, A_DOUT(6) => 
        \readData21[6]\, A_DOUT(5) => \readData21[5]\, A_DOUT(4)
         => \readData21[4]\, A_DOUT(3) => \readData21[3]\, 
        A_DOUT(2) => \readData21[2]\, A_DOUT(1) => 
        \readData21[1]\, A_DOUT(0) => \readData21[0]\, B_DOUT(17)
         => nc98, B_DOUT(16) => \readData21[34]\, B_DOUT(15) => 
        \readData21[33]\, B_DOUT(14) => \readData21[32]\, 
        B_DOUT(13) => \readData21[31]\, B_DOUT(12) => 
        \readData21[30]\, B_DOUT(11) => \readData21[29]\, 
        B_DOUT(10) => \readData21[28]\, B_DOUT(9) => 
        \readData21[27]\, B_DOUT(8) => nc89, B_DOUT(7) => 
        \readData21[25]\, B_DOUT(6) => \readData21[24]\, 
        B_DOUT(5) => \readData21[23]\, B_DOUT(4) => 
        \readData21[22]\, B_DOUT(3) => \readData21[21]\, 
        B_DOUT(2) => \readData21[20]\, B_DOUT(1) => 
        \readData21[19]\, B_DOUT(0) => \readData21[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a21_1[1]\, A_WEN(0) => \wen_a21_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b_m[1]\, 
        B_WEN(0) => \wen_b_m[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_1_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_258, D => N_162, Y => 
        \readData_31_am_1_1[16]_net_1\);
    
    \readData_31_bm_RNO_0[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[34]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[31]\, D => \readData11[34]\, Y => 
        N_881);
    
    block8 : RAM1K18
      port map(A_DOUT(17) => nc70, A_DOUT(16) => \readData8[16]\, 
        A_DOUT(15) => \readData8[15]\, A_DOUT(14) => 
        \readData8[14]\, A_DOUT(13) => \readData8[13]\, 
        A_DOUT(12) => \readData8[12]\, A_DOUT(11) => 
        \readData8[11]\, A_DOUT(10) => \readData8[10]\, A_DOUT(9)
         => \readData8[9]\, A_DOUT(8) => nc60, A_DOUT(7) => 
        \readData8[7]\, A_DOUT(6) => \readData8[6]\, A_DOUT(5)
         => \readData8[5]\, A_DOUT(4) => \readData8[4]\, 
        A_DOUT(3) => \readData8[3]\, A_DOUT(2) => \readData8[2]\, 
        A_DOUT(1) => \readData8[1]\, A_DOUT(0) => \readData8[0]\, 
        B_DOUT(17) => nc105, B_DOUT(16) => \readData8[34]\, 
        B_DOUT(15) => \readData8[33]\, B_DOUT(14) => 
        \readData8[32]\, B_DOUT(13) => \readData8[31]\, 
        B_DOUT(12) => \readData8[30]\, B_DOUT(11) => 
        \readData8[29]\, B_DOUT(10) => \readData8[28]\, B_DOUT(9)
         => \readData8[27]\, B_DOUT(8) => nc74, B_DOUT(7) => 
        \readData8[25]\, B_DOUT(6) => \readData8[24]\, B_DOUT(5)
         => \readData8[23]\, B_DOUT(4) => \readData8[22]\, 
        B_DOUT(3) => \readData8[21]\, B_DOUT(2) => 
        \readData8[20]\, B_DOUT(1) => \readData8[19]\, B_DOUT(0)
         => \readData8[18]\, BUSY => OPEN, A_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => N_375_i_0, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        N_72_i_0, A_DIN(15) => N_70_i_0, A_DIN(14) => N_68_i_0, 
        A_DIN(13) => N_66_i_0, A_DIN(12) => N_64_i_0, A_DIN(11)
         => N_58_i_0, A_DIN(10) => N_56_i_0, A_DIN(9) => N_54_i_0, 
        A_DIN(8) => GND_net_1, A_DIN(7) => N_52_i_0, A_DIN(6) => 
        N_50_i_0, A_DIN(5) => N_48_i_0, A_DIN(4) => N_46_i_0, 
        A_DIN(3) => N_44_i_0, A_DIN(2) => N_42_i_0, A_DIN(1) => 
        N_40_i_0, A_DIN(0) => N_38_i_0, A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a8_1[1]\, 
        A_WEN(0) => \wen_a8_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b8_1[1]\, 
        B_WEN(0) => \wen_b8_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block12_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem_m3(2), Y => \wen_b12_1[0]\);
    
    \readData_31_bm_RNO[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[28]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[25]\, D => \readData15[28]\, Y => 
        N_971);
    
    \readData_31_am_RNO_0[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[34]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[31]\, D => \readData10[34]\, Y => 
        N_401);
    
    \readData_31_bm_RNO_0[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[30]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[27]\, D => \readData11[30]\, Y => 
        N_877);
    
    \readData_31_bm[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_974, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[28]_net_1\, D => N_878, Y => 
        \readData_31_bm[28]_net_1\);
    
    \readData_31_am_RNO_2[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[16]\, D => \readData2[16]\, Y => 
        \readData_10_1_1[15]\);
    
    \readData_31_bm_RNO_0[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[21]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[19]\, D => \readData11[21]\, Y => 
        N_869);
    
    \readData_31_am_1_1_RNO_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[27]\, D => \readData4[27]\, Y => 
        \readData_6_1_1[24]\);
    
    block22 : RAM1K18
      port map(A_DOUT(17) => nc120, A_DOUT(16) => 
        \readData22[16]\, A_DOUT(15) => \readData22[15]\, 
        A_DOUT(14) => \readData22[14]\, A_DOUT(13) => 
        \readData22[13]\, A_DOUT(12) => \readData22[12]\, 
        A_DOUT(11) => \readData22[11]\, A_DOUT(10) => 
        \readData22[10]\, A_DOUT(9) => \readData22[9]\, A_DOUT(8)
         => nc119, A_DOUT(7) => \readData22[7]\, A_DOUT(6) => 
        \readData22[6]\, A_DOUT(5) => \readData22[5]\, A_DOUT(4)
         => \readData22[4]\, A_DOUT(3) => \readData22[3]\, 
        A_DOUT(2) => \readData22[2]\, A_DOUT(1) => 
        \readData22[1]\, A_DOUT(0) => \readData22[0]\, B_DOUT(17)
         => nc64, B_DOUT(16) => \readData22[34]\, B_DOUT(15) => 
        \readData22[33]\, B_DOUT(14) => \readData22[32]\, 
        B_DOUT(13) => \readData22[31]\, B_DOUT(12) => 
        \readData22[30]\, B_DOUT(11) => \readData22[29]\, 
        B_DOUT(10) => \readData22[28]\, B_DOUT(9) => 
        \readData22[27]\, B_DOUT(8) => nc110, B_DOUT(7) => 
        \readData22[25]\, B_DOUT(6) => \readData22[24]\, 
        B_DOUT(5) => \readData22[23]\, B_DOUT(4) => 
        \readData22[22]\, B_DOUT(3) => \readData22[21]\, 
        B_DOUT(2) => \readData22[20]\, B_DOUT(1) => 
        \readData22[19]\, B_DOUT(0) => \readData22[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a_m[1]\, A_WEN(0) => \wen_a_m[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b22_1[1]\, 
        B_WEN(0) => \wen_b22_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_ns[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[5]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[5]_net_1\, Y => 
        ram_rdata(5));
    
    \readData_31_ns[25]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[25]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[25]_net_1\, Y => 
        ram_rdata(25));
    
    \readData_31_am_RNO_0[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[6]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[6]\, D => \readData10[6]\, Y => N_376);
    
    \readData_31_bm_1_1_RNO_0[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[20]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[18]\, D => \readData9[20]\, Y => 
        N_644);
    
    \readData_31_am_RNO_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[16]\, D => \readData6[16]\, Y => 
        \readData_13_1_1[15]\);
    
    \readData_31_bm[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_959, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[13]_net_1\, D => N_863, Y => 
        \readData_31_bm[13]_net_1\);
    
    \readData_31_am_1_1_RNO[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[22]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[20]\, D => \readData12[22]\, Y => 
        N_262);
    
    \readData_31_am_1_1_RNO_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[10]\, D => \readData4[10]\, Y => 
        \readData_6_1_1[9]\);
    
    block23 : RAM1K18
      port map(A_DOUT(17) => nc9, A_DOUT(16) => \readData23[16]\, 
        A_DOUT(15) => \readData23[15]\, A_DOUT(14) => 
        \readData23[14]\, A_DOUT(13) => \readData23[13]\, 
        A_DOUT(12) => \readData23[12]\, A_DOUT(11) => 
        \readData23[11]\, A_DOUT(10) => \readData23[10]\, 
        A_DOUT(9) => \readData23[9]\, A_DOUT(8) => nc92, 
        A_DOUT(7) => \readData23[7]\, A_DOUT(6) => 
        \readData23[6]\, A_DOUT(5) => \readData23[5]\, A_DOUT(4)
         => \readData23[4]\, A_DOUT(3) => \readData23[3]\, 
        A_DOUT(2) => \readData23[2]\, A_DOUT(1) => 
        \readData23[1]\, A_DOUT(0) => \readData23[0]\, B_DOUT(17)
         => nc91, B_DOUT(16) => \readData23[34]\, B_DOUT(15) => 
        \readData23[33]\, B_DOUT(14) => \readData23[32]\, 
        B_DOUT(13) => \readData23[31]\, B_DOUT(12) => 
        \readData23[30]\, B_DOUT(11) => \readData23[29]\, 
        B_DOUT(10) => \readData23[28]\, B_DOUT(9) => 
        \readData23[27]\, B_DOUT(8) => nc13, B_DOUT(7) => 
        \readData23[25]\, B_DOUT(6) => \readData23[24]\, 
        B_DOUT(5) => \readData23[23]\, B_DOUT(4) => 
        \readData23[22]\, B_DOUT(3) => \readData23[21]\, 
        B_DOUT(2) => \readData23[20]\, B_DOUT(1) => 
        \readData23[19]\, B_DOUT(0) => \readData23[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a23_1[1]\, A_WEN(0) => \wen_a23_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b23_1[1]\, 
        B_WEN(0) => \wen_b23_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[5]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[5]\, D => \readData15[5]\, Y => N_951);
    
    \readData_31_bm_RNO_0[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[2]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[2]\, D => \readData11[2]\, Y => N_852);
    
    \readData_31_am_1_1_RNO[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[3]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[3]\, D => \readData12[3]\, Y => N_245);
    
    \readData_31_am_1_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_254, D => N_158, Y => 
        \readData_31_am_1_1[12]_net_1\);
    
    \readData_31_am[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_493, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[27]_net_1\, D => N_397, Y => 
        \readData_31_am[27]_net_1\);
    
    \readData_31_am_1_1_RNO_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[28]\, D => \readData4[28]\, Y => 
        \readData_6_1_1[25]\);
    
    \readData_31_bm_RNO_2[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[29]\, D => \readData3[29]\, Y => 
        \readData_25_1_1[26]\);
    
    block13_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem_m3(2), Y => 
        \wen_b13_1[0]\);
    
    \readData_31_am_1_1_RNO[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[10]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[9]\, D => \readData12[10]\, Y => 
        N_251);
    
    \readData_31_am_1_1_RNO_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[0]\, D => \readData4[0]\, Y => 
        \readData_6_1_1[0]\);
    
    \readData_31_am_1_1_RNO[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[14]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[13]\, D => \readData12[14]\, Y => 
        N_255);
    
    \readData_31_bm_RNO_2[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[19]\, D => \readData3[19]\, Y => 
        \readData_25_1_1[17]\);
    
    \readData_31_bm_1_1_RNO_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[4]\, D => \readData5[4]\, Y => 
        \readData_21_1_1[4]\);
    
    \readData_31_bm_RNO_0[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[24]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[22]\, D => \readData11[24]\, Y => 
        N_872);
    
    \readData_31_am_RNO[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[28]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[25]\, D => \readData14[28]\, Y => 
        N_491);
    
    \readData_31_am_1_1_RNO_0[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[31]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[28]\, D => \readData8[31]\, Y => 
        N_174);
    
    block28 : RAM1K18
      port map(A_DOUT(17) => nc23, A_DOUT(16) => \readData28[16]\, 
        A_DOUT(15) => \readData28[15]\, A_DOUT(14) => 
        \readData28[14]\, A_DOUT(13) => \readData28[13]\, 
        A_DOUT(12) => \readData28[12]\, A_DOUT(11) => 
        \readData28[11]\, A_DOUT(10) => \readData28[10]\, 
        A_DOUT(9) => \readData28[9]\, A_DOUT(8) => nc55, 
        A_DOUT(7) => \readData28[7]\, A_DOUT(6) => 
        \readData28[6]\, A_DOUT(5) => \readData28[5]\, A_DOUT(4)
         => \readData28[4]\, A_DOUT(3) => \readData28[3]\, 
        A_DOUT(2) => \readData28[2]\, A_DOUT(1) => 
        \readData28[1]\, A_DOUT(0) => \readData28[0]\, B_DOUT(17)
         => nc80, B_DOUT(16) => \readData28[34]\, B_DOUT(15) => 
        \readData28[33]\, B_DOUT(14) => \readData28[32]\, 
        B_DOUT(13) => \readData28[31]\, B_DOUT(12) => 
        \readData28[30]\, B_DOUT(11) => \readData28[29]\, 
        B_DOUT(10) => \readData28[28]\, B_DOUT(9) => 
        \readData28[27]\, B_DOUT(8) => nc33, B_DOUT(7) => 
        \readData28[25]\, B_DOUT(6) => \readData28[24]\, 
        B_DOUT(5) => \readData28[23]\, B_DOUT(4) => 
        \readData28[22]\, B_DOUT(3) => \readData28[21]\, 
        B_DOUT(2) => \readData28[20]\, B_DOUT(1) => 
        \readData28[19]\, B_DOUT(0) => \readData28[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a28_1[1]\, A_WEN(0) => \wen_a28_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b28_1[1]\, 
        B_WEN(0) => \wen_b28_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_2[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[32]\, D => \readData3[32]\, Y => 
        \readData_25_1_1[29]\);
    
    \readData_31_am[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_480, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[14]_net_1\, D => N_384, Y => 
        \readData_31_am[14]_net_1\);
    
    \readData_31_bm_RNO_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[19]\, D => \readData7[19]\, Y => 
        \readData_28_1_1[17]\);
    
    \readData_31_am_RNO_2[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[4]\, D => \readData2[4]\, Y => 
        \readData_10_1_1[4]\);
    
    \readData_31_bm_1_1_RNO_0[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[6]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[6]\, D => \readData9[6]\, Y => N_632);
    
    \readData_31_bm_RNO_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[34]\, D => \readData7[34]\, Y => 
        \readData_28_1_1[31]\);
    
    \readData_31_am_RNO_0[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[24]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[22]\, D => \readData10[24]\, Y => 
        N_392);
    
    \readData_31_bm_RNO[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[34]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[31]\, D => \readData15[34]\, Y => 
        N_977);
    
    \readData_31_am_RNO_2[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[6]\, D => \readData2[6]\, Y => 
        \readData_10_1_1[6]\);
    
    \readData_31_am_1_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_266, D => N_170, Y => 
        \readData_31_am_1_1[24]_net_1\);
    
    \readData_31_ns[16]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[16]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[16]_net_1\, Y => 
        ram_rdata(16));
    
    \readData_31_am_RNO_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[34]\, D => \readData6[34]\, Y => 
        \readData_13_1_1[31]\);
    
    \readData_31_bm_RNO_0[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[14]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[13]\, D => \readData11[14]\, Y => 
        N_863);
    
    \readData_31_bm[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_965, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[19]_net_1\, D => N_869, Y => 
        \readData_31_bm[19]_net_1\);
    
    \readData_31_bm_RNO_0[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[11]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[10]\, D => \readData11[11]\, Y => 
        N_860);
    
    \readData_31_bm_RNO_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[9]\, D => \readData7[9]\, Y => 
        \readData_28_1_1[8]\);
    
    \readData_31_am[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_478, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[12]_net_1\, D => N_382, Y => 
        \readData_31_am[12]_net_1\);
    
    \readData_31_am_1_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_261, D => N_165, Y => 
        \readData_31_am_1_1[19]_net_1\);
    
    \readData_31_bm_RNO_2[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[13]\, D => \readData3[13]\, Y => 
        \readData_25_1_1[12]\);
    
    \readData_31_bm_1_1_RNO[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[0]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[0]\, D => \readData13[0]\, Y => N_722);
    
    \readData_31_bm_1_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_744, D => N_648, Y => 
        \readData_31_bm_1_1[22]_net_1\);
    
    block24_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem_m3(2), Y => \wen_b24_1[0]\);
    
    \readData_31_bm_RNO_2[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[9]\, D => \readData3[9]\, Y => 
        \readData_25_1_1[8]\);
    
    \readData_31_am_1_1_RNO_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[9]\, D => \readData4[9]\, Y => 
        \readData_6_1_1[8]\);
    
    \readData_31_bm_RNO[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[14]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[13]\, D => \readData15[14]\, Y => 
        N_959);
    
    \readData_31_bm_RNO_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[13]\, D => \readData7[13]\, Y => 
        \readData_28_1_1[12]\);
    
    \readData_31_bm_RNO[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[33]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[30]\, D => \readData15[33]\, Y => 
        N_976);
    
    \readData_31_bm[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_958, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[12]_net_1\, D => N_862, Y => 
        \readData_31_bm[12]_net_1\);
    
    \readData_31_am_RNO_2[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[13]\, D => \readData2[13]\, Y => 
        \readData_10_1_1[12]\);
    
    \readData_31_am_1_1_RNO[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[25]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[23]\, D => \readData12[25]\, Y => 
        N_265);
    
    \readData_31_am_RNO_0[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[1]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[1]\, D => \readData10[1]\, Y => N_371);
    
    block17 : RAM1K18
      port map(A_DOUT(17) => nc84, A_DOUT(16) => \readData17[16]\, 
        A_DOUT(15) => \readData17[15]\, A_DOUT(14) => 
        \readData17[14]\, A_DOUT(13) => \readData17[13]\, 
        A_DOUT(12) => \readData17[12]\, A_DOUT(11) => 
        \readData17[11]\, A_DOUT(10) => \readData17[10]\, 
        A_DOUT(9) => \readData17[9]\, A_DOUT(8) => nc16, 
        A_DOUT(7) => \readData17[7]\, A_DOUT(6) => 
        \readData17[6]\, A_DOUT(5) => \readData17[5]\, A_DOUT(4)
         => \readData17[4]\, A_DOUT(3) => \readData17[3]\, 
        A_DOUT(2) => \readData17[2]\, A_DOUT(1) => 
        \readData17[1]\, A_DOUT(0) => \readData17[0]\, B_DOUT(17)
         => nc26, B_DOUT(16) => \readData17[34]\, B_DOUT(15) => 
        \readData17[33]\, B_DOUT(14) => \readData17[32]\, 
        B_DOUT(13) => \readData17[31]\, B_DOUT(12) => 
        \readData17[30]\, B_DOUT(11) => \readData17[29]\, 
        B_DOUT(10) => \readData17[28]\, B_DOUT(9) => 
        \readData17[27]\, B_DOUT(8) => nc45, B_DOUT(7) => 
        \readData17[25]\, B_DOUT(6) => \readData17[24]\, 
        B_DOUT(5) => \readData17[23]\, B_DOUT(4) => 
        \readData17[22]\, B_DOUT(3) => \readData17[21]\, 
        B_DOUT(2) => \readData17[20]\, B_DOUT(1) => 
        \readData17[19]\, B_DOUT(0) => \readData17[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a17_1[1]\, A_WEN(0) => \wen_a17_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b17_1[1]\, 
        B_WEN(0) => \wen_b17_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \readData_31_am_1_1_RNO_2[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[31]\, D => \readData0[31]\, Y => 
        \readData_3_1_1[28]\);
    
    \readData_31_bm_1_1_RNO_2[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[9]\, D => \readData1[9]\, Y => 
        \readData_18_1_1[8]\);
    
    \readData_31_am_RNO_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[13]\, D => \readData6[13]\, Y => 
        \readData_13_1_1[12]\);
    
    \readData_31_bm_RNO_2[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[25]\, D => \readData3[25]\, Y => 
        \readData_25_1_1[23]\);
    
    block21_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem_m3(2), Y => \wen_b_m[0]\);
    
    block30_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(1), Y => \wen_a30_1[1]\);
    
    \readData_31_ns[31]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[31]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[31]_net_1\, Y => 
        ram_rdata(31));
    
    \readData_31_am_1_1_RNO_0[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[4]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[4]\, D => \readData8[4]\, Y => N_150);
    
    \readData_31_bm_RNO_2[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[22]\, D => \readData3[22]\, Y => 
        \readData_25_1_1[20]\);
    
    \readData_31_am_1_1_RNO_2[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[19]\, D => \readData0[19]\, Y => 
        \readData_3_1_1[17]\);
    
    block21_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(0), Y => \wen_a21_1[0]\);
    
    \readData_31_bm_1_1_RNO_0[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[16]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[15]\, D => \readData9[16]\, Y => 
        N_641);
    
    \readData_31_am_1_1_RNO_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[19]\, D => \readData4[19]\, Y => 
        \readData_6_1_1[17]\);
    
    \readData_31_am_1_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_249, D => N_153, Y => \readData_31_am_1_1[7]_net_1\);
    
    block7_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(1), Y => \wen_a7_1[1]\);
    
    \readData_31_bm_RNO_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[28]\, D => \readData7[28]\, Y => 
        \readData_28_1_1[25]\);
    
    block22_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem_m3(3), Y => \wen_b22_1[1]\);
    
    \readData_31_bm_1_1_RNO_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[1]\, D => \readData5[1]\, Y => 
        \readData_21_1_1[1]\);
    
    \readData_31_bm[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_951, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[5]_net_1\, D => N_855, Y => 
        \readData_31_bm[5]_net_1\);
    
    block6_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem_m3(2), Y => \wen_b6_1[0]\);
    
    \readData_31_bm[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_973, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[27]_net_1\, D => N_877, Y => 
        \readData_31_bm[27]_net_1\);
    
    \readData_31_am_1_1_RNO_0[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[25]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[23]\, D => \readData8[25]\, Y => 
        N_169);
    
    \readData_31_bm_1_1_RNO[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[14]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[13]\, D => \readData13[14]\, Y => 
        N_735);
    
    block9_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem_m3(2), Y => \wen_b9_1[0]\);
    
    \readData_31_am_1_1_RNO_0[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[9]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[8]\, D => \readData8[9]\, Y => N_154);
    
    \readData_31_bm_1_1_RNO_2[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[5]\, D => \readData1[5]\, Y => 
        \readData_18_1_1[5]\);
    
    block24_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem_m3(3), Y => \wen_b24_1[1]\);
    
    \readData_31_bm_1_1_RNO_2[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[20]\, D => \readData1[20]\, Y => 
        \readData_18_1_1[18]\);
    
    \readData_31_bm_1_1_RNO[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[21]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[19]\, D => \readData13[21]\, Y => 
        N_741);
    
    \readData_31_am_1_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_242, D => N_146, Y => \readData_31_am_1_1[0]_net_1\);
    
    \readData_31_am_1_1_RNO[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[18]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[16]\, D => \readData12[18]\, Y => 
        N_258);
    
    \readData_31_bm_1_1_RNO_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[20]\, D => \readData5[20]\, Y => 
        \readData_21_1_1[18]\);
    
    \readData_31_am_RNO_2[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[5]\, D => \readData2[5]\, Y => 
        \readData_10_1_1[5]\);
    
    block16_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(1), Y => 
        \wen_a16_1[1]\);
    
    \readData_31_am_RNO[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[10]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[9]\, D => \readData14[10]\, Y => 
        N_475);
    
    \readData_31_bm_1_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_750, D => N_654, Y => 
        \readData_31_bm_1_1[28]_net_1\);
    
    \readData_31_am_1_1_RNO_2[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[4]\, D => \readData0[4]\, Y => 
        \readData_3_1_1[4]\);
    
    \readData_31_am_RNO[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[13]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[12]\, D => \readData14[13]\, Y => 
        N_478);
    
    \readData_31_am_1_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_257, D => N_161, Y => 
        \readData_31_am_1_1[15]_net_1\);
    
    \readData_31_bm_RNO[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[13]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[12]\, D => \readData15[13]\, Y => 
        N_958);
    
    \readData_31_am_RNO_0[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[4]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[4]\, D => \readData10[4]\, Y => N_374);
    
    block31 : RAM1K18
      port map(A_DOUT(17) => nc73, A_DOUT(16) => \readData31[16]\, 
        A_DOUT(15) => \readData31[15]\, A_DOUT(14) => 
        \readData31[14]\, A_DOUT(13) => \readData31[13]\, 
        A_DOUT(12) => \readData31[12]\, A_DOUT(11) => 
        \readData31[11]\, A_DOUT(10) => \readData31[10]\, 
        A_DOUT(9) => \readData31[9]\, A_DOUT(8) => nc58, 
        A_DOUT(7) => \readData31[7]\, A_DOUT(6) => 
        \readData31[6]\, A_DOUT(5) => \readData31[5]\, A_DOUT(4)
         => \readData31[4]\, A_DOUT(3) => \readData31[3]\, 
        A_DOUT(2) => \readData31[2]\, A_DOUT(1) => 
        \readData31[1]\, A_DOUT(0) => \readData31[0]\, B_DOUT(17)
         => nc63, B_DOUT(16) => \readData31[34]\, B_DOUT(15) => 
        \readData31[33]\, B_DOUT(14) => \readData31[32]\, 
        B_DOUT(13) => \readData31[31]\, B_DOUT(12) => 
        \readData31[30]\, B_DOUT(11) => \readData31[29]\, 
        B_DOUT(10) => \readData31[28]\, B_DOUT(9) => 
        \readData31[27]\, B_DOUT(8) => nc27, B_DOUT(7) => 
        \readData31[25]\, B_DOUT(6) => \readData31[24]\, 
        B_DOUT(5) => \readData31[23]\, B_DOUT(4) => 
        \readData31[22]\, B_DOUT(3) => \readData31[21]\, 
        B_DOUT(2) => \readData31[20]\, B_DOUT(1) => 
        \readData31[19]\, B_DOUT(0) => \readData31[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a31_1[1]\, A_WEN(0) => \wen_a31_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b31_1[1]\, 
        B_WEN(0) => \wen_b31_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_971, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[25]_net_1\, D => N_875, Y => 
        \readData_31_bm[25]_net_1\);
    
    \readData_31_am_RNO_0[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[33]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[30]\, D => \readData10[33]\, Y => 
        N_400);
    
    block13_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(0), Y => 
        \wen_a13_1[0]\);
    
    \readData_31_am_1_1_RNO_2[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[1]\, D => \readData0[1]\, Y => 
        \readData_3_1_1[1]\);
    
    block14_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(1), Y => \wen_a14_1[1]\);
    
    \readData_31_am_1_1_RNO_0[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[10]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[9]\, D => \readData8[10]\, Y => N_155);
    
    \readData_31_am_1_1_RNO_2[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[25]\, D => \readData0[25]\, Y => 
        \readData_3_1_1[23]\);
    
    \readData_31_ns[28]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[28]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[28]_net_1\, Y => 
        ram_rdata(28));
    
    \readData_31_bm_1_1_RNO[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[25]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[23]\, D => \readData13[25]\, Y => 
        N_745);
    
    block26 : RAM1K18
      port map(A_DOUT(17) => nc17, A_DOUT(16) => \readData26[16]\, 
        A_DOUT(15) => \readData26[15]\, A_DOUT(14) => 
        \readData26[14]\, A_DOUT(13) => \readData26[13]\, 
        A_DOUT(12) => \readData26[12]\, A_DOUT(11) => 
        \readData26[11]\, A_DOUT(10) => \readData26[10]\, 
        A_DOUT(9) => \readData26[9]\, A_DOUT(8) => nc127, 
        A_DOUT(7) => \readData26[7]\, A_DOUT(6) => 
        \readData26[6]\, A_DOUT(5) => \readData26[5]\, A_DOUT(4)
         => \readData26[4]\, A_DOUT(3) => \readData26[3]\, 
        A_DOUT(2) => \readData26[2]\, A_DOUT(1) => 
        \readData26[1]\, A_DOUT(0) => \readData26[0]\, B_DOUT(17)
         => nc99, B_DOUT(16) => \readData26[34]\, B_DOUT(15) => 
        \readData26[33]\, B_DOUT(14) => \readData26[32]\, 
        B_DOUT(13) => \readData26[31]\, B_DOUT(12) => 
        \readData26[30]\, B_DOUT(11) => \readData26[29]\, 
        B_DOUT(10) => \readData26[28]\, B_DOUT(9) => 
        \readData26[27]\, B_DOUT(8) => nc126, B_DOUT(7) => 
        \readData26[25]\, B_DOUT(6) => \readData26[24]\, 
        B_DOUT(5) => \readData26[23]\, B_DOUT(4) => 
        \readData26[22]\, B_DOUT(3) => \readData26[21]\, 
        B_DOUT(2) => \readData26[20]\, B_DOUT(1) => 
        \readData26[19]\, B_DOUT(0) => \readData26[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a26_1[1]\, A_WEN(0) => \wen_a26_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b26_1[1]\, 
        B_WEN(0) => \wen_b26_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_1_1_RNO_0[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[12]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[11]\, D => \readData8[12]\, Y => 
        N_157);
    
    \readData_31_ns[29]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[29]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[29]_net_1\, Y => 
        ram_rdata(29));
    
    block10_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(1), Y => \wen_a10_1[1]\);
    
    \readData_31_bm_RNO[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[1]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[1]\, D => \readData15[1]\, Y => N_947);
    
    \readData_31_bm_RNO[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[4]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[4]\, D => \readData15[4]\, Y => N_950);
    
    \readData_31_bm_1_1_RNO_0[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[11]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[10]\, D => \readData9[11]\, Y => 
        N_636);
    
    \readData_31_bm_1_1_RNO[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[32]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[29]\, D => \readData13[32]\, Y => 
        N_751);
    
    \readData_31_am_RNO[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[9]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[8]\, D => \readData14[9]\, Y => N_474);
    
    \readData_31_bm_RNO[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[32]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[29]\, D => \readData15[32]\, Y => 
        N_975);
    
    \readData_31_am_1_1_RNO_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[31]\, D => \readData4[31]\, Y => 
        \readData_6_1_1[28]\);
    
    \readData_31_am_1_1_RNO_0[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[1]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[1]\, D => \readData8[1]\, Y => N_147);
    
    \readData_31_bm_RNO_0[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[5]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[5]\, D => \readData11[5]\, Y => N_855);
    
    \readData_31_am_1_1_RNO[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[29]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[26]\, D => \readData12[29]\, Y => 
        N_268);
    
    \readData_31_am_1_1_RNO_0[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[33]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[30]\, D => \readData8[33]\, Y => 
        N_176);
    
    \readData_31_bm[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_960, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[14]_net_1\, D => N_864, Y => 
        \readData_31_bm[14]_net_1\);
    
    \readData_31_am_1_1_RNO[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[19]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[17]\, D => \readData12[19]\, Y => 
        N_259);
    
    \readData_31_am[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_496, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[30]_net_1\, D => N_400, Y => 
        \readData_31_am[30]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[12]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[11]\, D => \readData9[12]\, Y => 
        N_637);
    
    \readData_31_bm_RNO[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[3]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[3]\, D => \readData15[3]\, Y => N_949);
    
    \readData_31_am[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_477, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[11]_net_1\, D => N_381, Y => 
        \readData_31_am[11]_net_1\);
    
    block4_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem_m3(3), Y => \wen_b4_1[1]\);
    
    \readData_31_bm_1_1_RNO_0[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[19]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[17]\, D => \readData9[19]\, Y => 
        N_643);
    
    \readData_31_am[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_479, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[13]_net_1\, D => N_383, Y => 
        \readData_31_am[13]_net_1\);
    
    \readData_31_bm_RNO_0[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[23]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[21]\, D => \readData11[23]\, Y => 
        N_871);
    
    \readData_31_bm_1_1_RNO_0[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[3]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[3]\, D => \readData9[3]\, Y => N_629);
    
    \readData_31_bm[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_962, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[16]_net_1\, D => N_866, Y => 
        \readData_31_bm[16]_net_1\);
    
    \readData_31_am_RNO_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[33]\, D => \readData6[33]\, Y => 
        \readData_13_1_1[30]\);
    
    \readData_31_bm[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_977, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[31]_net_1\, D => N_881, Y => 
        \readData_31_bm[31]_net_1\);
    
    \readData_31_am_RNO[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[5]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[5]\, D => \readData14[5]\, Y => N_471);
    
    block31_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(1), Y => \wen_a31_1[1]\);
    
    \readData_31_am_RNO_0[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[23]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[21]\, D => \readData10[23]\, Y => 
        N_391);
    
    \readData_31_am_1_1_RNO_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[3]\, D => \readData4[3]\, Y => 
        \readData_6_1_1[3]\);
    
    readdata_xhdl1401_1_0 : CFG3
      generic map(INIT => x"40")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => ahbsram_addr(12), Y => readdata_xhdl1401_1);
    
    block6_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem_m3(3), Y => \wen_b6_1[1]\);
    
    block9_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(1), Y => \wen_a9_1[1]\);
    
    block18_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(14), C
         => readdata_xhdl1401_1, D => sram_wen_mem(1), Y => 
        \wen_a18_1[1]\);
    
    \readData_31_bm_1_1_RNO_2[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[16]\, D => \readData1[16]\, Y => 
        \readData_18_1_1[15]\);
    
    \readData_31_am[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_467, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[1]_net_1\, D => N_371, Y => 
        \readData_31_am[1]_net_1\);
    
    \readData_31_am_1_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_247, D => N_151, Y => \readData_31_am_1_1[5]_net_1\);
    
    \readData_31_am[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_472, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[6]_net_1\, D => N_376, Y => 
        \readData_31_am[6]_net_1\);
    
    block8_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(1), Y => \wen_a8_1[1]\);
    
    \readData_31_ns[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[6]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[6]_net_1\, Y => 
        ram_rdata(6));
    
    \readData_31_bm_RNO_2[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[2]\, D => \readData3[2]\, Y => 
        \readData_25_1_1[2]\);
    
    \readData_31_bm_1_1_RNO_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[16]\, D => \readData5[16]\, Y => 
        \readData_21_1_1[15]\);
    
    \readData_31_bm_RNO_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[10]\, D => \readData7[10]\, Y => 
        \readData_28_1_1[9]\);
    
    \readData_31_am_1_1_RNO[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[30]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[27]\, D => \readData12[30]\, Y => 
        N_269);
    
    \readData_31_am[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_469, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[3]_net_1\, D => N_373, Y => 
        \readData_31_am[3]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[10]\, D => \readData5[10]\, Y => 
        \readData_21_1_1[9]\);
    
    \readData_31_bm_RNO_2[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[12]\, D => \readData3[12]\, Y => 
        \readData_25_1_1[11]\);
    
    \readData_31_bm_RNO_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[31]\, D => \readData7[31]\, Y => 
        \readData_28_1_1[28]\);
    
    block15_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(1), Y => \wen_a15_1[1]\);
    
    block5 : RAM1K18
      port map(A_DOUT(17) => nc117, A_DOUT(16) => \readData5[16]\, 
        A_DOUT(15) => \readData5[15]\, A_DOUT(14) => 
        \readData5[14]\, A_DOUT(13) => \readData5[13]\, 
        A_DOUT(12) => \readData5[12]\, A_DOUT(11) => 
        \readData5[11]\, A_DOUT(10) => \readData5[10]\, A_DOUT(9)
         => \readData5[9]\, A_DOUT(8) => nc36, A_DOUT(7) => 
        \readData5[7]\, A_DOUT(6) => \readData5[6]\, A_DOUT(5)
         => \readData5[5]\, A_DOUT(4) => \readData5[4]\, 
        A_DOUT(3) => \readData5[3]\, A_DOUT(2) => \readData5[2]\, 
        A_DOUT(1) => \readData5[1]\, A_DOUT(0) => \readData5[0]\, 
        B_DOUT(17) => nc116, B_DOUT(16) => \readData5[34]\, 
        B_DOUT(15) => \readData5[33]\, B_DOUT(14) => 
        \readData5[32]\, B_DOUT(13) => \readData5[31]\, 
        B_DOUT(12) => \readData5[30]\, B_DOUT(11) => 
        \readData5[29]\, B_DOUT(10) => \readData5[28]\, B_DOUT(9)
         => \readData5[27]\, B_DOUT(8) => nc48, B_DOUT(7) => 
        \readData5[25]\, B_DOUT(6) => \readData5[24]\, B_DOUT(5)
         => \readData5[23]\, B_DOUT(4) => \readData5[22]\, 
        B_DOUT(3) => \readData5[21]\, B_DOUT(2) => 
        \readData5[20]\, B_DOUT(1) => \readData5[19]\, B_DOUT(0)
         => \readData5[18]\, BUSY => OPEN, A_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => N_375_i_0, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        N_72_i_0, A_DIN(15) => N_70_i_0, A_DIN(14) => N_68_i_0, 
        A_DIN(13) => N_66_i_0, A_DIN(12) => N_64_i_0, A_DIN(11)
         => N_58_i_0, A_DIN(10) => N_56_i_0, A_DIN(9) => N_54_i_0, 
        A_DIN(8) => GND_net_1, A_DIN(7) => N_52_i_0, A_DIN(6) => 
        N_50_i_0, A_DIN(5) => N_48_i_0, A_DIN(4) => N_46_i_0, 
        A_DIN(3) => N_44_i_0, A_DIN(2) => N_42_i_0, A_DIN(1) => 
        N_40_i_0, A_DIN(0) => N_38_i_0, A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a5_1[1]\, 
        A_WEN(0) => \wen_a5_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b5_1[1]\, 
        B_WEN(0) => \wen_b5_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block31_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem_m3(3), Y => \wen_b31_1[1]\);
    
    \readData_31_am_RNO_0[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[30]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[27]\, D => \readData10[30]\, Y => 
        N_397);
    
    readdata_xhdl1418_0_a2_0_0 : CFG3
      generic map(INIT => x"01")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => readdata_xhdl1419_0_a2_0);
    
    \readData_31_am_RNO_2[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[12]\, D => \readData2[12]\, Y => 
        \readData_10_1_1[11]\);
    
    \readData_31_ns[12]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[12]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[12]_net_1\, Y => 
        ram_rdata(12));
    
    \readData_31_bm_RNO_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[12]\, D => \readData7[12]\, Y => 
        \readData_28_1_1[11]\);
    
    \readData_31_bm_1_1_RNO[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[18]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[16]\, D => \readData13[18]\, Y => 
        N_738);
    
    \readData_31_am_RNO_0[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[16]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[15]\, D => \readData10[16]\, Y => 
        N_385);
    
    block25_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem_m3(2), Y => \wen_b25_1[0]\);
    
    \readData_31_bm_RNO_0[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[10]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[9]\, D => \readData11[10]\, Y => 
        N_859);
    
    \readData_31_bm_1_1_RNO_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[0]\, D => \readData5[0]\, Y => 
        \readData_21_1_1[0]\);
    
    \readData_31_am_RNO_0[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[31]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[28]\, D => \readData10[31]\, Y => 
        N_398);
    
    \readData_31_bm_1_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_751, D => N_655, Y => 
        \readData_31_bm_1_1[29]_net_1\);
    
    \readData_31_am_RNO_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[12]\, D => \readData6[12]\, Y => 
        \readData_13_1_1[11]\);
    
    \readData_31_bm_RNO_0[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[3]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[3]\, D => \readData11[3]\, Y => N_853);
    
    \readData_31_am_1_1_RNO_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[25]\, D => \readData4[25]\, Y => 
        \readData_6_1_1[23]\);
    
    \readData_31_am_RNO_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[1]\, D => \readData6[1]\, Y => 
        \readData_13_1_1[1]\);
    
    \readData_31_bm_1_1_RNO_0[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[25]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[23]\, D => \readData9[25]\, Y => 
        N_649);
    
    \readData_31_bm_1_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_743, D => N_647, Y => 
        \readData_31_bm_1_1[21]_net_1\);
    
    \readData_31_am_1_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_268, D => N_172, Y => 
        \readData_31_am_1_1[26]_net_1\);
    
    \readData_31_ns[21]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[21]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[21]_net_1\, Y => 
        ram_rdata(21));
    
    \readData_31_am_1_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_260, D => N_164, Y => 
        \readData_31_am_1_1[18]_net_1\);
    
    block29_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem_m3(3), Y => \wen_b29_1[1]\);
    
    \readData_31_am_RNO_2[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[19]\, D => \readData2[19]\, Y => 
        \readData_10_1_1[17]\);
    
    \readData_31_bm_1_1_RNO[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[7]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[7]\, D => \readData13[7]\, Y => N_729);
    
    block1_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem_m3(3), Y
         => \wen_b1_1[1]\);
    
    \readData_31_am_1_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_248, D => N_152, Y => \readData_31_am_1_1[6]_net_1\);
    
    \readData_31_bm_RNO_0[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[19]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[17]\, D => \readData11[19]\, Y => 
        N_867);
    
    \readData_31_am_RNO[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[14]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[13]\, D => \readData14[14]\, Y => 
        N_479);
    
    \readData_31_am_RNO_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[19]\, D => \readData6[19]\, Y => 
        \readData_13_1_1[17]\);
    
    \readData_31_am_RNO_2[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[20]\, D => \readData2[20]\, Y => 
        \readData_10_1_1[18]\);
    
    \readData_31_am_1_1_RNO_2[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[12]\, D => \readData0[12]\, Y => 
        \readData_3_1_1[11]\);
    
    \readData_31_am_RNO_2[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[28]\, D => \readData2[28]\, Y => 
        \readData_10_1_1[25]\);
    
    block11_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(1), Y => \wen_a11_1[1]\);
    
    \readData_31_bm_1_1_RNO_2[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[11]\, D => \readData1[11]\, Y => 
        \readData_18_1_1[10]\);
    
    \readData_31_bm_RNO_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[7]\, D => \readData7[7]\, Y => 
        \readData_28_1_1[7]\);
    
    \readData_31_am_1_1_RNO_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[12]\, D => \readData4[12]\, Y => 
        \readData_6_1_1[11]\);
    
    \readData_31_am_1_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_264, D => N_168, Y => 
        \readData_31_am_1_1[22]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[9]\, D => \readData5[9]\, Y => 
        \readData_21_1_1[8]\);
    
    \readData_31_bm_1_1_RNO[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[29]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[26]\, D => \readData13[29]\, Y => 
        N_748);
    
    block7_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(0), Y => \wen_a7_1[0]\);
    
    \readData_31_am_RNO_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[20]\, D => \readData6[20]\, Y => 
        \readData_13_1_1[18]\);
    
    \readData_31_am_1_1_RNO_0[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[32]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[29]\, D => \readData8[32]\, Y => 
        N_175);
    
    \readData_31_bm_1_1_RNO_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[11]\, D => \readData5[11]\, Y => 
        \readData_21_1_1[10]\);
    
    \readData_31_bm[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_964, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[18]_net_1\, D => N_868, Y => 
        \readData_31_bm[18]_net_1\);
    
    \readData_31_bm_RNO[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[27]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[24]\, D => \readData15[27]\, Y => 
        N_970);
    
    \readData_31_am_RNO_2[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[10]\, D => \readData2[10]\, Y => 
        \readData_10_1_1[9]\);
    
    \readData_31_bm_1_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_753, D => N_657, Y => 
        \readData_31_bm_1_1[31]_net_1\);
    
    block23_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(0), Y => \wen_a23_1[0]\);
    
    \readData_31_am_1_1_RNO[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[0]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[0]\, D => \readData12[0]\, Y => N_242);
    
    \readData_31_bm_1_1_RNO_0[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[32]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[29]\, D => \readData9[32]\, Y => 
        N_655);
    
    \readData_31_bm_1_1_RNO_2[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[25]\, D => \readData1[25]\, Y => 
        \readData_18_1_1[23]\);
    
    \readData_31_am[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_483, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[17]_net_1\, D => N_387, Y => 
        \readData_31_am[17]_net_1\);
    
    \readData_31_bm_RNO_0[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[13]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[12]\, D => \readData11[13]\, Y => 
        N_862);
    
    \readData_31_bm_1_1_RNO_2[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[12]\, D => \readData1[12]\, Y => 
        \readData_18_1_1[11]\);
    
    \readData_31_bm_1_1_RNO_0[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[4]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[4]\, D => \readData9[4]\, Y => N_630);
    
    block15_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(0), Y => \wen_a15_1[0]\);
    
    block12_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(0), Y => \wen_a12_1[0]\);
    
    \readData_31_bm_RNO_2[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[30]\, D => \readData3[30]\, Y => 
        \readData_25_1_1[27]\);
    
    \readData_31_am_RNO[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[31]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[28]\, D => \readData14[31]\, Y => 
        N_494);
    
    block11_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem_m3(3), Y => \wen_b11_1[1]\);
    
    \readData_31_bm_1_1_RNO_2[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[19]\, D => \readData1[19]\, Y => 
        \readData_18_1_1[17]\);
    
    block20_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem_m3(2), Y => \wen_b20_1[0]\);
    
    \readData_31_bm_1_1_RNO_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[12]\, D => \readData5[12]\, Y => 
        \readData_21_1_1[11]\);
    
    \readData_31_am_RNO_0[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[13]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[12]\, D => \readData10[13]\, Y => 
        N_382);
    
    \readData_31_ns[15]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[15]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[15]_net_1\, Y => 
        ram_rdata(15));
    
    \readData_31_bm[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_966, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[20]_net_1\, D => N_870, Y => 
        \readData_31_bm[20]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[19]\, D => \readData5[19]\, Y => 
        \readData_21_1_1[17]\);
    
    \readData_31_am_RNO[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[33]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[30]\, D => \readData14[33]\, Y => 
        N_496);
    
    \readData_31_am_RNO_2[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[3]\, D => \readData2[3]\, Y => 
        \readData_10_1_1[3]\);
    
    \readData_31_bm_RNO_0[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[0]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[0]\, D => \readData11[0]\, Y => N_850);
    
    \readData_31_am_RNO[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[15]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[14]\, D => \readData14[15]\, Y => 
        N_480);
    
    \readData_31_am_1_1_RNO_2[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[3]\, D => \readData0[3]\, Y => 
        \readData_3_1_1[3]\);
    
    \readData_31_am[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_470, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[4]_net_1\, D => N_374, Y => 
        \readData_31_am[4]_net_1\);
    
    block30_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(0), Y => \wen_a30_1[0]\);
    
    \readData_31_am_1_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_271, D => N_175, Y => 
        \readData_31_am_1_1[29]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[18]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[16]\, D => \readData9[18]\, Y => 
        N_642);
    
    block20 : RAM1K18
      port map(A_DOUT(17) => nc37, A_DOUT(16) => \readData20[16]\, 
        A_DOUT(15) => \readData20[15]\, A_DOUT(14) => 
        \readData20[14]\, A_DOUT(13) => \readData20[13]\, 
        A_DOUT(12) => \readData20[12]\, A_DOUT(11) => 
        \readData20[11]\, A_DOUT(10) => \readData20[10]\, 
        A_DOUT(9) => \readData20[9]\, A_DOUT(8) => nc5, A_DOUT(7)
         => \readData20[7]\, A_DOUT(6) => \readData20[6]\, 
        A_DOUT(5) => \readData20[5]\, A_DOUT(4) => 
        \readData20[4]\, A_DOUT(3) => \readData20[3]\, A_DOUT(2)
         => \readData20[2]\, A_DOUT(1) => \readData20[1]\, 
        A_DOUT(0) => \readData20[0]\, B_DOUT(17) => nc103, 
        B_DOUT(16) => \readData20[34]\, B_DOUT(15) => 
        \readData20[33]\, B_DOUT(14) => \readData20[32]\, 
        B_DOUT(13) => \readData20[31]\, B_DOUT(12) => 
        \readData20[30]\, B_DOUT(11) => \readData20[29]\, 
        B_DOUT(10) => \readData20[28]\, B_DOUT(9) => 
        \readData20[27]\, B_DOUT(8) => nc101, B_DOUT(7) => 
        \readData20[25]\, B_DOUT(6) => \readData20[24]\, 
        B_DOUT(5) => \readData20[23]\, B_DOUT(4) => 
        \readData20[22]\, B_DOUT(3) => \readData20[21]\, 
        B_DOUT(2) => \readData20[20]\, B_DOUT(1) => 
        \readData20[19]\, B_DOUT(0) => \readData20[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a20_1[1]\, A_WEN(0) => \wen_a20_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b20_1[1]\, 
        B_WEN(0) => \wen_b20_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_1_1_RNO_2[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[32]\, D => \readData0[32]\, Y => 
        \readData_3_1_1[29]\);
    
    \readData_31_bm_1_1_RNO_0[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[9]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[8]\, D => \readData9[9]\, Y => N_634);
    
    \readData_31_bm_RNO_2[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[24]\, D => \readData3[24]\, Y => 
        \readData_25_1_1[22]\);
    
    \readData_31_bm_1_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_730, D => N_634, Y => \readData_31_bm_1_1[8]_net_1\);
    
    \readData_31_bm_1_1_RNO[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[16]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[15]\, D => \readData13[16]\, Y => 
        N_737);
    
    \readData_31_bm_1_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_732, D => N_636, Y => 
        \readData_31_bm_1_1[10]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[32]\, D => \readData1[32]\, Y => 
        \readData_18_1_1[29]\);
    
    \readData_31_am_1_1_RNO_2[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[10]\, D => \readData0[10]\, Y => 
        \readData_3_1_1[9]\);
    
    \readData_31_am_RNO[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[19]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[17]\, D => \readData14[19]\, Y => 
        N_483);
    
    \readData_31_bm_1_1_RNO_2[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[4]\, D => \readData1[4]\, Y => 
        \readData_18_1_1[4]\);
    
    \readData_31_am_RNO_2[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[7]\, D => \readData2[7]\, Y => 
        \readData_10_1_1[7]\);
    
    \readData_31_am_RNO_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[29]\, D => \readData6[29]\, Y => 
        \readData_13_1_1[26]\);
    
    \readData_31_am_RNO_2[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[24]\, D => \readData2[24]\, Y => 
        \readData_10_1_1[22]\);
    
    \readData_31_am_1_1_RNO_0[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[13]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[12]\, D => \readData8[13]\, Y => 
        N_158);
    
    \readData_31_bm_RNO[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[30]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[27]\, D => \readData15[30]\, Y => 
        N_973);
    
    \readData_31_bm_1_1_RNO[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[12]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[11]\, D => \readData13[12]\, Y => 
        N_733);
    
    \readData_31_am[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_475, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[9]_net_1\, D => N_379, Y => 
        \readData_31_am[9]_net_1\);
    
    \readData_31_am_RNO[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[1]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[1]\, D => \readData14[1]\, Y => N_467);
    
    \readData_31_am_RNO[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[4]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[4]\, D => \readData14[4]\, Y => N_470);
    
    block22_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(1), Y => \wen_a_m[1]\);
    
    \readData_31_am_RNO_0[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[22]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[20]\, D => \readData10[22]\, Y => 
        N_390);
    
    \readData_31_am_RNO[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[18]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[16]\, D => \readData14[18]\, Y => 
        N_482);
    
    \readData_31_ns[27]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[27]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[27]_net_1\, Y => 
        ram_rdata(27));
    
    \readData_31_am_RNO[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[23]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[21]\, D => \readData14[23]\, Y => 
        N_487);
    
    \readData_31_bm_1_1_RNO_0[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[13]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[12]\, D => \readData9[13]\, Y => 
        N_638);
    
    block0_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem_m3(3), Y
         => \wen_b0_1[1]\);
    
    \readData_31_bm_RNO_0[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[6]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[6]\, D => \readData11[6]\, Y => N_856);
    
    \readData_31_bm[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_947, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[1]_net_1\, D => N_851, Y => 
        \readData_31_bm[1]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[1]\, D => \readData1[1]\, Y => 
        \readData_18_1_1[1]\);
    
    \readData_31_bm[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_952, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[6]_net_1\, D => N_856, Y => 
        \readData_31_bm[6]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[10]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[9]\, D => \readData9[10]\, Y => 
        N_635);
    
    \readData_31_bm_RNO[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[2]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[2]\, D => \readData15[2]\, Y => N_948);
    
    block5_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem_m3(3), Y => 
        \wen_b5_1[1]\);
    
    block10_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(0), Y => \wen_a10_1[0]\);
    
    \readData_31_bm_RNO[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[31]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[28]\, D => \readData15[31]\, Y => 
        N_974);
    
    \readData_31_bm[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_949, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[3]_net_1\, D => N_853, Y => 
        \readData_31_bm[3]_net_1\);
    
    \readData_31_am_RNO_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[32]\, D => \readData6[32]\, Y => 
        \readData_13_1_1[29]\);
    
    block18_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(14), C
         => readdata_xhdl1401_1, D => sram_wen_mem_m3(3), Y => 
        \wen_b18_1[1]\);
    
    \readData_31_am_1_1_RNO_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[6]\, D => \readData4[6]\, Y => 
        \readData_6_1_1[6]\);
    
    \readData_31_am_RNO[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[3]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[3]\, D => \readData14[3]\, Y => N_469);
    
    block14_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem(0), Y => \wen_a14_1[0]\);
    
    \readData_31_am_RNO_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[27]\, D => \readData6[27]\, Y => 
        \readData_13_1_1[24]\);
    
    \readData_31_bm_1_1_RNO[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[28]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[25]\, D => \readData13[28]\, Y => 
        N_747);
    
    \readData_31_am_RNO_2[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[11]\, D => \readData2[11]\, Y => 
        \readData_10_1_1[10]\);
    
    block0_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem_m3(2), Y
         => \wen_b0_1[0]\);
    
    \readData_31_bm_1_1_RNO_0[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[1]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[1]\, D => \readData9[1]\, Y => N_627);
    
    \readData_31_am_1_1_RNO_0[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[5]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[5]\, D => \readData8[5]\, Y => N_151);
    
    block28_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem_m3(2), Y => \wen_b28_1[0]\);
    
    \readData_31_bm_1_1_RNO_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[25]\, D => \readData5[25]\, Y => 
        \readData_21_1_1[23]\);
    
    \readData_31_bm_RNO[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[12]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[11]\, D => \readData15[12]\, Y => 
        N_957);
    
    \readData_31_bm_RNO_2[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[4]\, D => \readData3[4]\, Y => 
        \readData_25_1_1[4]\);
    
    \readData_31_bm[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_963, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[17]_net_1\, D => N_867, Y => 
        \readData_31_bm[17]_net_1\);
    
    \readData_31_am_RNO_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[11]\, D => \readData6[11]\, Y => 
        \readData_13_1_1[10]\);
    
    \readData_31_bm_1_1_RNO[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[23]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[21]\, D => \readData13[23]\, Y => 
        N_743);
    
    \readData_31_bm_1_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_724, D => N_628, Y => \readData_31_bm_1_1[2]_net_1\);
    
    \readData_31_am_1_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_267, D => N_171, Y => 
        \readData_31_am_1_1[25]_net_1\);
    
    \readData_31_bm_RNO_2[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[6]\, D => \readData3[6]\, Y => 
        \readData_25_1_1[6]\);
    
    \readData_31_bm_RNO_2[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[33]\, D => \readData3[33]\, Y => 
        \readData_25_1_1[30]\);
    
    \readData_31_ns[30]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[30]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[30]_net_1\, Y => 
        ram_rdata(30));
    
    \readData_31_am_1_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_251, D => N_155, Y => \readData_31_am_1_1[9]_net_1\);
    
    \readData_31_am_1_1_RNO_0[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[18]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[16]\, D => \readData8[18]\, Y => 
        N_162);
    
    \readData_31_am_RNO_0[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[25]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[23]\, D => \readData10[25]\, Y => 
        N_393);
    
    \readData_31_am_1_1_RNO_0[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[30]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[27]\, D => \readData8[30]\, Y => 
        N_173);
    
    \readData_31_bm_RNO[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[18]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[16]\, D => \readData15[18]\, Y => 
        N_962);
    
    \readData_31_am_1_1_RNO_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[32]\, D => \readData4[32]\, Y => 
        \readData_6_1_1[29]\);
    
    \readData_31_bm_1_1_RNO_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[3]\, D => \readData5[3]\, Y => 
        \readData_21_1_1[3]\);
    
    \readData_31_bm_RNO[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[11]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[10]\, D => \readData15[11]\, Y => 
        N_956);
    
    \readData_31_bm[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_961, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[15]_net_1\, D => N_865, Y => 
        \readData_31_bm[15]_net_1\);
    
    \readData_31_am_1_1[11]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_253, D => N_157, Y => 
        \readData_31_am_1_1[11]_net_1\);
    
    block16_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem_m3(3), Y => 
        \wen_b16_1[1]\);
    
    block13_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem_m3(3), Y => 
        \wen_b13_1[1]\);
    
    \readData_31_bm_RNO_0[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[1]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[1]\, D => \readData11[1]\, Y => N_851);
    
    \readData_31_bm_1_1_RNO_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[32]\, D => \readData5[32]\, Y => 
        \readData_21_1_1[29]\);
    
    \readData_31_am_RNO_0[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[9]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[8]\, D => \readData10[9]\, Y => N_378);
    
    \readData_31_am_RNO_2[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[14]\, D => \readData2[14]\, Y => 
        \readData_10_1_1[13]\);
    
    \readData_31_bm_1_1_RNO_2[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[18]\, D => \readData1[18]\, Y => 
        \readData_18_1_1[16]\);
    
    block27 : RAM1K18
      port map(A_DOUT(17) => nc52, A_DOUT(16) => \readData27[16]\, 
        A_DOUT(15) => \readData27[15]\, A_DOUT(14) => 
        \readData27[14]\, A_DOUT(13) => \readData27[13]\, 
        A_DOUT(12) => \readData27[12]\, A_DOUT(11) => 
        \readData27[11]\, A_DOUT(10) => \readData27[10]\, 
        A_DOUT(9) => \readData27[9]\, A_DOUT(8) => nc76, 
        A_DOUT(7) => \readData27[7]\, A_DOUT(6) => 
        \readData27[6]\, A_DOUT(5) => \readData27[5]\, A_DOUT(4)
         => \readData27[4]\, A_DOUT(3) => \readData27[3]\, 
        A_DOUT(2) => \readData27[2]\, A_DOUT(1) => 
        \readData27[1]\, A_DOUT(0) => \readData27[0]\, B_DOUT(17)
         => nc51, B_DOUT(16) => \readData27[34]\, B_DOUT(15) => 
        \readData27[33]\, B_DOUT(14) => \readData27[32]\, 
        B_DOUT(13) => \readData27[31]\, B_DOUT(12) => 
        \readData27[30]\, B_DOUT(11) => \readData27[29]\, 
        B_DOUT(10) => \readData27[28]\, B_DOUT(9) => 
        \readData27[27]\, B_DOUT(8) => nc66, B_DOUT(7) => 
        \readData27[25]\, B_DOUT(6) => \readData27[24]\, 
        B_DOUT(5) => \readData27[23]\, B_DOUT(4) => 
        \readData27[22]\, B_DOUT(3) => \readData27[21]\, 
        B_DOUT(2) => \readData27[20]\, B_DOUT(1) => 
        \readData27[19]\, B_DOUT(0) => \readData27[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a27_1[1]\, A_WEN(0) => \wen_a27_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b27_1[1]\, 
        B_WEN(0) => \wen_b27_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block25_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(0), Y => \wen_a25_1[0]\);
    
    block22_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(0), Y => \wen_a_m[0]\);
    
    \readData_31_bm_RNO_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[29]\, D => \readData7[29]\, Y => 
        \readData_28_1_1[26]\);
    
    \readData_31_bm_1_1_RNO_0[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[31]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[28]\, D => \readData9[31]\, Y => 
        N_654);
    
    \readData_31_bm_RNO_0[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[27]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[24]\, D => \readData11[27]\, Y => 
        N_874);
    
    \readData_31_bm_1_1_RNO_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[18]\, D => \readData5[18]\, Y => 
        \readData_21_1_1[16]\);
    
    \readData_31_am_RNO_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[14]\, D => \readData6[14]\, Y => 
        \readData_13_1_1[13]\);
    
    \readData_31_am_1_1_RNO[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[33]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[30]\, D => \readData12[33]\, Y => 
        N_272);
    
    block13_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(1), Y => 
        \wen_a13_1[1]\);
    
    \readData_31_bm_RNO_1[29]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[32]\, D => \readData7[32]\, Y => 
        \readData_28_1_1[29]\);
    
    \readData_31_am_1_1_RNO_2[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[30]\, D => \readData0[30]\, Y => 
        \readData_3_1_1[27]\);
    
    block27_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(1), Y => \wen_a27_1[1]\);
    
    \readData_31_am_1_1_RNO_2[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[13]\, D => \readData0[13]\, Y => 
        \readData_3_1_1[12]\);
    
    \readData_31_ns[18]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[18]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[18]_net_1\, Y => 
        ram_rdata(18));
    
    \readData_31_bm_RNO_0[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[12]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[11]\, D => \readData11[12]\, Y => 
        N_861);
    
    \readData_31_bm_RNO[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[7]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[7]\, D => \readData15[7]\, Y => N_953);
    
    \readData_31_ns[19]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[19]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[19]_net_1\, Y => 
        ram_rdata(19));
    
    \readData_31_am_1_1_RNO_2[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[2]\, D => \readData0[2]\, Y => 
        \readData_3_1_1[2]\);
    
    \readData_31_am_1_1_RNO_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[13]\, D => \readData4[13]\, Y => 
        \readData_6_1_1[12]\);
    
    \readData_31_bm_1_1_RNO_2[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[13]\, D => \readData1[13]\, Y => 
        \readData_18_1_1[12]\);
    
    \readData_31_am_RNO_0[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[12]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[11]\, D => \readData10[12]\, Y => 
        N_381);
    
    \readData_31_bm_RNO_2[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[15]\, D => \readData3[15]\, Y => 
        \readData_25_1_1[14]\);
    
    \readData_31_bm[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_950, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[4]_net_1\, D => N_854, Y => 
        \readData_31_bm[4]_net_1\);
    
    \readData_31_bm_1_1_RNO_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[13]\, D => \readData5[13]\, Y => 
        \readData_21_1_1[12]\);
    
    block30 : RAM1K18
      port map(A_DOUT(17) => nc77, A_DOUT(16) => \readData30[16]\, 
        A_DOUT(15) => \readData30[15]\, A_DOUT(14) => 
        \readData30[14]\, A_DOUT(13) => \readData30[13]\, 
        A_DOUT(12) => \readData30[12]\, A_DOUT(11) => 
        \readData30[11]\, A_DOUT(10) => \readData30[10]\, 
        A_DOUT(9) => \readData30[9]\, A_DOUT(8) => nc67, 
        A_DOUT(7) => \readData30[7]\, A_DOUT(6) => 
        \readData30[6]\, A_DOUT(5) => \readData30[5]\, A_DOUT(4)
         => \readData30[4]\, A_DOUT(3) => \readData30[3]\, 
        A_DOUT(2) => \readData30[2]\, A_DOUT(1) => 
        \readData30[1]\, A_DOUT(0) => \readData30[0]\, B_DOUT(17)
         => nc4, B_DOUT(16) => \readData30[34]\, B_DOUT(15) => 
        \readData30[33]\, B_DOUT(14) => \readData30[32]\, 
        B_DOUT(13) => \readData30[31]\, B_DOUT(12) => 
        \readData30[30]\, B_DOUT(11) => \readData30[29]\, 
        B_DOUT(10) => \readData30[28]\, B_DOUT(9) => 
        \readData30[27]\, B_DOUT(8) => nc124, B_DOUT(7) => 
        \readData30[25]\, B_DOUT(6) => \readData30[24]\, 
        B_DOUT(5) => \readData30[23]\, B_DOUT(4) => 
        \readData30[22]\, B_DOUT(3) => \readData30[21]\, 
        B_DOUT(2) => \readData30[20]\, B_DOUT(1) => 
        \readData30[19]\, B_DOUT(0) => \readData30[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a30_1[1]\, A_WEN(0) => \wen_a30_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b30_1[1]\, 
        B_WEN(0) => \wen_b30_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_RNO_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[2]\, D => \readData6[2]\, Y => 
        \readData_13_1_1[2]\);
    
    \readData_31_bm_RNO_2[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[5]\, D => \readData3[5]\, Y => 
        \readData_25_1_1[5]\);
    
    block8_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem_m3(3), Y => \wen_b8_1[1]\);
    
    \readData_31_bm_RNO_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[15]\, D => \readData7[15]\, Y => 
        \readData_28_1_1[14]\);
    
    \readData_31_bm_1_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_726, D => N_630, Y => \readData_31_bm_1_1[4]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[15]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[14]\, D => \readData9[15]\, Y => 
        N_640);
    
    \readData_31_bm_1_1_RNO_2[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[31]\, D => \readData1[31]\, Y => 
        \readData_18_1_1[28]\);
    
    \readData_31_am_1_1_RNO_2[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[6]\, D => \readData0[6]\, Y => 
        \readData_3_1_1[6]\);
    
    \readData_31_bm_RNO_0[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[4]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[4]\, D => \readData11[4]\, Y => N_854);
    
    \readData_31_bm_RNO[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[25]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[23]\, D => \readData15[25]\, Y => 
        N_969);
    
    \readData_31_am_1_1_RNO[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[7]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[7]\, D => \readData12[7]\, Y => N_249);
    
    \readData_31_ns[23]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[23]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[23]_net_1\, Y => 
        ram_rdata(23));
    
    \readData_31_am_1_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_255, D => N_159, Y => 
        \readData_31_am_1_1[13]_net_1\);
    
    block31_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem_m3(2), Y => \wen_b31_1[0]\);
    
    block29_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(1), Y => \wen_a29_1[1]\);
    
    \readData_31_bm[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_955, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[9]_net_1\, D => N_859, Y => 
        \readData_31_bm[9]_net_1\);
    
    \readData_31_bm_RNO_2[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[23]\, D => \readData3[23]\, Y => 
        \readData_25_1_1[21]\);
    
    \readData_31_am_RNO_0[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[19]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[17]\, D => \readData10[19]\, Y => 
        N_387);
    
    \readData_31_bm_RNO_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[25]\, D => \readData7[25]\, Y => 
        \readData_28_1_1[23]\);
    
    block4 : RAM1K18
      port map(A_DOUT(17) => nc109, A_DOUT(16) => \readData4[16]\, 
        A_DOUT(15) => \readData4[15]\, A_DOUT(14) => 
        \readData4[14]\, A_DOUT(13) => \readData4[13]\, 
        A_DOUT(12) => \readData4[12]\, A_DOUT(11) => 
        \readData4[11]\, A_DOUT(10) => \readData4[10]\, A_DOUT(9)
         => \readData4[9]\, A_DOUT(8) => nc42, A_DOUT(7) => 
        \readData4[7]\, A_DOUT(6) => \readData4[6]\, A_DOUT(5)
         => \readData4[5]\, A_DOUT(4) => \readData4[4]\, 
        A_DOUT(3) => \readData4[3]\, A_DOUT(2) => \readData4[2]\, 
        A_DOUT(1) => \readData4[1]\, A_DOUT(0) => \readData4[0]\, 
        B_DOUT(17) => nc114, B_DOUT(16) => \readData4[34]\, 
        B_DOUT(15) => \readData4[33]\, B_DOUT(14) => 
        \readData4[32]\, B_DOUT(13) => \readData4[31]\, 
        B_DOUT(12) => \readData4[30]\, B_DOUT(11) => 
        \readData4[29]\, B_DOUT(10) => \readData4[28]\, B_DOUT(9)
         => \readData4[27]\, B_DOUT(8) => nc100, B_DOUT(7) => 
        \readData4[25]\, B_DOUT(6) => \readData4[24]\, B_DOUT(5)
         => \readData4[23]\, B_DOUT(4) => \readData4[22]\, 
        B_DOUT(3) => \readData4[21]\, B_DOUT(2) => 
        \readData4[20]\, B_DOUT(1) => \readData4[19]\, B_DOUT(0)
         => \readData4[18]\, BUSY => OPEN, A_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => N_375_i_0, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        N_72_i_0, A_DIN(15) => N_70_i_0, A_DIN(14) => N_68_i_0, 
        A_DIN(13) => N_66_i_0, A_DIN(12) => N_64_i_0, A_DIN(11)
         => N_58_i_0, A_DIN(10) => N_56_i_0, A_DIN(9) => N_54_i_0, 
        A_DIN(8) => GND_net_1, A_DIN(7) => N_52_i_0, A_DIN(6) => 
        N_50_i_0, A_DIN(5) => N_48_i_0, A_DIN(4) => N_46_i_0, 
        A_DIN(3) => N_44_i_0, A_DIN(2) => N_42_i_0, A_DIN(1) => 
        N_40_i_0, A_DIN(0) => N_38_i_0, A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a4_1[1]\, 
        A_WEN(0) => \wen_a4_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b4_1[1]\, 
        B_WEN(0) => \wen_b4_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block20_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(0), Y => \wen_a20_1[0]\);
    
    \readData_31_am_RNO_2[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[23]\, D => \readData2[23]\, Y => 
        \readData_10_1_1[21]\);
    
    \readData_31_bm_RNO_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[22]\, D => \readData7[22]\, Y => 
        \readData_28_1_1[20]\);
    
    \readData_31_am_1_1_RNO_2[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[7]\, D => \readData0[7]\, Y => 
        \readData_3_1_1[7]\);
    
    \readData_31_am_RNO_0[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[20]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[18]\, D => \readData10[20]\, Y => 
        N_388);
    
    \readData_31_am_1_1_RNO_0[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[11]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[10]\, D => \readData8[11]\, Y => 
        N_156);
    
    \wen_a_m_30_0_a2_0[1]\ : CFG3
      generic map(INIT => x"20")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1144);
    
    block24_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(0), Y => \wen_a24_1[0]\);
    
    \readData_31_am_1_1_RNO_2[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[18]\, D => \readData0[18]\, Y => 
        \readData_3_1_1[16]\);
    
    \readData_31_am_1_1_RNO[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[20]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[18]\, D => \readData12[20]\, Y => 
        N_260);
    
    \readData_31_bm_1_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_739, D => N_643, Y => 
        \readData_31_bm_1_1[17]_net_1\);
    
    \readData_31_am_RNO[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[21]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[19]\, D => \readData14[21]\, Y => 
        N_485);
    
    \readData_31_am_1_1_RNO_2[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[34]\, D => \readData0[34]\, Y => 
        \readData_3_1_1[31]\);
    
    \readData_31_am_1_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_270, D => N_174, Y => 
        \readData_31_am_1_1[28]_net_1\);
    
    \readData_31_am_1_1_RNO_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[18]\, D => \readData4[18]\, Y => 
        \readData_6_1_1[16]\);
    
    block27_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem_m3(3), Y => \wen_b27_1[1]\);
    
    \readData_31_am_1_1_RNO_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[34]\, D => \readData4[34]\, Y => 
        \readData_6_1_1[31]\);
    
    \readData_31_bm_1_1_RNO_2[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[33]\, D => \readData1[33]\, Y => 
        \readData_18_1_1[30]\);
    
    \readData_31_bm_1_1_RNO_0[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[28]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[25]\, D => \readData9[28]\, Y => 
        N_651);
    
    block1 : RAM1K18
      port map(A_DOUT(17) => nc83, A_DOUT(16) => \readData1[16]\, 
        A_DOUT(15) => \readData1[15]\, A_DOUT(14) => 
        \readData1[14]\, A_DOUT(13) => \readData1[13]\, 
        A_DOUT(12) => \readData1[12]\, A_DOUT(11) => 
        \readData1[11]\, A_DOUT(10) => \readData1[10]\, A_DOUT(9)
         => \readData1[9]\, A_DOUT(8) => nc41, A_DOUT(7) => 
        \readData1[7]\, A_DOUT(6) => \readData1[6]\, A_DOUT(5)
         => \readData1[5]\, A_DOUT(4) => \readData1[4]\, 
        A_DOUT(3) => \readData1[3]\, A_DOUT(2) => \readData1[2]\, 
        A_DOUT(1) => \readData1[1]\, A_DOUT(0) => \readData1[0]\, 
        B_DOUT(17) => nc90, B_DOUT(16) => \readData1[34]\, 
        B_DOUT(15) => \readData1[33]\, B_DOUT(14) => 
        \readData1[32]\, B_DOUT(13) => \readData1[31]\, 
        B_DOUT(12) => \readData1[30]\, B_DOUT(11) => 
        \readData1[29]\, B_DOUT(10) => \readData1[28]\, B_DOUT(9)
         => \readData1[27]\, B_DOUT(8) => nc94, B_DOUT(7) => 
        \readData1[25]\, B_DOUT(6) => \readData1[24]\, B_DOUT(5)
         => \readData1[23]\, B_DOUT(4) => \readData1[22]\, 
        B_DOUT(3) => \readData1[21]\, B_DOUT(2) => 
        \readData1[20]\, B_DOUT(1) => \readData1[19]\, B_DOUT(0)
         => \readData1[18]\, BUSY => OPEN, A_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => N_375_i_0, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        N_72_i_0, A_DIN(15) => N_70_i_0, A_DIN(14) => N_68_i_0, 
        A_DIN(13) => N_66_i_0, A_DIN(12) => N_64_i_0, A_DIN(11)
         => N_58_i_0, A_DIN(10) => N_56_i_0, A_DIN(9) => N_54_i_0, 
        A_DIN(8) => GND_net_1, A_DIN(7) => N_52_i_0, A_DIN(6) => 
        N_50_i_0, A_DIN(5) => N_48_i_0, A_DIN(4) => N_46_i_0, 
        A_DIN(3) => N_44_i_0, A_DIN(2) => N_42_i_0, A_DIN(1) => 
        N_40_i_0, A_DIN(0) => N_38_i_0, A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a1_1[1]\, 
        A_WEN(0) => \wen_a1_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b1_1[1]\, 
        B_WEN(0) => \wen_b1_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_1_1_RNO_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[33]\, D => \readData5[33]\, Y => 
        \readData_21_1_1[30]\);
    
    block5_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(0), Y => 
        \wen_a5_1[0]\);
    
    \readData_31_bm_1_1_RNO_2[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[3]\, D => \readData1[3]\, Y => 
        \readData_18_1_1[3]\);
    
    \readData_31_am_RNO_2[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[30]\, D => \readData2[30]\, Y => 
        \readData_10_1_1[27]\);
    
    \readData_31_am_1_1_RNO[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[21]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[19]\, D => \readData12[21]\, Y => 
        N_261);
    
    block27_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem_m3(2), Y => \wen_b27_1[0]\);
    
    \readData_31_am_RNO_2[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[31]\, D => \readData2[31]\, Y => 
        \readData_10_1_1[28]\);
    
    \readData_31_am_1_1_RNO_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[30]\, D => \readData4[30]\, Y => 
        \readData_6_1_1[27]\);
    
    readdata_xhdl1400_0_a2_0 : CFG3
      generic map(INIT => x"02")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1168);
    
    \readData_31_bm_1_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_736, D => N_640, Y => 
        \readData_31_bm_1_1[14]_net_1\);
    
    \readData_31_am_RNO_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[5]\, D => \readData6[5]\, Y => 
        \readData_13_1_1[5]\);
    
    block14_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem_m3(2), Y => \wen_b14_1[0]\);
    
    \readData_31_bm_1_1_RNO_2[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[34]\, D => \readData1[34]\, Y => 
        \readData_18_1_1[31]\);
    
    \readData_31_am_1_1_RNO_0[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[0]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[0]\, D => \readData8[0]\, Y => N_146);
    
    \readData_31_am_RNO[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[24]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[22]\, D => \readData14[24]\, Y => 
        N_488);
    
    \readData_31_bm_RNO[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[24]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[22]\, D => \readData15[24]\, Y => 
        N_968);
    
    \readData_31_bm_1_1_RNO_2[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[10]\, D => \readData1[10]\, Y => 
        \readData_18_1_1[9]\);
    
    \readData_31_bm_1_1_RNO[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[11]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[10]\, D => \readData13[11]\, Y => 
        N_732);
    
    \readData_31_bm_1_1_RNO_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[34]\, D => \readData5[34]\, Y => 
        \readData_21_1_1[31]\);
    
    \readData_31_am_RNO[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[2]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[2]\, D => \readData14[2]\, Y => N_468);
    
    block5_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem(1), Y => 
        \wen_a5_1[1]\);
    
    \readData_31_am_1_1_RNO[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[12]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[11]\, D => \readData12[12]\, Y => 
        N_253);
    
    block19 : RAM1K18
      port map(A_DOUT(17) => nc122, A_DOUT(16) => 
        \readData19[16]\, A_DOUT(15) => \readData19[15]\, 
        A_DOUT(14) => \readData19[14]\, A_DOUT(13) => 
        \readData19[13]\, A_DOUT(12) => \readData19[12]\, 
        A_DOUT(11) => \readData19[11]\, A_DOUT(10) => 
        \readData19[10]\, A_DOUT(9) => \readData19[9]\, A_DOUT(8)
         => nc112, A_DOUT(7) => \readData19[7]\, A_DOUT(6) => 
        \readData19[6]\, A_DOUT(5) => \readData19[5]\, A_DOUT(4)
         => \readData19[4]\, A_DOUT(3) => \readData19[3]\, 
        A_DOUT(2) => \readData19[2]\, A_DOUT(1) => 
        \readData19[1]\, A_DOUT(0) => \readData19[0]\, B_DOUT(17)
         => nc86, B_DOUT(16) => \readData19[34]\, B_DOUT(15) => 
        \readData19[33]\, B_DOUT(14) => \readData19[32]\, 
        B_DOUT(13) => \readData19[31]\, B_DOUT(12) => 
        \readData19[30]\, B_DOUT(11) => \readData19[29]\, 
        B_DOUT(10) => \readData19[28]\, B_DOUT(9) => 
        \readData19[27]\, B_DOUT(8) => nc59, B_DOUT(7) => 
        \readData19[25]\, B_DOUT(6) => \readData19[24]\, 
        B_DOUT(5) => \readData19[23]\, B_DOUT(4) => 
        \readData19[22]\, B_DOUT(3) => \readData19[21]\, 
        B_DOUT(2) => \readData19[20]\, B_DOUT(1) => 
        \readData19[19]\, B_DOUT(0) => \readData19[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a19_1[1]\, A_WEN(0) => \wen_a19_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b19_1[1]\, 
        B_WEN(0) => \wen_b19_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    readdata_xhdl1406_1 : CFG3
      generic map(INIT => x"20")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => ahbsram_addr(13), Y => readdata_xhdl1414_1);
    
    \readData_31_am_1_1_RNO[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[31]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[28]\, D => \readData12[31]\, Y => 
        N_270);
    
    \readData_31_ns[11]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[11]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[11]_net_1\, Y => 
        ram_rdata(11));
    
    \readData_31_ns[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[1]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[1]_net_1\, Y => 
        ram_rdata(1));
    
    block0_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem(1), Y => 
        \wen_a0_1[1]\);
    
    \readData_31_bm_RNO_0[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[28]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[25]\, D => \readData11[28]\, Y => 
        N_875);
    
    block11_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem_m3(2), Y => \wen_b11_1[0]\);
    
    \readData_31_ns[20]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[20]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[20]_net_1\, Y => 
        ram_rdata(20));
    
    \readData_31_bm_1_1_RNO[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[20]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[18]\, D => \readData13[20]\, Y => 
        N_740);
    
    \readData_31_ns[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[7]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[7]_net_1\, Y => 
        ram_rdata(7));
    
    \readData_31_bm_1_1_RNO_2[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[28]\, D => \readData1[28]\, Y => 
        \readData_18_1_1[25]\);
    
    \readData_31_bm_1_1_RNO_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[31]\, D => \readData5[31]\, Y => 
        \readData_21_1_1[28]\);
    
    block2_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem_m3(2), Y => \wen_b2_1[0]\);
    
    \readData_31_am_1_1_RNO[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[32]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[29]\, D => \readData12[32]\, Y => 
        N_271);
    
    block5_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => readdata_xhdl1414_1, D => sram_wen_mem_m3(2), Y => 
        \wen_b5_1[0]\);
    
    block14 : RAM1K18
      port map(A_DOUT(17) => nc25, A_DOUT(16) => \readData14[16]\, 
        A_DOUT(15) => \readData14[15]\, A_DOUT(14) => 
        \readData14[14]\, A_DOUT(13) => \readData14[13]\, 
        A_DOUT(12) => \readData14[12]\, A_DOUT(11) => 
        \readData14[11]\, A_DOUT(10) => \readData14[10]\, 
        A_DOUT(9) => \readData14[9]\, A_DOUT(8) => nc15, 
        A_DOUT(7) => \readData14[7]\, A_DOUT(6) => 
        \readData14[6]\, A_DOUT(5) => \readData14[5]\, A_DOUT(4)
         => \readData14[4]\, A_DOUT(3) => \readData14[3]\, 
        A_DOUT(2) => \readData14[2]\, A_DOUT(1) => 
        \readData14[1]\, A_DOUT(0) => \readData14[0]\, B_DOUT(17)
         => nc87, B_DOUT(16) => \readData14[34]\, B_DOUT(15) => 
        \readData14[33]\, B_DOUT(14) => \readData14[32]\, 
        B_DOUT(13) => \readData14[31]\, B_DOUT(12) => 
        \readData14[30]\, B_DOUT(11) => \readData14[29]\, 
        B_DOUT(10) => \readData14[28]\, B_DOUT(9) => 
        \readData14[27]\, B_DOUT(8) => nc35, B_DOUT(7) => 
        \readData14[25]\, B_DOUT(6) => \readData14[24]\, 
        B_DOUT(5) => \readData14[23]\, B_DOUT(4) => 
        \readData14[22]\, B_DOUT(3) => \readData14[21]\, 
        B_DOUT(2) => \readData14[20]\, B_DOUT(1) => 
        \readData14[19]\, B_DOUT(0) => \readData14[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a14_1[1]\, A_WEN(0) => \wen_a14_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b14_1[1]\, 
        B_WEN(0) => \wen_b14_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[6]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[6]\, D => \readData15[6]\, Y => N_952);
    
    \readData_31_ns[9]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[9]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[9]_net_1\, Y => 
        ram_rdata(9));
    
    block12_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem_m3(3), Y => \wen_b12_1[1]\);
    
    \readData_31_bm_1_1_RNO_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[6]\, D => \readData5[6]\, Y => 
        \readData_21_1_1[6]\);
    
    \readData_31_am_1_1_RNO_0[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[23]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[21]\, D => \readData8[23]\, Y => 
        N_167);
    
    \readData_31_am[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_497, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[31]_net_1\, D => N_401, Y => 
        \readData_31_am[31]_net_1\);
    
    \readData_31_bm_1_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_725, D => N_629, Y => \readData_31_bm_1_1[3]_net_1\);
    
    \readData_31_am[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_492, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[26]_net_1\, D => N_396, Y => 
        \readData_31_am[26]_net_1\);
    
    \readData_31_bm_RNO_2[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[16]\, D => \readData3[16]\, Y => 
        \readData_25_1_1[15]\);
    
    \readData_31_bm_1_1_RNO_0[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[5]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[5]\, D => \readData9[5]\, Y => N_631);
    
    \readData_31_bm_1_1_RNO_0[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[22]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[20]\, D => \readData9[22]\, Y => 
        N_646);
    
    \readData_31_bm_1_1_RNO_2[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[15]\, D => \readData1[15]\, Y => 
        \readData_18_1_1[14]\);
    
    \readData_31_bm[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_956, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[10]_net_1\, D => N_860, Y => 
        \readData_31_bm[10]_net_1\);
    
    \readData_31_am[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_495, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[29]_net_1\, D => N_399, Y => 
        \readData_31_am[29]_net_1\);
    
    block29_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem_m3(2), Y => \wen_b29_1[0]\);
    
    \readData_31_bm_RNO_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[1]\, D => \readData7[1]\, Y => 
        \readData_28_1_1[1]\);
    
    \readData_31_bm_1_1_RNO[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[22]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[20]\, D => \readData13[22]\, Y => 
        N_742);
    
    block14_RNO_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem_m3(3), Y => \wen_b14_1[1]\);
    
    \readData_31_ns[24]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[24]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[24]_net_1\, Y => 
        ram_rdata(24));
    
    \readData_31_bm_1_1_RNO_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[15]\, D => \readData5[15]\, Y => 
        \readData_21_1_1[14]\);
    
    block15 : RAM1K18
      port map(A_DOUT(17) => nc49, A_DOUT(16) => \readData15[16]\, 
        A_DOUT(15) => \readData15[15]\, A_DOUT(14) => 
        \readData15[14]\, A_DOUT(13) => \readData15[13]\, 
        A_DOUT(12) => \readData15[12]\, A_DOUT(11) => 
        \readData15[11]\, A_DOUT(10) => \readData15[10]\, 
        A_DOUT(9) => \readData15[9]\, A_DOUT(8) => nc28, 
        A_DOUT(7) => \readData15[7]\, A_DOUT(6) => 
        \readData15[6]\, A_DOUT(5) => \readData15[5]\, A_DOUT(4)
         => \readData15[4]\, A_DOUT(3) => \readData15[3]\, 
        A_DOUT(2) => \readData15[2]\, A_DOUT(1) => 
        \readData15[1]\, A_DOUT(0) => \readData15[0]\, B_DOUT(17)
         => nc18, B_DOUT(16) => \readData15[34]\, B_DOUT(15) => 
        \readData15[33]\, B_DOUT(14) => \readData15[32]\, 
        B_DOUT(13) => \readData15[31]\, B_DOUT(12) => 
        \readData15[30]\, B_DOUT(11) => \readData15[29]\, 
        B_DOUT(10) => \readData15[28]\, B_DOUT(9) => 
        \readData15[27]\, B_DOUT(8) => nc128, B_DOUT(7) => 
        \readData15[25]\, B_DOUT(6) => \readData15[24]\, 
        B_DOUT(5) => \readData15[23]\, B_DOUT(4) => 
        \readData15[22]\, B_DOUT(3) => \readData15[21]\, 
        B_DOUT(2) => \readData15[20]\, B_DOUT(1) => 
        \readData15[19]\, B_DOUT(0) => \readData15[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a15_1[1]\, A_WEN(0) => \wen_a15_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b15_1[1]\, 
        B_WEN(0) => \wen_b15_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[16]\, D => \readData7[16]\, Y => 
        \readData_28_1_1[15]\);
    
    \readData_31_bm_1_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_742, D => N_646, Y => 
        \readData_31_bm_1_1[20]_net_1\);
    
    \readData_31_am_1_1_RNO[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[23]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[21]\, D => \readData12[23]\, Y => 
        N_263);
    
    \readData_31_am_1_1_RNO_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[2]\, D => \readData4[2]\, Y => 
        \readData_6_1_1[2]\);
    
    \readData_31_bm_1_1_RNO[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[31]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[28]\, D => \readData13[31]\, Y => 
        N_750);
    
    readdata_xhdl1388_0_a2_1 : CFG3
      generic map(INIT => x"80")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1148);
    
    \readData_31_bm_1_1_RNO_0[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[23]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[21]\, D => \readData9[23]\, Y => 
        N_647);
    
    \readData_31_am_RNO_0[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[11]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[10]\, D => \readData10[11]\, Y => 
        N_380);
    
    \readData_31_bm_1_1[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_723, D => N_627, Y => \readData_31_bm_1_1[1]_net_1\);
    
    \readData_31_am_1_1_RNO_0[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[15]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[14]\, D => \readData8[15]\, Y => 
        N_160);
    
    \readData_31_am_1_1_RNO_2[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[11]\, D => \readData0[11]\, Y => 
        \readData_3_1_1[10]\);
    
    \readData_31_bm_1_1_RNO_0[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[30]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[27]\, D => \readData9[30]\, Y => 
        N_653);
    
    \readData_31_am_1_1_RNO_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[11]\, D => \readData4[11]\, Y => 
        \readData_6_1_1[10]\);
    
    block20_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem_m3(3), Y => \wen_b20_1[1]\);
    
    \readData_31_am_1_1_RNO_0[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[16]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[15]\, D => \readData8[16]\, Y => 
        N_161);
    
    block3_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem_m3(3), Y => \wen_b3_1[1]\);
    
    \readData_31_am_1_1_RNO_2[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[23]\, D => \readData0[23]\, Y => 
        \readData_3_1_1[21]\);
    
    \readData_31_bm_RNO_2[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[10]\, D => \readData3[10]\, Y => 
        \readData_25_1_1[9]\);
    
    \readData_31_am[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_491, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[25]_net_1\, D => N_395, Y => 
        \readData_31_am[25]_net_1\);
    
    readdata_xhdl1402_0 : CFG3
      generic map(INIT => x"01")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => readdata_xhdl1403_0);
    
    \readData_31_bm_1_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_752, D => N_656, Y => 
        \readData_31_bm_1_1[30]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[22]\, D => \readData1[22]\, Y => 
        \readData_18_1_1[20]\);
    
    block3_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(1), Y => \wen_a3_1[1]\);
    
    block25_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem_m3(3), Y => \wen_b25_1[1]\);
    
    block26_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem_m3(2), Y => \wen_b26_1[0]\);
    
    \readData_31_bm_1_1_RNO[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[13]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[12]\, D => \readData13[13]\, Y => 
        N_734);
    
    \readData_31_am_1_1_RNO_0[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[2]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[2]\, D => \readData8[2]\, Y => N_148);
    
    \readData_31_am_RNO[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[7]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[7]\, D => \readData14[7]\, Y => N_473);
    
    \readData_31_am_RNO_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[4]\, D => \readData6[4]\, Y => 
        \readData_13_1_1[4]\);
    
    \readData_31_am_RNO_2[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[22]\, D => \readData2[22]\, Y => 
        \readData_10_1_1[20]\);
    
    \readData_31_ns[17]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[17]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[17]_net_1\, Y => 
        ram_rdata(17));
    
    readdata_xhdl1407_0_a2_1 : CFG3
      generic map(INIT => x"40")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1149);
    
    \readData_31_am_RNO[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[11]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[10]\, D => \readData14[11]\, Y => 
        N_476);
    
    \readData_31_am_RNO_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[6]\, D => \readData6[6]\, Y => 
        \readData_13_1_1[6]\);
    
    \readData_31_bm_1_1_RNO_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[28]\, D => \readData5[28]\, Y => 
        \readData_21_1_1[25]\);
    
    \readData_31_bm_1_1_RNO_2[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[23]\, D => \readData1[23]\, Y => 
        \readData_18_1_1[21]\);
    
    \readData_31_am[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_494, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[28]_net_1\, D => N_398, Y => 
        \readData_31_am[28]_net_1\);
    
    \readData_31_bm_RNO_2[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[3]\, D => \readData3[3]\, Y => 
        \readData_25_1_1[3]\);
    
    \readData_31_bm_1_1_RNO_2[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[30]\, D => \readData1[30]\, Y => 
        \readData_18_1_1[27]\);
    
    \readData_31_am_RNO_0[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[14]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[13]\, D => \readData10[14]\, Y => 
        N_383);
    
    \readData_31_am_RNO_0[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[7]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[7]\, D => \readData10[7]\, Y => N_377);
    
    \readData_31_am_1_1_RNO_0[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[7]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[7]\, D => \readData8[7]\, Y => N_153);
    
    \readData_31_bm_1_1_RNO_2[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[2]\, D => \readData1[2]\, Y => 
        \readData_18_1_1[2]\);
    
    \readData_31_am[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_486, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[20]_net_1\, D => N_390, Y => 
        \readData_31_am[20]_net_1\);
    
    \readData_31_am_RNO[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[25]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[23]\, D => \readData14[25]\, Y => 
        N_489);
    
    block17_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(0), Y => 
        \wen_a17_1[0]\);
    
    \readData_31_am_1_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_263, D => N_167, Y => 
        \readData_31_am_1_1[21]_net_1\);
    
    \readData_31_bm_1_1_RNO[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[24]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[22]\, D => \readData13[24]\, Y => 
        N_744);
    
    \readData_31_am_RNO_1[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[28]\, D => \readData6[28]\, Y => 
        \readData_13_1_1[25]\);
    
    \readData_31_bm_RNO_0[28]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[31]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[28]\, D => \readData11[31]\, Y => 
        N_878);
    
    block22_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem_m3(2), Y => \wen_b22_1[0]\);
    
    \readData_31_bm_RNO_2[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[7]\, D => \readData3[7]\, Y => 
        \readData_25_1_1[7]\);
    
    \readData_31_bm_1_1_RNO_2[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[6]\, D => \readData1[6]\, Y => 
        \readData_18_1_1[6]\);
    
    \readData_31_bm[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_967, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[21]_net_1\, D => N_871, Y => 
        \readData_31_bm[21]_net_1\);
    
    \readData_31_am_RNO_2[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[25]\, D => \readData2[25]\, Y => 
        \readData_10_1_1[23]\);
    
    \readData_31_am_1_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_252, D => N_156, Y => 
        \readData_31_am_1_1[10]_net_1\);
    
    \readData_31_bm_RNO_0[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[15]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[14]\, D => \readData11[15]\, Y => 
        N_864);
    
    block4_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(0), Y => \wen_a4_1[0]\);
    
    block30_RNO_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem_m3(2), Y => \wen_b30_1[0]\);
    
    \readData_31_am_1_1_RNO[12]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[13]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[12]\, D => \readData12[13]\, Y => 
        N_254);
    
    \readData_31_bm_1_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_735, D => N_639, Y => 
        \readData_31_bm_1_1[13]_net_1\);
    
    \readData_31_bm_RNO_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[30]\, D => \readData7[30]\, Y => 
        \readData_28_1_1[27]\);
    
    \readData_31_bm_1_1_RNO_2[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[7]\, D => \readData1[7]\, Y => 
        \readData_18_1_1[7]\);
    
    block15_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem_m3(2), Y => \wen_b15_1[0]\);
    
    \readData_31_bm_RNO_2[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[20]\, D => \readData3[20]\, Y => 
        \readData_25_1_1[18]\);
    
    \readData_31_am_1_1[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_273, D => N_177, Y => 
        \readData_31_am_1_1[31]_net_1\);
    
    \readData_31_am_1_1_RNO_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[23]\, D => \readData4[23]\, Y => 
        \readData_6_1_1[21]\);
    
    block23_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem_m3(2), Y => \wen_b23_1[0]\);
    
    \readData_31_bm_1_1_RNO[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[5]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[5]\, D => \readData13[5]\, Y => N_727);
    
    \readData_31_bm_1_1_RNO_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[22]\, D => \readData5[22]\, Y => 
        \readData_21_1_1[20]\);
    
    block9_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(0), Y => \wen_a9_1[0]\);
    
    \readData_31_bm_RNO_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[20]\, D => \readData7[20]\, Y => 
        \readData_28_1_1[18]\);
    
    \readData_31_am_RNO_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[3]\, D => \readData6[3]\, Y => 
        \readData_13_1_1[3]\);
    
    \readData_31_am_1_1_RNO_2[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[15]\, D => \readData0[15]\, Y => 
        \readData_3_1_1[14]\);
    
    \readData_31_am_1_1_RNO_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[5]\, D => \readData4[5]\, Y => 
        \readData_6_1_1[5]\);
    
    \readData_31_am_1_1[17]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_259, D => N_163, Y => 
        \readData_31_am_1_1[17]_net_1\);
    
    \readData_31_am_RNO[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[27]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[24]\, D => \readData14[27]\, Y => 
        N_490);
    
    \readData_31_am_1_1_RNO_2[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[0]\, D => \readData0[0]\, Y => 
        \readData_3_1_1[0]\);
    
    block19_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem_m3(3), Y => \wen_b19_1[1]\);
    
    \readData_31_am_1_1_RNO_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[15]\, D => \readData4[15]\, Y => 
        \readData_6_1_1[14]\);
    
    block6 : RAM1K18
      port map(A_DOUT(17) => nc107, A_DOUT(16) => \readData6[16]\, 
        A_DOUT(15) => \readData6[15]\, A_DOUT(14) => 
        \readData6[14]\, A_DOUT(13) => \readData6[13]\, 
        A_DOUT(12) => \readData6[12]\, A_DOUT(11) => 
        \readData6[11]\, A_DOUT(10) => \readData6[10]\, A_DOUT(9)
         => \readData6[9]\, A_DOUT(8) => nc118, A_DOUT(7) => 
        \readData6[7]\, A_DOUT(6) => \readData6[6]\, A_DOUT(5)
         => \readData6[5]\, A_DOUT(4) => \readData6[4]\, 
        A_DOUT(3) => \readData6[3]\, A_DOUT(2) => \readData6[2]\, 
        A_DOUT(1) => \readData6[1]\, A_DOUT(0) => \readData6[0]\, 
        B_DOUT(17) => nc106, B_DOUT(16) => \readData6[34]\, 
        B_DOUT(15) => \readData6[33]\, B_DOUT(14) => 
        \readData6[32]\, B_DOUT(13) => \readData6[31]\, 
        B_DOUT(12) => \readData6[30]\, B_DOUT(11) => 
        \readData6[29]\, B_DOUT(10) => \readData6[28]\, B_DOUT(9)
         => \readData6[27]\, B_DOUT(8) => nc75, B_DOUT(7) => 
        \readData6[25]\, B_DOUT(6) => \readData6[24]\, B_DOUT(5)
         => \readData6[23]\, B_DOUT(4) => \readData6[22]\, 
        B_DOUT(3) => \readData6[21]\, B_DOUT(2) => 
        \readData6[20]\, B_DOUT(1) => \readData6[19]\, B_DOUT(0)
         => \readData6[18]\, BUSY => OPEN, A_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => N_375_i_0, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        N_72_i_0, A_DIN(15) => N_70_i_0, A_DIN(14) => N_68_i_0, 
        A_DIN(13) => N_66_i_0, A_DIN(12) => N_64_i_0, A_DIN(11)
         => N_58_i_0, A_DIN(10) => N_56_i_0, A_DIN(9) => N_54_i_0, 
        A_DIN(8) => GND_net_1, A_DIN(7) => N_52_i_0, A_DIN(6) => 
        N_50_i_0, A_DIN(5) => N_48_i_0, A_DIN(4) => N_46_i_0, 
        A_DIN(3) => N_44_i_0, A_DIN(2) => N_42_i_0, A_DIN(1) => 
        N_40_i_0, A_DIN(0) => N_38_i_0, A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a6_1[1]\, 
        A_WEN(0) => \wen_a6_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b6_1[1]\, 
        B_WEN(0) => \wen_b6_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_2[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[27]\, D => \readData3[27]\, Y => 
        \readData_25_1_1[24]\);
    
    \readData_31_am_1_1_RNO_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[7]\, D => \readData4[7]\, Y => 
        \readData_6_1_1[7]\);
    
    \readData_31_am_1_1_RNO_2[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[16]\, D => \readData0[16]\, Y => 
        \readData_3_1_1[15]\);
    
    \readData_31_am_RNO_2[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[0]\, D => \readData2[0]\, Y => 
        \readData_10_1_1[0]\);
    
    \readData_31_bm_RNO_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[24]\, D => \readData7[24]\, Y => 
        \readData_28_1_1[22]\);
    
    \readData_31_am_1_1_RNO_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[16]\, D => \readData4[16]\, Y => 
        \readData_6_1_1[15]\);
    
    \readData_31_bm_1_1_RNO_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[23]\, D => \readData5[23]\, Y => 
        \readData_21_1_1[21]\);
    
    readdata_xhdl1399_0_a2_0 : CFG3
      generic map(INIT => x"10")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1150);
    
    \readData_31_bm_1_1_RNO_0[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[29]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[26]\, D => \readData9[29]\, Y => 
        N_652);
    
    \readData_31_am_RNO_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[0]\, D => \readData6[0]\, Y => 
        \readData_13_1_1[0]\);
    
    \readData_31_am_1_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_265, D => N_169, Y => 
        \readData_31_am_1_1[23]_net_1\);
    
    \readData_31_bm_1_1_RNO[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[2]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[2]\, D => \readData13[2]\, Y => N_724);
    
    \readData_31_bm_1_1_RNO_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[30]\, D => \readData5[30]\, Y => 
        \readData_21_1_1[27]\);
    
    \readData_31_am_RNO[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[30]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[27]\, D => \readData14[30]\, Y => 
        N_493);
    
    \readData_31_bm_1_1_RNO_0[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[0]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[0]\, D => \readData9[0]\, Y => N_626);
    
    \readData_31_am_1_1_RNO[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[24]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[22]\, D => \readData12[24]\, Y => 
        N_264);
    
    \readData_31_am[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_468, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[2]_net_1\, D => N_372, Y => 
        \readData_31_am[2]_net_1\);
    
    \readData_31_bm_RNO[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[16]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[15]\, D => \readData15[16]\, Y => 
        N_961);
    
    \readData_31_am_RNO_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[24]\, D => \readData6[24]\, Y => 
        \readData_13_1_1[22]\);
    
    \readData_31_bm_RNO_0[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[33]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[30]\, D => \readData11[33]\, Y => 
        N_880);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    block3_RNO : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(0), Y => \wen_a3_1[0]\);
    
    \readData_31_am_RNO[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[29]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[26]\, D => \readData14[29]\, Y => 
        N_492);
    
    \readData_31_am_RNO[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[6]\, B => ahbsram_addr(14), C => 
        \readData_13_1_1[6]\, D => \readData14[6]\, Y => N_472);
    
    \readData_31_am_RNO[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[34]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[31]\, D => \readData14[34]\, Y => 
        N_497);
    
    \readData_31_ns[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[4]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[4]_net_1\, Y => 
        ram_rdata(4));
    
    \wen_a_m_10_0_a2_0[1]\ : CFG3
      generic map(INIT => x"04")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1143);
    
    \readData_31_am_1_1_RNO_0[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[24]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[22]\, D => \readData8[24]\, Y => 
        N_168);
    
    block2_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(1), Y => \wen_a2_1[1]\);
    
    \readData_31_bm_RNO_0[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[9]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[8]\, D => \readData11[9]\, Y => N_858);
    
    block1_RNO_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem(1), Y => 
        \wen_a1_1[1]\);
    
    \readData_31_bm_1_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_749, D => N_653, Y => 
        \readData_31_bm_1_1[27]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[24]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[22]\, D => \readData9[24]\, Y => 
        N_648);
    
    \readData_31_am_1_1_RNO_0[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[20]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[18]\, D => \readData8[20]\, Y => 
        N_164);
    
    \readData_31_am[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_474, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[8]_net_1\, D => N_378, Y => 
        \readData_31_am[8]_net_1\);
    
    \readData_31_bm_1_1_RNO[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[4]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[4]\, D => \readData13[4]\, Y => N_726);
    
    block10_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem_m3(2), Y => \wen_b10_1[0]\);
    
    \readData_31_bm_1_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_738, D => N_642, Y => 
        \readData_31_bm_1_1[16]_net_1\);
    
    \readData_31_bm_1_1_RNO[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[15]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[14]\, D => \readData13[15]\, Y => 
        N_736);
    
    \readData_31_am_1_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_250, D => N_154, Y => \readData_31_am_1_1[8]_net_1\);
    
    \readData_31_ns[13]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[13]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[13]_net_1\, Y => 
        ram_rdata(13));
    
    \readData_31_am_RNO[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[16]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[15]\, D => \readData14[16]\, Y => 
        N_481);
    
    \readData_31_bm_1_1_RNO_2[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[29]\, D => \readData1[29]\, Y => 
        \readData_18_1_1[26]\);
    
    \readData_31_bm_RNO_2[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[34]\, D => \readData3[34]\, Y => 
        \readData_25_1_1[31]\);
    
    block4_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem_m3(2), Y => \wen_b4_1[0]\);
    
    \readData_31_am_RNO_0[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[29]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[26]\, D => \readData10[29]\, Y => 
        N_396);
    
    \readData_31_bm_RNO[21]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[23]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[21]\, D => \readData15[23]\, Y => 
        N_967);
    
    \readData_31_bm_1_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_746, D => N_650, Y => 
        \readData_31_bm_1_1[24]_net_1\);
    
    \readData_31_bm_1_1_RNO[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[6]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[6]\, D => \readData13[6]\, Y => N_728);
    
    block11 : RAM1K18
      port map(A_DOUT(17) => nc65, A_DOUT(16) => \readData11[16]\, 
        A_DOUT(15) => \readData11[15]\, A_DOUT(14) => 
        \readData11[14]\, A_DOUT(13) => \readData11[13]\, 
        A_DOUT(12) => \readData11[12]\, A_DOUT(11) => 
        \readData11[11]\, A_DOUT(10) => \readData11[10]\, 
        A_DOUT(9) => \readData11[9]\, A_DOUT(8) => nc38, 
        A_DOUT(7) => \readData11[7]\, A_DOUT(6) => 
        \readData11[6]\, A_DOUT(5) => \readData11[5]\, A_DOUT(4)
         => \readData11[4]\, A_DOUT(3) => \readData11[3]\, 
        A_DOUT(2) => \readData11[2]\, A_DOUT(1) => 
        \readData11[1]\, A_DOUT(0) => \readData11[0]\, B_DOUT(17)
         => nc93, B_DOUT(16) => \readData11[34]\, B_DOUT(15) => 
        \readData11[33]\, B_DOUT(14) => \readData11[32]\, 
        B_DOUT(13) => \readData11[31]\, B_DOUT(12) => 
        \readData11[30]\, B_DOUT(11) => \readData11[29]\, 
        B_DOUT(10) => \readData11[28]\, B_DOUT(9) => 
        \readData11[27]\, B_DOUT(8) => nc1, B_DOUT(7) => 
        \readData11[25]\, B_DOUT(6) => \readData11[24]\, 
        B_DOUT(5) => \readData11[23]\, B_DOUT(4) => 
        \readData11[22]\, B_DOUT(3) => \readData11[21]\, 
        B_DOUT(2) => \readData11[20]\, B_DOUT(1) => 
        \readData11[19]\, B_DOUT(0) => \readData11[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a11_1[1]\, A_WEN(0) => \wen_a11_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b11_1[1]\, 
        B_WEN(0) => \wen_b11_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_RNO_2[31]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[34]\, D => \readData2[34]\, Y => 
        \readData_10_1_1[31]\);
    
    \readData_31_am_1_1_RNO[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[16]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[15]\, D => \readData12[16]\, Y => 
        N_257);
    
    \readData_31_am_RNO_2[1]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[1]\, D => \readData2[1]\, Y => 
        \readData_10_1_1[1]\);
    
    \readData_31_bm_RNO_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[33]\, D => \readData7[33]\, Y => 
        \readData_28_1_1[30]\);
    
    \readData_31_am_1_1_RNO_2[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[24]\, D => \readData0[24]\, Y => 
        \readData_3_1_1[22]\);
    
    block7_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem_m3(3), Y => \wen_b7_1[1]\);
    
    \readData_31_bm_1_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_729, D => N_633, Y => \readData_31_bm_1_1[7]_net_1\);
    
    block27_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(0), Y => \wen_a27_1[0]\);
    
    \readData_31_bm_1_1_RNO_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[2]\, D => \readData5[2]\, Y => 
        \readData_21_1_1[2]\);
    
    block12 : RAM1K18
      port map(A_DOUT(17) => nc2, A_DOUT(16) => \readData12[16]\, 
        A_DOUT(15) => \readData12[15]\, A_DOUT(14) => 
        \readData12[14]\, A_DOUT(13) => \readData12[13]\, 
        A_DOUT(12) => \readData12[12]\, A_DOUT(11) => 
        \readData12[11]\, A_DOUT(10) => \readData12[10]\, 
        A_DOUT(9) => \readData12[9]\, A_DOUT(8) => nc50, 
        A_DOUT(7) => \readData12[7]\, A_DOUT(6) => 
        \readData12[6]\, A_DOUT(5) => \readData12[5]\, A_DOUT(4)
         => \readData12[4]\, A_DOUT(3) => \readData12[3]\, 
        A_DOUT(2) => \readData12[2]\, A_DOUT(1) => 
        \readData12[1]\, A_DOUT(0) => \readData12[0]\, B_DOUT(17)
         => nc22, B_DOUT(16) => \readData12[34]\, B_DOUT(15) => 
        \readData12[33]\, B_DOUT(14) => \readData12[32]\, 
        B_DOUT(13) => \readData12[31]\, B_DOUT(12) => 
        \readData12[30]\, B_DOUT(11) => \readData12[29]\, 
        B_DOUT(10) => \readData12[28]\, B_DOUT(9) => 
        \readData12[27]\, B_DOUT(8) => nc12, B_DOUT(7) => 
        \readData12[25]\, B_DOUT(6) => \readData12[24]\, 
        B_DOUT(5) => \readData12[23]\, B_DOUT(4) => 
        \readData12[22]\, B_DOUT(3) => \readData12[21]\, 
        B_DOUT(2) => \readData12[20]\, B_DOUT(1) => 
        \readData12[19]\, B_DOUT(0) => \readData12[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a12_1[1]\, A_WEN(0) => \wen_a12_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b12_1[1]\, 
        B_WEN(0) => \wen_b12_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[2]\, D => \readData7[2]\, Y => 
        \readData_28_1_1[2]\);
    
    block26_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1147, D => sram_wen_mem(1), Y => \wen_a26_1[1]\);
    
    block12_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(1), Y => \wen_a12_1[1]\);
    
    \readData_31_bm_1_1_RNO_2[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[24]\, D => \readData1[24]\, Y => 
        \readData_18_1_1[22]\);
    
    \readData_31_bm_1_1_RNO[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[34]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[31]\, D => \readData13[34]\, Y => 
        N_753);
    
    \readData_31_bm_RNO_0[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[16]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[15]\, D => \readData11[16]\, Y => 
        N_865);
    
    \readData_31_bm_RNO[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[29]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[26]\, D => \readData15[29]\, Y => 
        N_972);
    
    block13 : RAM1K18
      port map(A_DOUT(17) => nc21, A_DOUT(16) => \readData13[16]\, 
        A_DOUT(15) => \readData13[15]\, A_DOUT(14) => 
        \readData13[14]\, A_DOUT(13) => \readData13[13]\, 
        A_DOUT(12) => \readData13[12]\, A_DOUT(11) => 
        \readData13[11]\, A_DOUT(10) => \readData13[10]\, 
        A_DOUT(9) => \readData13[9]\, A_DOUT(8) => nc11, 
        A_DOUT(7) => \readData13[7]\, A_DOUT(6) => 
        \readData13[6]\, A_DOUT(5) => \readData13[5]\, A_DOUT(4)
         => \readData13[4]\, A_DOUT(3) => \readData13[3]\, 
        A_DOUT(2) => \readData13[2]\, A_DOUT(1) => 
        \readData13[1]\, A_DOUT(0) => \readData13[0]\, B_DOUT(17)
         => nc78, B_DOUT(16) => \readData13[34]\, B_DOUT(15) => 
        \readData13[33]\, B_DOUT(14) => \readData13[32]\, 
        B_DOUT(13) => \readData13[31]\, B_DOUT(12) => 
        \readData13[30]\, B_DOUT(11) => \readData13[29]\, 
        B_DOUT(10) => \readData13[28]\, B_DOUT(9) => 
        \readData13[27]\, B_DOUT(8) => nc54, B_DOUT(7) => 
        \readData13[25]\, B_DOUT(6) => \readData13[24]\, 
        B_DOUT(5) => \readData13[23]\, B_DOUT(4) => 
        \readData13[22]\, B_DOUT(3) => \readData13[21]\, 
        B_DOUT(2) => \readData13[20]\, B_DOUT(1) => 
        \readData13[19]\, B_DOUT(0) => \readData13[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a13_1[1]\, A_WEN(0) => \wen_a13_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b13_1[1]\, 
        B_WEN(0) => \wen_b13_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_RNO_0[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[32]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[29]\, D => \readData10[32]\, Y => 
        N_399);
    
    \readData_31_am_1_1_RNO_0[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[29]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[26]\, D => \readData8[29]\, Y => 
        N_172);
    
    \readData_31_bm_1_1_RNO[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[27]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[24]\, D => \readData13[27]\, Y => 
        N_746);
    
    \readData_31_bm_RNO[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[22]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[20]\, D => \readData15[22]\, Y => 
        N_966);
    
    \readData_31_am_RNO_2[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[18]\, D => \readData2[18]\, Y => 
        \readData_10_1_1[16]\);
    
    \readData_31_bm_1_1_RNO[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[1]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[1]\, D => \readData13[1]\, Y => N_723);
    
    \readData_31_am_RNO_0[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[27]\, B => ahbsram_addr(14), C
         => \readData_10_1_1[24]\, D => \readData10[27]\, Y => 
        N_394);
    
    \readData_31_am_RNO_0[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[2]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[2]\, D => \readData10[2]\, Y => N_372);
    
    \readData_31_am_RNO_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[18]\, D => \readData6[18]\, Y => 
        \readData_13_1_1[16]\);
    
    block0_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem(0), Y => 
        \wen_a0_1[0]\);
    
    \readData_31_bm_1_1[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_722, D => N_626, Y => \readData_31_bm_1_1[0]_net_1\);
    
    \readData_31_am_1_1[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_244, D => N_148, Y => \readData_31_am_1_1[2]_net_1\);
    
    block24_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(1), Y => \wen_a24_1[1]\);
    
    block18 : RAM1K18
      port map(A_DOUT(17) => nc68, A_DOUT(16) => \readData18[16]\, 
        A_DOUT(15) => \readData18[15]\, A_DOUT(14) => 
        \readData18[14]\, A_DOUT(13) => \readData18[13]\, 
        A_DOUT(12) => \readData18[12]\, A_DOUT(11) => 
        \readData18[11]\, A_DOUT(10) => \readData18[10]\, 
        A_DOUT(9) => \readData18[9]\, A_DOUT(8) => nc3, A_DOUT(7)
         => \readData18[7]\, A_DOUT(6) => \readData18[6]\, 
        A_DOUT(5) => \readData18[5]\, A_DOUT(4) => 
        \readData18[4]\, A_DOUT(3) => \readData18[3]\, A_DOUT(2)
         => \readData18[2]\, A_DOUT(1) => \readData18[1]\, 
        A_DOUT(0) => \readData18[0]\, B_DOUT(17) => nc32, 
        B_DOUT(16) => \readData18[34]\, B_DOUT(15) => 
        \readData18[33]\, B_DOUT(14) => \readData18[32]\, 
        B_DOUT(13) => \readData18[31]\, B_DOUT(12) => 
        \readData18[30]\, B_DOUT(11) => \readData18[29]\, 
        B_DOUT(10) => \readData18[28]\, B_DOUT(9) => 
        \readData18[27]\, B_DOUT(8) => nc104, B_DOUT(7) => 
        \readData18[25]\, B_DOUT(6) => \readData18[24]\, 
        B_DOUT(5) => \readData18[23]\, B_DOUT(4) => 
        \readData18[22]\, B_DOUT(3) => \readData18[21]\, 
        B_DOUT(2) => \readData18[20]\, B_DOUT(1) => 
        \readData18[19]\, B_DOUT(0) => \readData18[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a18_1[1]\, A_WEN(0) => \wen_a18_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b18_1[1]\, 
        B_WEN(0) => \wen_b18_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_1_1_RNO[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[28]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[25]\, D => \readData12[28]\, Y => 
        N_267);
    
    \readData_31_bm_1_1_RNO_0[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[2]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[2]\, D => \readData9[2]\, Y => N_628);
    
    \readData_31_am[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_466, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[0]_net_1\, D => N_370, Y => 
        \readData_31_am[0]_net_1\);
    
    \readData_31_am_1_1_RNO_0[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[14]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[13]\, D => \readData8[14]\, Y => 
        N_159);
    
    \readData_31_bm_1_1[15]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_737, D => N_641, Y => 
        \readData_31_bm_1_1[15]_net_1\);
    
    block20_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(1), Y => \wen_a20_1[1]\);
    
    \readData_31_am_RNO_2[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[21]\, D => \readData2[21]\, Y => 
        \readData_10_1_1[19]\);
    
    block18_RNO_1 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(14), C
         => readdata_xhdl1401_1, D => sram_wen_mem_m3(2), Y => 
        \wen_b18_1[0]\);
    
    \readData_31_bm_RNO_2[25]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[28]\, D => \readData3[28]\, Y => 
        \readData_25_1_1[25]\);
    
    block9_RNO_2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem_m3(3), Y => \wen_b9_1[1]\);
    
    \readData_31_am_1_1_RNO_2[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[33]\, D => \readData0[33]\, Y => 
        \readData_3_1_1[30]\);
    
    \readData_31_ns[10]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[10]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[10]_net_1\, Y => 
        ram_rdata(10));
    
    \readData_31_am_RNO_2[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[15]\, D => \readData2[15]\, Y => 
        \readData_10_1_1[14]\);
    
    \readData_31_am_RNO_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[21]\, D => \readData6[21]\, Y => 
        \readData_13_1_1[19]\);
    
    \readData_31_am_1_1_RNO_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[33]\, D => \readData4[33]\, Y => 
        \readData_6_1_1[30]\);
    
    \readData_31_am[16]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_482, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[16]_net_1\, D => N_386, Y => 
        \readData_31_am[16]_net_1\);
    
    \readData_31_bm_1_1_RNO[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[9]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[8]\, D => \readData13[9]\, Y => N_730);
    
    \readData_31_am[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_485, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[19]_net_1\, D => N_389, Y => 
        \readData_31_am[19]_net_1\);
    
    \readData_31_am_1_1_RNO_2[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[29]\, D => \readData0[29]\, Y => 
        \readData_3_1_1[26]\);
    
    \readData_31_am_RNO_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[15]\, D => \readData6[15]\, Y => 
        \readData_13_1_1[14]\);
    
    \readData_31_bm_1_1_RNO_0[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[7]\, B => ahbsram_addr(14), C => 
        \readData_18_1_1[7]\, D => \readData9[7]\, Y => N_633);
    
    block2 : RAM1K18
      port map(A_DOUT(17) => nc40, A_DOUT(16) => \readData2[16]\, 
        A_DOUT(15) => \readData2[15]\, A_DOUT(14) => 
        \readData2[14]\, A_DOUT(13) => \readData2[13]\, 
        A_DOUT(12) => \readData2[12]\, A_DOUT(11) => 
        \readData2[11]\, A_DOUT(10) => \readData2[10]\, A_DOUT(9)
         => \readData2[9]\, A_DOUT(8) => nc31, A_DOUT(7) => 
        \readData2[7]\, A_DOUT(6) => \readData2[6]\, A_DOUT(5)
         => \readData2[5]\, A_DOUT(4) => \readData2[4]\, 
        A_DOUT(3) => \readData2[3]\, A_DOUT(2) => \readData2[2]\, 
        A_DOUT(1) => \readData2[1]\, A_DOUT(0) => \readData2[0]\, 
        B_DOUT(17) => nc96, B_DOUT(16) => \readData2[34]\, 
        B_DOUT(15) => \readData2[33]\, B_DOUT(14) => 
        \readData2[32]\, B_DOUT(13) => \readData2[31]\, 
        B_DOUT(12) => \readData2[30]\, B_DOUT(11) => 
        \readData2[29]\, B_DOUT(10) => \readData2[28]\, B_DOUT(9)
         => \readData2[27]\, B_DOUT(8) => nc44, B_DOUT(7) => 
        \readData2[25]\, B_DOUT(6) => \readData2[24]\, B_DOUT(5)
         => \readData2[23]\, B_DOUT(4) => \readData2[22]\, 
        B_DOUT(3) => \readData2[21]\, B_DOUT(2) => 
        \readData2[20]\, B_DOUT(1) => \readData2[19]\, B_DOUT(0)
         => \readData2[18]\, BUSY => OPEN, A_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => N_375_i_0, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        N_72_i_0, A_DIN(15) => N_70_i_0, A_DIN(14) => N_68_i_0, 
        A_DIN(13) => N_66_i_0, A_DIN(12) => N_64_i_0, A_DIN(11)
         => N_58_i_0, A_DIN(10) => N_56_i_0, A_DIN(9) => N_54_i_0, 
        A_DIN(8) => GND_net_1, A_DIN(7) => N_52_i_0, A_DIN(6) => 
        N_50_i_0, A_DIN(5) => N_48_i_0, A_DIN(4) => N_46_i_0, 
        A_DIN(3) => N_44_i_0, A_DIN(2) => N_42_i_0, A_DIN(1) => 
        N_40_i_0, A_DIN(0) => N_38_i_0, A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a2_1[1]\, 
        A_WEN(0) => \wen_a2_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b2_1[1]\, 
        B_WEN(0) => \wen_b2_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_am_RNO_1[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[9]\, D => \readData6[9]\, Y => 
        \readData_13_1_1[8]\);
    
    \readData_31_bm_1_1_RNO_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[29]\, D => \readData5[29]\, Y => 
        \readData_21_1_1[26]\);
    
    \readData_31_bm_RNO[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[0]\, B => ahbsram_addr(14), C => 
        \readData_28_1_1[0]\, D => \readData15[0]\, Y => N_946);
    
    block0 : RAM1K18
      port map(A_DOUT(17) => nc7, A_DOUT(16) => \readData0[16]\, 
        A_DOUT(15) => \readData0[15]\, A_DOUT(14) => 
        \readData0[14]\, A_DOUT(13) => \readData0[13]\, 
        A_DOUT(12) => \readData0[12]\, A_DOUT(11) => 
        \readData0[11]\, A_DOUT(10) => \readData0[10]\, A_DOUT(9)
         => \readData0[9]\, A_DOUT(8) => nc97, A_DOUT(7) => 
        \readData0[7]\, A_DOUT(6) => \readData0[6]\, A_DOUT(5)
         => \readData0[5]\, A_DOUT(4) => \readData0[4]\, 
        A_DOUT(3) => \readData0[3]\, A_DOUT(2) => \readData0[2]\, 
        A_DOUT(1) => \readData0[1]\, A_DOUT(0) => \readData0[0]\, 
        B_DOUT(17) => nc85, B_DOUT(16) => \readData0[34]\, 
        B_DOUT(15) => \readData0[33]\, B_DOUT(14) => 
        \readData0[32]\, B_DOUT(13) => \readData0[31]\, 
        B_DOUT(12) => \readData0[30]\, B_DOUT(11) => 
        \readData0[29]\, B_DOUT(10) => \readData0[28]\, B_DOUT(9)
         => \readData0[27]\, B_DOUT(8) => nc72, B_DOUT(7) => 
        \readData0[25]\, B_DOUT(6) => \readData0[24]\, B_DOUT(5)
         => \readData0[23]\, B_DOUT(4) => \readData0[22]\, 
        B_DOUT(3) => \readData0[21]\, B_DOUT(2) => 
        \readData0[20]\, B_DOUT(1) => \readData0[19]\, B_DOUT(0)
         => \readData0[18]\, BUSY => OPEN, A_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => N_375_i_0, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        N_72_i_0, A_DIN(15) => N_70_i_0, A_DIN(14) => N_68_i_0, 
        A_DIN(13) => N_66_i_0, A_DIN(12) => N_64_i_0, A_DIN(11)
         => N_58_i_0, A_DIN(10) => N_56_i_0, A_DIN(9) => N_54_i_0, 
        A_DIN(8) => GND_net_1, A_DIN(7) => N_52_i_0, A_DIN(6) => 
        N_50_i_0, A_DIN(5) => N_48_i_0, A_DIN(4) => N_46_i_0, 
        A_DIN(3) => N_44_i_0, A_DIN(2) => N_42_i_0, A_DIN(1) => 
        N_40_i_0, A_DIN(0) => N_38_i_0, A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a0_1[1]\, 
        A_WEN(0) => \wen_a0_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b0_1[1]\, 
        B_WEN(0) => \wen_b0_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[5]\, D => \readData7[5]\, Y => 
        \readData_28_1_1[5]\);
    
    \readData_31_am[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_473, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[7]_net_1\, D => N_377, Y => 
        \readData_31_am[7]_net_1\);
    
    \readData_31_am_RNO_2[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[9]\, D => \readData2[9]\, Y => 
        \readData_10_1_1[8]\);
    
    \readData_31_am_1_1_RNO_2[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[20]\, D => \readData0[20]\, Y => 
        \readData_3_1_1[18]\);
    
    \readData_31_bm_RNO_0[26]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[29]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[26]\, D => \readData11[29]\, Y => 
        N_876);
    
    \readData_31_am_1_1_RNO_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[20]\, D => \readData4[20]\, Y => 
        \readData_6_1_1[18]\);
    
    \readData_31_ns[14]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[14]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[14]_net_1\, Y => 
        ram_rdata(14));
    
    \readData_31_bm[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_969, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[23]_net_1\, D => N_873, Y => 
        \readData_31_bm[23]_net_1\);
    
    \readData_31_am_1_1_RNO_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[24]\, D => \readData4[24]\, Y => 
        \readData_6_1_1[22]\);
    
    block28_RNO_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(1), Y => \wen_a28_1[1]\);
    
    \readData_31_bm[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_948, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[2]_net_1\, D => N_852, Y => 
        \readData_31_bm[2]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[27]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[24]\, D => \readData9[27]\, Y => 
        N_650);
    
    \readData_31_am_1_1_RNO[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[15]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[14]\, D => \readData12[15]\, Y => 
        N_256);
    
    \readData_31_bm_RNO_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[23]\, D => \readData7[23]\, Y => 
        \readData_28_1_1[21]\);
    
    \readData_31_bm_RNO_0[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[32]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[29]\, D => \readData11[32]\, Y => 
        N_879);
    
    \readData_31_am[15]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_481, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[15]_net_1\, D => N_385, Y => 
        \readData_31_am[15]_net_1\);
    
    block29 : RAM1K18
      port map(A_DOUT(17) => nc6, A_DOUT(16) => \readData29[16]\, 
        A_DOUT(15) => \readData29[15]\, A_DOUT(14) => 
        \readData29[14]\, A_DOUT(13) => \readData29[13]\, 
        A_DOUT(12) => \readData29[12]\, A_DOUT(11) => 
        \readData29[11]\, A_DOUT(10) => \readData29[10]\, 
        A_DOUT(9) => \readData29[9]\, A_DOUT(8) => nc71, 
        A_DOUT(7) => \readData29[7]\, A_DOUT(6) => 
        \readData29[6]\, A_DOUT(5) => \readData29[5]\, A_DOUT(4)
         => \readData29[4]\, A_DOUT(3) => \readData29[3]\, 
        A_DOUT(2) => \readData29[2]\, A_DOUT(1) => 
        \readData29[1]\, A_DOUT(0) => \readData29[0]\, B_DOUT(17)
         => nc62, B_DOUT(16) => \readData29[34]\, B_DOUT(15) => 
        \readData29[33]\, B_DOUT(14) => \readData29[32]\, 
        B_DOUT(13) => \readData29[31]\, B_DOUT(12) => 
        \readData29[30]\, B_DOUT(11) => \readData29[29]\, 
        B_DOUT(10) => \readData29[28]\, B_DOUT(9) => 
        \readData29[27]\, B_DOUT(8) => nc61, B_DOUT(7) => 
        \readData29[25]\, B_DOUT(6) => \readData29[24]\, 
        B_DOUT(5) => \readData29[23]\, B_DOUT(4) => 
        \readData29[22]\, B_DOUT(3) => \readData29[21]\, 
        B_DOUT(2) => \readData29[20]\, B_DOUT(1) => 
        \readData29[19]\, B_DOUT(0) => \readData29[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a29_1[1]\, A_WEN(0) => \wen_a29_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b29_1[1]\, 
        B_WEN(0) => \wen_b29_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_1_1_RNO_1[22]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[24]\, D => \readData5[24]\, Y => 
        \readData_21_1_1[22]\);
    
    \readData_31_am_RNO_1[21]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[23]\, D => \readData6[23]\, Y => 
        \readData_13_1_1[21]\);
    
    block19_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(0), Y => \wen_a19_1[0]\);
    
    \readData_31_ns[26]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[26]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[26]_net_1\, Y => 
        ram_rdata(26));
    
    \readData_31_bm_RNO_2[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[18]\, D => \readData3[18]\, Y => 
        \readData_25_1_1[16]\);
    
    block7 : RAM1K18
      port map(A_DOUT(17) => nc125, A_DOUT(16) => \readData7[16]\, 
        A_DOUT(15) => \readData7[15]\, A_DOUT(14) => 
        \readData7[14]\, A_DOUT(13) => \readData7[13]\, 
        A_DOUT(12) => \readData7[12]\, A_DOUT(11) => 
        \readData7[11]\, A_DOUT(10) => \readData7[10]\, A_DOUT(9)
         => \readData7[9]\, A_DOUT(8) => nc115, A_DOUT(7) => 
        \readData7[7]\, A_DOUT(6) => \readData7[6]\, A_DOUT(5)
         => \readData7[5]\, A_DOUT(4) => \readData7[4]\, 
        A_DOUT(3) => \readData7[3]\, A_DOUT(2) => \readData7[2]\, 
        A_DOUT(1) => \readData7[1]\, A_DOUT(0) => \readData7[0]\, 
        B_DOUT(17) => nc102, B_DOUT(16) => \readData7[34]\, 
        B_DOUT(15) => \readData7[33]\, B_DOUT(14) => 
        \readData7[32]\, B_DOUT(13) => \readData7[31]\, 
        B_DOUT(12) => \readData7[30]\, B_DOUT(11) => 
        \readData7[29]\, B_DOUT(10) => \readData7[28]\, B_DOUT(9)
         => \readData7[27]\, B_DOUT(8) => nc19, B_DOUT(7) => 
        \readData7[25]\, B_DOUT(6) => \readData7[24]\, B_DOUT(5)
         => \readData7[23]\, B_DOUT(4) => \readData7[22]\, 
        B_DOUT(3) => \readData7[21]\, B_DOUT(2) => 
        \readData7[20]\, B_DOUT(1) => \readData7[19]\, B_DOUT(0)
         => \readData7[18]\, BUSY => OPEN, A_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => N_375_i_0, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        N_72_i_0, A_DIN(15) => N_70_i_0, A_DIN(14) => N_68_i_0, 
        A_DIN(13) => N_66_i_0, A_DIN(12) => N_64_i_0, A_DIN(11)
         => N_58_i_0, A_DIN(10) => N_56_i_0, A_DIN(9) => N_54_i_0, 
        A_DIN(8) => GND_net_1, A_DIN(7) => N_52_i_0, A_DIN(6) => 
        N_50_i_0, A_DIN(5) => N_48_i_0, A_DIN(4) => N_46_i_0, 
        A_DIN(3) => N_44_i_0, A_DIN(2) => N_42_i_0, A_DIN(1) => 
        N_40_i_0, A_DIN(0) => N_38_i_0, A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a7_1[1]\, 
        A_WEN(0) => \wen_a7_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b7_1[1]\, 
        B_WEN(0) => \wen_b7_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block25_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(1), Y => \wen_a25_1[1]\);
    
    \readData_31_bm_RNO[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[21]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[19]\, D => \readData15[21]\, Y => 
        N_965);
    
    \readData_31_bm[8]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_954, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[8]_net_1\, D => N_858, Y => 
        \readData_31_bm[8]_net_1\);
    
    block17_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(1), Y => 
        \wen_a17_1[1]\);
    
    \readData_31_am[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_490, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[24]_net_1\, D => N_394, Y => 
        \readData_31_am[24]_net_1\);
    
    \readData_31_am_RNO[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[32]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[29]\, D => \readData14[32]\, Y => 
        N_495);
    
    \readData_31_bm_RNO_1[16]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[18]\, D => \readData7[18]\, Y => 
        \readData_28_1_1[16]\);
    
    \readData_31_bm_1_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_727, D => N_631, Y => \readData_31_bm_1_1[5]_net_1\);
    
    \readData_31_am_1_1_RNO_0[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[22]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[20]\, D => \readData8[22]\, Y => 
        N_166);
    
    \readData_31_am_1_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_246, D => N_150, Y => \readData_31_am_1_1[4]_net_1\);
    
    block24 : RAM1K18
      port map(A_DOUT(17) => nc29, A_DOUT(16) => \readData24[16]\, 
        A_DOUT(15) => \readData24[15]\, A_DOUT(14) => 
        \readData24[14]\, A_DOUT(13) => \readData24[13]\, 
        A_DOUT(12) => \readData24[12]\, A_DOUT(11) => 
        \readData24[11]\, A_DOUT(10) => \readData24[10]\, 
        A_DOUT(9) => \readData24[9]\, A_DOUT(8) => nc88, 
        A_DOUT(7) => \readData24[7]\, A_DOUT(6) => 
        \readData24[6]\, A_DOUT(5) => \readData24[5]\, A_DOUT(4)
         => \readData24[4]\, A_DOUT(3) => \readData24[3]\, 
        A_DOUT(2) => \readData24[2]\, A_DOUT(1) => 
        \readData24[1]\, A_DOUT(0) => \readData24[0]\, B_DOUT(17)
         => nc53, B_DOUT(16) => \readData24[34]\, B_DOUT(15) => 
        \readData24[33]\, B_DOUT(14) => \readData24[32]\, 
        B_DOUT(13) => \readData24[31]\, B_DOUT(12) => 
        \readData24[30]\, B_DOUT(11) => \readData24[29]\, 
        B_DOUT(10) => \readData24[28]\, B_DOUT(9) => 
        \readData24[27]\, B_DOUT(8) => nc39, B_DOUT(7) => 
        \readData24[25]\, B_DOUT(6) => \readData24[24]\, 
        B_DOUT(5) => \readData24[23]\, B_DOUT(4) => 
        \readData24[22]\, B_DOUT(3) => \readData24[21]\, 
        B_DOUT(2) => \readData24[20]\, B_DOUT(1) => 
        \readData24[19]\, B_DOUT(0) => \readData24[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a24_1[1]\, A_WEN(0) => \wen_a24_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b24_1[1]\, 
        B_WEN(0) => \wen_b24_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_2[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[21]\, D => \readData3[21]\, Y => 
        \readData_25_1_1[19]\);
    
    \readData_31_bm_1_1_RNO_1[5]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[5]\, D => \readData5[5]\, Y => 
        \readData_21_1_1[5]\);
    
    \readData_31_am[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_484, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[18]_net_1\, D => N_388, Y => 
        \readData_31_am[18]_net_1\);
    
    \readData_31_bm[29]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_975, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[29]_net_1\, D => N_879, Y => 
        \readData_31_bm[29]_net_1\);
    
    \readData_31_bm_1_1_RNO_2[0]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[0]\, D => \readData1[0]\, Y => 
        \readData_18_1_1[0]\);
    
    \readData_31_am_RNO_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[30]\, D => \readData6[30]\, Y => 
        \readData_13_1_1[27]\);
    
    \readData_31_ns[8]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[8]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[8]_net_1\, Y => 
        ram_rdata(8));
    
    \readData_31_am_1_1_RNO[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[5]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[5]\, D => \readData12[5]\, Y => N_247);
    
    block8_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1143, D => sram_wen_mem(0), Y => \wen_a8_1[0]\);
    
    \readData_31_bm_RNO_1[19]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[21]\, D => \readData7[21]\, Y => 
        \readData_28_1_1[19]\);
    
    \readData_31_ns[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[2]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[2]_net_1\, Y => 
        ram_rdata(2));
    
    \readData_31_bm_1_1_RNO_1[7]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[7]\, D => \readData5[7]\, Y => 
        \readData_21_1_1[7]\);
    
    block18_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(14), C
         => readdata_xhdl1401_1, D => sram_wen_mem(0), Y => 
        \wen_a18_1[0]\);
    
    \readData_31_am[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_488, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[22]_net_1\, D => N_392, Y => 
        \readData_31_am[22]_net_1\);
    
    \readData_31_bm_RNO_0[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[20]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[18]\, D => \readData11[20]\, Y => 
        N_868);
    
    \readData_31_bm_1_1_RNO_2[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData17[27]\, D => \readData1[27]\, Y => 
        \readData_18_1_1[24]\);
    
    \readData_31_am_1_1_RNO[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[27]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[24]\, D => \readData12[27]\, Y => 
        N_266);
    
    \readData_31_am[10]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_476, B => ahbsram_addr(12), C => 
        \readData_31_am_1_1[10]_net_1\, D => N_380, Y => 
        \readData_31_am[10]_net_1\);
    
    \readData_31_am_RNO_1[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[31]\, D => \readData6[31]\, Y => 
        \readData_13_1_1[28]\);
    
    \readData_31_am_RNO_2[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[33]\, D => \readData2[33]\, Y => 
        \readData_10_1_1[30]\);
    
    block25 : RAM1K18
      port map(A_DOUT(17) => nc8, A_DOUT(16) => \readData25[16]\, 
        A_DOUT(15) => \readData25[15]\, A_DOUT(14) => 
        \readData25[14]\, A_DOUT(13) => \readData25[13]\, 
        A_DOUT(12) => \readData25[12]\, A_DOUT(11) => 
        \readData25[11]\, A_DOUT(10) => \readData25[10]\, 
        A_DOUT(9) => \readData25[9]\, A_DOUT(8) => nc82, 
        A_DOUT(7) => \readData25[7]\, A_DOUT(6) => 
        \readData25[6]\, A_DOUT(5) => \readData25[5]\, A_DOUT(4)
         => \readData25[4]\, A_DOUT(3) => \readData25[3]\, 
        A_DOUT(2) => \readData25[2]\, A_DOUT(1) => 
        \readData25[1]\, A_DOUT(0) => \readData25[0]\, B_DOUT(17)
         => nc108, B_DOUT(16) => \readData25[34]\, B_DOUT(15) => 
        \readData25[33]\, B_DOUT(14) => \readData25[32]\, 
        B_DOUT(13) => \readData25[31]\, B_DOUT(12) => 
        \readData25[30]\, B_DOUT(11) => \readData25[29]\, 
        B_DOUT(10) => \readData25[28]\, B_DOUT(9) => 
        \readData25[27]\, B_DOUT(8) => nc81, B_DOUT(7) => 
        \readData25[25]\, B_DOUT(6) => \readData25[24]\, 
        B_DOUT(5) => \readData25[23]\, B_DOUT(4) => 
        \readData25[22]\, B_DOUT(3) => \readData25[21]\, 
        B_DOUT(2) => \readData25[20]\, B_DOUT(1) => 
        \readData25[19]\, B_DOUT(0) => \readData25[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a25_1[1]\, A_WEN(0) => \wen_a25_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b25_1[1]\, 
        B_WEN(0) => \wen_b25_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    block1_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1419_0_a2_0, D => sram_wen_mem_m3(2), Y
         => \wen_b1_1[0]\);
    
    \readData_31_bm_RNO_0[23]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[25]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[23]\, D => \readData11[25]\, Y => 
        N_873);
    
    \readData_31_am_1_1[14]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_256, D => N_160, Y => 
        \readData_31_am_1_1[14]_net_1\);
    
    block6_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1144, D => sram_wen_mem(0), Y => \wen_a6_1[0]\);
    
    \readData_31_bm_1_1_RNO[3]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[3]\, B => ahbsram_addr(14), C => 
        \readData_21_1_1[3]\, D => \readData13[3]\, Y => N_725);
    
    \readData_31_am_1_1_RNO_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[29]\, D => \readData4[29]\, Y => 
        \readData_6_1_1[26]\);
    
    \readData_31_bm_RNO_0[20]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[22]\, B => ahbsram_addr(14), C
         => \readData_25_1_1[20]\, D => \readData11[22]\, Y => 
        N_870);
    
    \readData_31_bm[22]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_968, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[22]_net_1\, D => N_872, Y => 
        \readData_31_bm[22]_net_1\);
    
    \readData_31_am_1_1[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_262, D => N_166, Y => 
        \readData_31_am_1_1[20]_net_1\);
    
    block19_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem(1), Y => \wen_a19_1[1]\);
    
    \readData_31_am_1_1_RNO_2[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[14]\, D => \readData0[14]\, Y => 
        \readData_3_1_1[13]\);
    
    block21_RNO_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(1), Y => \wen_a21_1[1]\);
    
    block16 : RAM1K18
      port map(A_DOUT(17) => nc79, A_DOUT(16) => \readData16[16]\, 
        A_DOUT(15) => \readData16[15]\, A_DOUT(14) => 
        \readData16[14]\, A_DOUT(13) => \readData16[13]\, 
        A_DOUT(12) => \readData16[12]\, A_DOUT(11) => 
        \readData16[11]\, A_DOUT(10) => \readData16[10]\, 
        A_DOUT(9) => \readData16[9]\, A_DOUT(8) => nc43, 
        A_DOUT(7) => \readData16[7]\, A_DOUT(6) => 
        \readData16[6]\, A_DOUT(5) => \readData16[5]\, A_DOUT(4)
         => \readData16[4]\, A_DOUT(3) => \readData16[3]\, 
        A_DOUT(2) => \readData16[2]\, A_DOUT(1) => 
        \readData16[1]\, A_DOUT(0) => \readData16[0]\, B_DOUT(17)
         => nc69, B_DOUT(16) => \readData16[34]\, B_DOUT(15) => 
        \readData16[33]\, B_DOUT(14) => \readData16[32]\, 
        B_DOUT(13) => \readData16[31]\, B_DOUT(12) => 
        \readData16[30]\, B_DOUT(11) => \readData16[29]\, 
        B_DOUT(10) => \readData16[28]\, B_DOUT(9) => 
        \readData16[27]\, B_DOUT(8) => nc56, B_DOUT(7) => 
        \readData16[25]\, B_DOUT(6) => \readData16[24]\, 
        B_DOUT(5) => \readData16[23]\, B_DOUT(4) => 
        \readData16[22]\, B_DOUT(3) => \readData16[21]\, 
        B_DOUT(2) => \readData16[20]\, B_DOUT(1) => 
        \readData16[19]\, B_DOUT(0) => \readData16[18]\, BUSY => 
        OPEN, A_CLK => CertificationSystem_sb_0_FAB_CCC_GL0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_375_i_0, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => N_72_i_0, A_DIN(15) => N_70_i_0, 
        A_DIN(14) => N_68_i_0, A_DIN(13) => N_66_i_0, A_DIN(12)
         => N_64_i_0, A_DIN(11) => N_58_i_0, A_DIN(10) => 
        N_56_i_0, A_DIN(9) => N_54_i_0, A_DIN(8) => GND_net_1, 
        A_DIN(7) => N_52_i_0, A_DIN(6) => N_50_i_0, A_DIN(5) => 
        N_48_i_0, A_DIN(4) => N_46_i_0, A_DIN(3) => N_44_i_0, 
        A_DIN(2) => N_42_i_0, A_DIN(1) => N_40_i_0, A_DIN(0) => 
        N_38_i_0, A_ADDR(13) => ahbsram_addr(10), A_ADDR(12) => 
        ahbsram_addr(9), A_ADDR(11) => ahbsram_addr(8), 
        A_ADDR(10) => ahbsram_addr(7), A_ADDR(9) => 
        ahbsram_addr(6), A_ADDR(8) => ahbsram_addr(5), A_ADDR(7)
         => ahbsram_addr(4), A_ADDR(6) => ahbsram_addr(3), 
        A_ADDR(5) => ahbsram_addr(2), A_ADDR(4) => GND_net_1, 
        A_ADDR(3) => GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1)
         => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1) => 
        \wen_a16_1[1]\, A_WEN(0) => \wen_a16_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b16_1[1]\, 
        B_WEN(0) => \wen_b16_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_1_1_RNO[9]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[10]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[9]\, D => \readData13[10]\, Y => 
        N_731);
    
    \readData_31_bm[11]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_957, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[11]_net_1\, D => N_861, Y => 
        \readData_31_bm[11]_net_1\);
    
    \readData_31_am_1_1_RNO_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[14]\, D => \readData4[14]\, Y => 
        \readData_6_1_1[13]\);
    
    \readData_31_bm_1_1_RNO[17]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[19]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[17]\, D => \readData13[19]\, Y => 
        N_739);
    
    \readData_31_bm_1_1[23]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_745, D => N_649, Y => 
        \readData_31_bm_1_1[23]_net_1\);
    
    \readData_31_bm_1_1[12]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_734, D => N_638, Y => 
        \readData_31_bm_1_1[12]_net_1\);
    
    \readData_31_am_1_1_RNO_2[20]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[22]\, D => \readData0[22]\, Y => 
        \readData_3_1_1[20]\);
    
    \readData_31_am_1_1_RNO[2]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[2]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[2]\, D => \readData12[2]\, Y => N_244);
    
    \readData_31_bm_1_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_728, D => N_632, Y => \readData_31_bm_1_1[6]_net_1\);
    
    block4_RNO_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem(1), Y => \wen_a4_1[1]\);
    
    block16_RNO : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem(0), Y => 
        \wen_a16_1[0]\);
    
    \readData_31_bm_RNO_2[28]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[31]\, D => \readData3[31]\, Y => 
        \readData_25_1_1[28]\);
    
    \readData_31_bm_RNO_2[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[14]\, D => \readData3[14]\, Y => 
        \readData_25_1_1[13]\);
    
    \readData_31_bm[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_976, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[30]_net_1\, D => N_880, Y => 
        \readData_31_bm[30]_net_1\);
    
    block9 : RAM1K18
      port map(A_DOUT(17) => nc20, A_DOUT(16) => \readData9[16]\, 
        A_DOUT(15) => \readData9[15]\, A_DOUT(14) => 
        \readData9[14]\, A_DOUT(13) => \readData9[13]\, 
        A_DOUT(12) => \readData9[12]\, A_DOUT(11) => 
        \readData9[11]\, A_DOUT(10) => \readData9[10]\, A_DOUT(9)
         => \readData9[9]\, A_DOUT(8) => nc10, A_DOUT(7) => 
        \readData9[7]\, A_DOUT(6) => \readData9[6]\, A_DOUT(5)
         => \readData9[5]\, A_DOUT(4) => \readData9[4]\, 
        A_DOUT(3) => \readData9[3]\, A_DOUT(2) => \readData9[2]\, 
        A_DOUT(1) => \readData9[1]\, A_DOUT(0) => \readData9[0]\, 
        B_DOUT(17) => nc57, B_DOUT(16) => \readData9[34]\, 
        B_DOUT(15) => \readData9[33]\, B_DOUT(14) => 
        \readData9[32]\, B_DOUT(13) => \readData9[31]\, 
        B_DOUT(12) => \readData9[30]\, B_DOUT(11) => 
        \readData9[29]\, B_DOUT(10) => \readData9[28]\, B_DOUT(9)
         => \readData9[27]\, B_DOUT(8) => nc95, B_DOUT(7) => 
        \readData9[25]\, B_DOUT(6) => \readData9[24]\, B_DOUT(5)
         => \readData9[23]\, B_DOUT(4) => \readData9[22]\, 
        B_DOUT(3) => \readData9[21]\, B_DOUT(2) => 
        \readData9[20]\, B_DOUT(1) => \readData9[19]\, B_DOUT(0)
         => \readData9[18]\, BUSY => OPEN, A_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => N_375_i_0, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        N_72_i_0, A_DIN(15) => N_70_i_0, A_DIN(14) => N_68_i_0, 
        A_DIN(13) => N_66_i_0, A_DIN(12) => N_64_i_0, A_DIN(11)
         => N_58_i_0, A_DIN(10) => N_56_i_0, A_DIN(9) => N_54_i_0, 
        A_DIN(8) => GND_net_1, A_DIN(7) => N_52_i_0, A_DIN(6) => 
        N_50_i_0, A_DIN(5) => N_48_i_0, A_DIN(4) => N_46_i_0, 
        A_DIN(3) => N_44_i_0, A_DIN(2) => N_42_i_0, A_DIN(1) => 
        N_40_i_0, A_DIN(0) => N_38_i_0, A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a9_1[1]\, 
        A_WEN(0) => \wen_a9_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b9_1[1]\, 
        B_WEN(0) => \wen_b9_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_bm_RNO_2[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData19[11]\, D => \readData3[11]\, Y => 
        \readData_25_1_1[10]\);
    
    \readData_31_am_1_1_RNO_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData20[4]\, D => \readData4[4]\, Y => 
        \readData_6_1_1[4]\);
    
    \readData_31_am_RNO_0[5]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData26[5]\, B => ahbsram_addr(14), C => 
        \readData_10_1_1[5]\, D => \readData10[5]\, Y => N_375);
    
    \readData_31_am_1_1[27]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_269, D => N_173, Y => 
        \readData_31_am_1_1[27]_net_1\);
    
    \readData_31_bm_1_1_RNO_0[13]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[14]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[13]\, D => \readData9[14]\, Y => 
        N_639);
    
    \readData_31_bm_RNO_1[13]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[14]\, D => \readData7[14]\, Y => 
        \readData_28_1_1[13]\);
    
    block17_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem_m3(3), Y => 
        \wen_b17_1[1]\);
    
    \readData_31_bm_RNO_1[4]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[4]\, D => \readData7[4]\, Y => 
        \readData_28_1_1[4]\);
    
    \readData_31_am_1_1_RNO_0[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[34]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[31]\, D => \readData8[34]\, Y => 
        N_177);
    
    block21_RNO_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1150, D => sram_wen_mem_m3(3), Y => \wen_b_m[1]\);
    
    \readData_31_am_1_1[30]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_272, D => N_176, Y => 
        \readData_31_am_1_1[30]_net_1\);
    
    \readData_31_bm_RNO_1[10]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[11]\, D => \readData7[11]\, Y => 
        \readData_28_1_1[10]\);
    
    \readData_31_am_1_1_RNO_0[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[6]\, B => ahbsram_addr(14), C => 
        \readData_3_1_1[6]\, D => \readData8[6]\, Y => N_152);
    
    \readData_31_bm_1_1_RNO_0[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[33]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[30]\, D => \readData9[33]\, Y => 
        N_656);
    
    \readData_31_bm[0]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_946, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[0]_net_1\, D => N_850, Y => 
        \readData_31_bm[0]_net_1\);
    
    \readData_31_bm_RNO_1[6]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData23[6]\, D => \readData7[6]\, Y => 
        \readData_28_1_1[6]\);
    
    \readData_31_am_1_1_RNO[4]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[4]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[4]\, D => \readData12[4]\, Y => N_246);
    
    block17_RNO_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => readdata_xhdl1403_0, D => sram_wen_mem_m3(2), Y => 
        \wen_b17_1[0]\);
    
    \readData_31_bm_RNO_0[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData27[7]\, B => ahbsram_addr(14), C => 
        \readData_25_1_1[7]\, D => \readData11[7]\, Y => N_857);
    
    \readData_31_bm_1_1_RNO[27]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[30]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[27]\, D => \readData13[30]\, Y => 
        N_749);
    
    \readData_31_am_1_1_RNO_0[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[21]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[19]\, D => \readData8[21]\, Y => 
        N_165);
    
    \readData_31_bm_1_1_RNO_0[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[34]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[31]\, D => \readData9[34]\, Y => 
        N_657);
    
    \readData_31_am_1_1_RNO[6]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[6]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[6]\, D => \readData12[6]\, Y => N_248);
    
    block30_RNO_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1148, D => sram_wen_mem_m3(3), Y => \wen_b30_1[1]\);
    
    \readData_31_bm_1_1_RNO[30]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData29[33]\, B => ahbsram_addr(14), C
         => \readData_21_1_1[30]\, D => \readData13[33]\, Y => 
        N_752);
    
    block3 : RAM1K18
      port map(A_DOUT(17) => nc24, A_DOUT(16) => \readData3[16]\, 
        A_DOUT(15) => \readData3[15]\, A_DOUT(14) => 
        \readData3[14]\, A_DOUT(13) => \readData3[13]\, 
        A_DOUT(12) => \readData3[12]\, A_DOUT(11) => 
        \readData3[11]\, A_DOUT(10) => \readData3[10]\, A_DOUT(9)
         => \readData3[9]\, A_DOUT(8) => nc14, A_DOUT(7) => 
        \readData3[7]\, A_DOUT(6) => \readData3[6]\, A_DOUT(5)
         => \readData3[5]\, A_DOUT(4) => \readData3[4]\, 
        A_DOUT(3) => \readData3[3]\, A_DOUT(2) => \readData3[2]\, 
        A_DOUT(1) => \readData3[1]\, A_DOUT(0) => \readData3[0]\, 
        B_DOUT(17) => nc46, B_DOUT(16) => \readData3[34]\, 
        B_DOUT(15) => \readData3[33]\, B_DOUT(14) => 
        \readData3[32]\, B_DOUT(13) => \readData3[31]\, 
        B_DOUT(12) => \readData3[30]\, B_DOUT(11) => 
        \readData3[29]\, B_DOUT(10) => \readData3[28]\, B_DOUT(9)
         => \readData3[27]\, B_DOUT(8) => nc30, B_DOUT(7) => 
        \readData3[25]\, B_DOUT(6) => \readData3[24]\, B_DOUT(5)
         => \readData3[23]\, B_DOUT(4) => \readData3[22]\, 
        B_DOUT(3) => \readData3[21]\, B_DOUT(2) => 
        \readData3[20]\, B_DOUT(1) => \readData3[19]\, B_DOUT(0)
         => \readData3[18]\, BUSY => OPEN, A_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => MSS_READY, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => N_375_i_0, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        N_72_i_0, A_DIN(15) => N_70_i_0, A_DIN(14) => N_68_i_0, 
        A_DIN(13) => N_66_i_0, A_DIN(12) => N_64_i_0, A_DIN(11)
         => N_58_i_0, A_DIN(10) => N_56_i_0, A_DIN(9) => N_54_i_0, 
        A_DIN(8) => GND_net_1, A_DIN(7) => N_52_i_0, A_DIN(6) => 
        N_50_i_0, A_DIN(5) => N_48_i_0, A_DIN(4) => N_46_i_0, 
        A_DIN(3) => N_44_i_0, A_DIN(2) => N_42_i_0, A_DIN(1) => 
        N_40_i_0, A_DIN(0) => N_38_i_0, A_ADDR(13) => 
        ahbsram_addr(10), A_ADDR(12) => ahbsram_addr(9), 
        A_ADDR(11) => ahbsram_addr(8), A_ADDR(10) => 
        ahbsram_addr(7), A_ADDR(9) => ahbsram_addr(6), A_ADDR(8)
         => ahbsram_addr(5), A_ADDR(7) => ahbsram_addr(4), 
        A_ADDR(6) => ahbsram_addr(3), A_ADDR(5) => 
        ahbsram_addr(2), A_ADDR(4) => GND_net_1, A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => \wen_a3_1[1]\, 
        A_WEN(0) => \wen_a3_1[0]\, B_CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => MSS_READY, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        N_63_i_0, B_DIN(15) => N_62_i_0, B_DIN(14) => N_60_i_0, 
        B_DIN(13) => N_98_i_0, B_DIN(12) => N_96_i_0, B_DIN(11)
         => N_94_i_0, B_DIN(10) => N_92_i_0, B_DIN(9) => N_90_i_0, 
        B_DIN(8) => GND_net_1, B_DIN(7) => N_88_i_0, B_DIN(6) => 
        N_86_i_0, B_DIN(5) => N_84_i_0, B_DIN(4) => N_82_i_0, 
        B_DIN(3) => N_80_i_0, B_DIN(2) => N_78_i_0, B_DIN(1) => 
        N_76_i_0, B_DIN(0) => N_74_i_0, B_ADDR(13) => 
        ahbsram_addr(10), B_ADDR(12) => ahbsram_addr(9), 
        B_ADDR(11) => ahbsram_addr(8), B_ADDR(10) => 
        ahbsram_addr(7), B_ADDR(9) => ahbsram_addr(6), B_ADDR(8)
         => ahbsram_addr(5), B_ADDR(7) => ahbsram_addr(4), 
        B_ADDR(6) => ahbsram_addr(3), B_ADDR(5) => 
        ahbsram_addr(2), B_ADDR(4) => GND_net_1, B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => \wen_b3_1[1]\, 
        B_WEN(0) => \wen_b3_1[0]\, A_EN => VCC_net_1, A_DOUT_LAT
         => VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, 
        B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2)
         => VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \readData_31_ns[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[0]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[0]_net_1\, Y => 
        ram_rdata(0));
    
    \readData_31_am_1_1_RNO[31]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[34]\, B => ahbsram_addr(14), C
         => \readData_6_1_1[31]\, D => \readData12[34]\, Y => 
        N_273);
    
    \readData_31_bm_1_1_RNO_0[19]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData25[21]\, B => ahbsram_addr(14), C
         => \readData_18_1_1[19]\, D => \readData9[21]\, Y => 
        N_645);
    
    \readData_31_bm[7]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => N_953, B => ahbsram_addr(12), C => 
        \readData_31_bm_1_1[7]_net_1\, D => N_857, Y => 
        \readData_31_bm[7]_net_1\);
    
    \readData_31_am_RNO_2[2]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData18[2]\, D => \readData2[2]\, Y => 
        \readData_10_1_1[2]\);
    
    \readData_31_bm_1_1_RNO_1[24]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData21[27]\, D => \readData5[27]\, Y => 
        \readData_21_1_1[24]\);
    
    \readData_31_bm_RNO[14]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData31[15]\, B => ahbsram_addr(14), C
         => \readData_28_1_1[14]\, D => \readData15[15]\, Y => 
        N_960);
    
    \readData_31_am_RNO_1[9]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData22[10]\, D => \readData6[10]\, Y => 
        \readData_13_1_1[9]\);
    
    \readData_31_bm_1_1[18]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_740, D => N_644, Y => 
        \readData_31_bm_1_1[18]_net_1\);
    
    \readData_31_am_1_1[3]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_245, D => N_149, Y => \readData_31_am_1_1[3]_net_1\);
    
    \readData_31_am_1_1_RNO_2[8]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(15), B => ahbsram_addr(14), C
         => \readData16[9]\, D => \readData0[9]\, Y => 
        \readData_3_1_1[8]\);
    
    \readData_31_am_1_1_RNO_0[24]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[27]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[24]\, D => \readData8[27]\, Y => 
        N_170);
    
    \readData_31_bm_1_1[26]\ : CFG4
      generic map(INIT => x"4657")

      port map(A => ahbsram_addr(13), B => ahbsram_addr(12), C
         => N_748, D => N_652, Y => 
        \readData_31_bm_1_1[26]_net_1\);
    
    \wen_a_m_12_0_a2_0[1]\ : CFG3
      generic map(INIT => x"08")

      port map(A => ahbsram_addr(12), B => ahbsram_addr(14), C
         => ahbsram_addr(13), Y => N_1147);
    
    block29_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1149, D => sram_wen_mem(0), Y => \wen_a29_1[0]\);
    
    block3_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => ahbsram_addr(11), B => ahbsram_addr(15), C
         => N_1168, D => sram_wen_mem_m3(2), Y => \wen_b3_1[0]\);
    
    \readData_31_ns[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \readData_31_am[3]_net_1\, B => 
        ahbsram_addr(11), C => \readData_31_bm[3]_net_1\, Y => 
        ram_rdata(3));
    
    \readData_31_am_1_1_RNO_0[25]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData24[28]\, B => ahbsram_addr(14), C
         => \readData_3_1_1[25]\, D => \readData8[28]\, Y => 
        N_171);
    
    \readData_31_am_1_1_RNO[1]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData28[1]\, B => ahbsram_addr(14), C => 
        \readData_6_1_1[1]\, D => \readData12[1]\, Y => N_243);
    
    \readData_31_am_RNO[18]\ : CFG4
      generic map(INIT => x"CB0B")

      port map(A => \readData30[20]\, B => ahbsram_addr(14), C
         => \readData_13_1_1[18]\, D => \readData14[20]\, Y => 
        N_484);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf is

    port( CoreAHBLite_0_AHBmslave3_HRDATA      : out   std_logic_vector(31 downto 0);
          sramcurr_state                       : out   std_logic_vector(1 downto 0);
          ahbsram_size                         : in    std_logic_vector(1 downto 0);
          ahbcurr_state                        : in    std_logic_vector(1 downto 0);
          ahbsram_addr                         : in    std_logic_vector(15 downto 0);
          MSS_READY                            : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic;
          sram_done                            : out   std_logic;
          HWRITE_d                             : in    std_logic;
          ahbsram_req_d1                       : in    std_logic;
          N_38_i_0                             : in    std_logic;
          N_40_i_0                             : in    std_logic;
          N_42_i_0                             : in    std_logic;
          N_44_i_0                             : in    std_logic;
          N_46_i_0                             : in    std_logic;
          N_48_i_0                             : in    std_logic;
          N_50_i_0                             : in    std_logic;
          N_52_i_0                             : in    std_logic;
          N_54_i_0                             : in    std_logic;
          N_56_i_0                             : in    std_logic;
          N_58_i_0                             : in    std_logic;
          N_64_i_0                             : in    std_logic;
          N_66_i_0                             : in    std_logic;
          N_68_i_0                             : in    std_logic;
          N_70_i_0                             : in    std_logic;
          N_72_i_0                             : in    std_logic;
          N_74_i_0                             : in    std_logic;
          N_76_i_0                             : in    std_logic;
          N_78_i_0                             : in    std_logic;
          N_80_i_0                             : in    std_logic;
          N_82_i_0                             : in    std_logic;
          N_84_i_0                             : in    std_logic;
          N_86_i_0                             : in    std_logic;
          N_88_i_0                             : in    std_logic;
          N_90_i_0                             : in    std_logic;
          N_92_i_0                             : in    std_logic;
          N_94_i_0                             : in    std_logic;
          N_96_i_0                             : in    std_logic;
          N_98_i_0                             : in    std_logic;
          N_60_i_0                             : in    std_logic;
          N_62_i_0                             : in    std_logic;
          N_63_i_0                             : in    std_logic
        );

end CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf;

architecture DEF_ARCH of 
        CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component 
        CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8
    port( ram_rdata                            : out   std_logic_vector(31 downto 0);
          sram_wen_mem_m3                      : in    std_logic_vector(3 downto 2) := (others => 'U');
          sram_wen_mem                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          ahbsram_addr                         : in    std_logic_vector(15 downto 2) := (others => 'U');
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U';
          N_375_i_0                            : in    std_logic := 'U';
          N_38_i_0                             : in    std_logic := 'U';
          N_40_i_0                             : in    std_logic := 'U';
          N_42_i_0                             : in    std_logic := 'U';
          N_44_i_0                             : in    std_logic := 'U';
          N_46_i_0                             : in    std_logic := 'U';
          N_48_i_0                             : in    std_logic := 'U';
          N_50_i_0                             : in    std_logic := 'U';
          N_52_i_0                             : in    std_logic := 'U';
          N_54_i_0                             : in    std_logic := 'U';
          N_56_i_0                             : in    std_logic := 'U';
          N_58_i_0                             : in    std_logic := 'U';
          N_64_i_0                             : in    std_logic := 'U';
          N_66_i_0                             : in    std_logic := 'U';
          N_68_i_0                             : in    std_logic := 'U';
          N_70_i_0                             : in    std_logic := 'U';
          N_72_i_0                             : in    std_logic := 'U';
          N_74_i_0                             : in    std_logic := 'U';
          N_76_i_0                             : in    std_logic := 'U';
          N_78_i_0                             : in    std_logic := 'U';
          N_80_i_0                             : in    std_logic := 'U';
          N_82_i_0                             : in    std_logic := 'U';
          N_84_i_0                             : in    std_logic := 'U';
          N_86_i_0                             : in    std_logic := 'U';
          N_88_i_0                             : in    std_logic := 'U';
          N_90_i_0                             : in    std_logic := 'U';
          N_92_i_0                             : in    std_logic := 'U';
          N_94_i_0                             : in    std_logic := 'U';
          N_96_i_0                             : in    std_logic := 'U';
          N_98_i_0                             : in    std_logic := 'U';
          N_60_i_0                             : in    std_logic := 'U';
          N_62_i_0                             : in    std_logic := 'U';
          N_63_i_0                             : in    std_logic := 'U'
        );
  end component;

    signal VCC_net_1, \ram_rdata[20]\, \sram_ren_d\, GND_net_1, 
        \ram_rdata[21]\, \ram_rdata[22]\, \ram_rdata[23]\, 
        \ram_rdata[24]\, \ram_rdata[25]\, \ram_rdata[26]\, 
        \ram_rdata[27]\, \ram_rdata[28]\, \ram_rdata[29]\, 
        \ram_rdata[30]\, \ram_rdata[31]\, \ram_rdata[5]\, 
        \ram_rdata[6]\, \ram_rdata[7]\, \ram_rdata[8]\, 
        \ram_rdata[9]\, \ram_rdata[10]\, \ram_rdata[11]\, 
        \ram_rdata[12]\, \ram_rdata[13]\, \ram_rdata[14]\, 
        \ram_rdata[15]\, \ram_rdata[16]\, \ram_rdata[17]\, 
        \ram_rdata[18]\, \ram_rdata[19]\, \ram_rdata[0]\, 
        \ram_rdata[1]\, \ram_rdata[2]\, \ram_rdata[3]\, 
        \ram_rdata[4]\, \sramcurr_state[0]_net_1\, N_374_i_0, 
        \sramcurr_state[1]_net_1\, N_373_i_0, sram_done_net_1, 
        N_5_i_0, N_375_i_0, N_380, N_396, N_402, N_382, N_388, 
        N_385, \sram_wen_mem_m3[3]_net_1\, 
        \sram_wen_mem_m3[2]_net_1\, \sram_wen_mem[1]_net_1\, 
        \sram_wen_mem[0]_net_1\ : std_logic;

    for all : CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8
	Use entity work.
        CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8(DEF_ARCH);
begin 

    sramcurr_state(1) <= \sramcurr_state[1]_net_1\;
    sramcurr_state(0) <= \sramcurr_state[0]_net_1\;
    sram_done <= sram_done_net_1;

    \sramahb_rdata_xhdl2[25]\ : SLE
      port map(D => \ram_rdata[25]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(25));
    
    \sramahb_rdata_xhdl2[16]\ : SLE
      port map(D => \ram_rdata[16]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(16));
    
    \sram_wen_mem_m3_i_o4[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_382, B => N_380, Y => N_385);
    
    \sramahb_rdata_xhdl2[24]\ : SLE
      port map(D => \ram_rdata[24]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(24));
    
    \sram_wen_mem_m3[3]\ : CFG4
      generic map(INIT => x"080F")

      port map(A => ahbsram_addr(1), B => ahbsram_addr(0), C => 
        N_385, D => N_396, Y => \sram_wen_mem_m3[3]_net_1\);
    
    \sramahb_rdata_xhdl2[8]\ : SLE
      port map(D => \ram_rdata[8]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(8));
    
    sram_ren_1_sqmuxa_0_a2_i_o4 : CFG4
      generic map(INIT => x"FFF1")

      port map(A => ahbcurr_state(0), B => ahbcurr_state(1), C
         => HWRITE_d, D => ahbsram_req_d1, Y => N_388);
    
    \sramahb_rdata_xhdl2[13]\ : SLE
      port map(D => \ram_rdata[13]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(13));
    
    \sramahb_rdata_xhdl2[9]\ : SLE
      port map(D => \ram_rdata[9]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(9));
    
    \sramahb_rdata_xhdl2[2]\ : SLE
      port map(D => \ram_rdata[2]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(2));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sramahb_rdata_xhdl2[22]\ : SLE
      port map(D => \ram_rdata[22]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(22));
    
    \sram_wen_mem[0]\ : CFG4
      generic map(INIT => x"010F")

      port map(A => ahbsram_addr(1), B => ahbsram_addr(0), C => 
        N_385, D => N_402, Y => \sram_wen_mem[0]_net_1\);
    
    \sramahb_rdata_xhdl2[5]\ : SLE
      port map(D => \ram_rdata[5]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(5));
    
    \sramahb_rdata_xhdl2[19]\ : SLE
      port map(D => \ram_rdata[19]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(19));
    
    \sramahb_rdata_xhdl2[4]\ : SLE
      port map(D => \ram_rdata[4]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(4));
    
    \sramahb_rdata_xhdl2[21]\ : SLE
      port map(D => \ram_rdata[21]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(21));
    
    \sramahb_rdata_xhdl2[18]\ : SLE
      port map(D => \ram_rdata[18]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(18));
    
    \sramahb_rdata_xhdl2[20]\ : SLE
      port map(D => \ram_rdata[20]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(20));
    
    \sramahb_rdata_xhdl2[15]\ : SLE
      port map(D => \ram_rdata[15]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(15));
    
    \sramcurr_state[0]\ : SLE
      port map(D => N_374_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sramcurr_state[0]_net_1\);
    
    \sramahb_rdata_xhdl2[14]\ : SLE
      port map(D => \ram_rdata[14]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(14));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sram_done\ : SLE
      port map(D => N_5_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => sram_done_net_1);
    
    \sramahb_rdata_xhdl2[0]\ : SLE
      port map(D => \ram_rdata[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(0));
    
    sram_wen_mems2_i_a4 : CFG3
      generic map(INIT => x"51")

      port map(A => ahbsram_size(1), B => ahbsram_size(0), C => 
        ahbsram_addr(1), Y => N_402);
    
    sram_done_RNO : CFG4
      generic map(INIT => x"0302")

      port map(A => ahbcurr_state(0), B => ahbsram_req_d1, C => 
        N_380, D => ahbcurr_state(1), Y => N_5_i_0);
    
    \sramcurr_state_ns_1_0_.N_373_i\ : CFG4
      generic map(INIT => x"0407")

      port map(A => sram_done_net_1, B => 
        \sramcurr_state[1]_net_1\, C => \sramcurr_state[0]_net_1\, 
        D => N_388, Y => N_373_i_0);
    
    \sram_wen_mem_m3[2]\ : CFG4
      generic map(INIT => x"020F")

      port map(A => ahbsram_addr(1), B => ahbsram_addr(0), C => 
        N_385, D => N_396, Y => \sram_wen_mem_m3[2]_net_1\);
    
    \sramahb_rdata_xhdl2[27]\ : SLE
      port map(D => \ram_rdata[27]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(27));
    
    \S0.byte_0\ : 
        CertificationSystem_sb_COREAHBLSRAM_0_0_lsram_2048to139264x8
      port map(ram_rdata(31) => \ram_rdata[31]\, ram_rdata(30)
         => \ram_rdata[30]\, ram_rdata(29) => \ram_rdata[29]\, 
        ram_rdata(28) => \ram_rdata[28]\, ram_rdata(27) => 
        \ram_rdata[27]\, ram_rdata(26) => \ram_rdata[26]\, 
        ram_rdata(25) => \ram_rdata[25]\, ram_rdata(24) => 
        \ram_rdata[24]\, ram_rdata(23) => \ram_rdata[23]\, 
        ram_rdata(22) => \ram_rdata[22]\, ram_rdata(21) => 
        \ram_rdata[21]\, ram_rdata(20) => \ram_rdata[20]\, 
        ram_rdata(19) => \ram_rdata[19]\, ram_rdata(18) => 
        \ram_rdata[18]\, ram_rdata(17) => \ram_rdata[17]\, 
        ram_rdata(16) => \ram_rdata[16]\, ram_rdata(15) => 
        \ram_rdata[15]\, ram_rdata(14) => \ram_rdata[14]\, 
        ram_rdata(13) => \ram_rdata[13]\, ram_rdata(12) => 
        \ram_rdata[12]\, ram_rdata(11) => \ram_rdata[11]\, 
        ram_rdata(10) => \ram_rdata[10]\, ram_rdata(9) => 
        \ram_rdata[9]\, ram_rdata(8) => \ram_rdata[8]\, 
        ram_rdata(7) => \ram_rdata[7]\, ram_rdata(6) => 
        \ram_rdata[6]\, ram_rdata(5) => \ram_rdata[5]\, 
        ram_rdata(4) => \ram_rdata[4]\, ram_rdata(3) => 
        \ram_rdata[3]\, ram_rdata(2) => \ram_rdata[2]\, 
        ram_rdata(1) => \ram_rdata[1]\, ram_rdata(0) => 
        \ram_rdata[0]\, sram_wen_mem_m3(3) => 
        \sram_wen_mem_m3[3]_net_1\, sram_wen_mem_m3(2) => 
        \sram_wen_mem_m3[2]_net_1\, sram_wen_mem(1) => 
        \sram_wen_mem[1]_net_1\, sram_wen_mem(0) => 
        \sram_wen_mem[0]_net_1\, ahbsram_addr(15) => 
        ahbsram_addr(15), ahbsram_addr(14) => ahbsram_addr(14), 
        ahbsram_addr(13) => ahbsram_addr(13), ahbsram_addr(12)
         => ahbsram_addr(12), ahbsram_addr(11) => 
        ahbsram_addr(11), ahbsram_addr(10) => ahbsram_addr(10), 
        ahbsram_addr(9) => ahbsram_addr(9), ahbsram_addr(8) => 
        ahbsram_addr(8), ahbsram_addr(7) => ahbsram_addr(7), 
        ahbsram_addr(6) => ahbsram_addr(6), ahbsram_addr(5) => 
        ahbsram_addr(5), ahbsram_addr(4) => ahbsram_addr(4), 
        ahbsram_addr(3) => ahbsram_addr(3), ahbsram_addr(2) => 
        ahbsram_addr(2), CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, MSS_READY => 
        MSS_READY, N_375_i_0 => N_375_i_0, N_38_i_0 => N_38_i_0, 
        N_40_i_0 => N_40_i_0, N_42_i_0 => N_42_i_0, N_44_i_0 => 
        N_44_i_0, N_46_i_0 => N_46_i_0, N_48_i_0 => N_48_i_0, 
        N_50_i_0 => N_50_i_0, N_52_i_0 => N_52_i_0, N_54_i_0 => 
        N_54_i_0, N_56_i_0 => N_56_i_0, N_58_i_0 => N_58_i_0, 
        N_64_i_0 => N_64_i_0, N_66_i_0 => N_66_i_0, N_68_i_0 => 
        N_68_i_0, N_70_i_0 => N_70_i_0, N_72_i_0 => N_72_i_0, 
        N_74_i_0 => N_74_i_0, N_76_i_0 => N_76_i_0, N_78_i_0 => 
        N_78_i_0, N_80_i_0 => N_80_i_0, N_82_i_0 => N_82_i_0, 
        N_84_i_0 => N_84_i_0, N_86_i_0 => N_86_i_0, N_88_i_0 => 
        N_88_i_0, N_90_i_0 => N_90_i_0, N_92_i_0 => N_92_i_0, 
        N_94_i_0 => N_94_i_0, N_96_i_0 => N_96_i_0, N_98_i_0 => 
        N_98_i_0, N_60_i_0 => N_60_i_0, N_62_i_0 => N_62_i_0, 
        N_63_i_0 => N_63_i_0);
    
    \sramahb_rdata_xhdl2[26]\ : SLE
      port map(D => \ram_rdata[26]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(26));
    
    \sram_wen_mem_m3_i_o3[0]\ : CFG4
      generic map(INIT => x"FF1F")

      port map(A => ahbcurr_state(0), B => ahbcurr_state(1), C
         => HWRITE_d, D => ahbsram_req_d1, Y => N_382);
    
    \sramcurr_state_ns_1_0_.N_374_i\ : CFG4
      generic map(INIT => x"1013")

      port map(A => sram_done_net_1, B => 
        \sramcurr_state[1]_net_1\, C => \sramcurr_state[0]_net_1\, 
        D => N_382, Y => N_374_i_0);
    
    \sramahb_rdata_xhdl2[12]\ : SLE
      port map(D => \ram_rdata[12]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(12));
    
    \sramahb_rdata_xhdl2[31]\ : SLE
      port map(D => \ram_rdata[31]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(31));
    
    \sramahb_rdata_xhdl2[23]\ : SLE
      port map(D => \ram_rdata[23]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(23));
    
    \sramahb_rdata_xhdl2[30]\ : SLE
      port map(D => \ram_rdata[30]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(30));
    
    \sram_wen_mem[1]\ : CFG4
      generic map(INIT => x"040F")

      port map(A => ahbsram_addr(1), B => ahbsram_addr(0), C => 
        N_385, D => N_402, Y => \sram_wen_mem[1]_net_1\);
    
    sram_ren_d : SLE
      port map(D => N_375_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sram_ren_d\);
    
    \sramahb_rdata_xhdl2[11]\ : SLE
      port map(D => \ram_rdata[11]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(11));
    
    sram_ren_0_sqmuxa_0_a2_i_o4_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \sramcurr_state[0]_net_1\, B => 
        \sramcurr_state[1]_net_1\, Y => N_380);
    
    \sramahb_rdata_xhdl2[10]\ : SLE
      port map(D => \ram_rdata[10]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(10));
    
    \sramcurr_state[1]\ : SLE
      port map(D => N_373_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sramcurr_state[1]_net_1\);
    
    \sramahb_rdata_xhdl2[6]\ : SLE
      port map(D => \ram_rdata[6]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(6));
    
    \sramahb_rdata_xhdl2[7]\ : SLE
      port map(D => \ram_rdata[7]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(7));
    
    \sramahb_rdata_xhdl2[1]\ : SLE
      port map(D => \ram_rdata[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(1));
    
    \sramahb_rdata_xhdl2[29]\ : SLE
      port map(D => \ram_rdata[29]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(29));
    
    \sramahb_rdata_xhdl2[28]\ : SLE
      port map(D => \ram_rdata[28]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(28));
    
    \sramahb_rdata_xhdl2[17]\ : SLE
      port map(D => \ram_rdata[17]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(17));
    
    sram_ren_1_sqmuxa_0_a2_i_o4_RNIIG8E : CFG2
      generic map(INIT => x"1")

      port map(A => N_388, B => N_380, Y => N_375_i_0);
    
    \sramahb_rdata_xhdl2[3]\ : SLE
      port map(D => \ram_rdata[3]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \sram_ren_d\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAHBLite_0_AHBmslave3_HRDATA(3));
    
    sram_wen_mem_ss3_i_0_a4 : CFG3
      generic map(INIT => x"15")

      port map(A => ahbsram_size(1), B => ahbsram_size(0), C => 
        ahbsram_addr(1), Y => N_396);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf is

    port( ahbsram_size                                            : out   std_logic_vector(1 downto 0);
          CoreAHBLite_0_AHBmslave3_HADDR                          : in    std_logic_vector(11 to 11);
          ahbsram_addr                                            : out   std_logic_vector(15 downto 0);
          ahbcurr_state                                           : out   std_logic_vector(1 downto 0);
          sramcurr_state                                          : in    std_logic_vector(1 downto 0);
          arbRegSMCurrentState                                    : in    std_logic_vector(15 to 15);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP : in    std_logic_vector(0 to 0);
          xhdl1222_2                                              : in    std_logic;
          xhdl1222_0                                              : in    std_logic;
          SDATASELInt_9                                           : in    std_logic;
          SDATASELInt_8                                           : in    std_logic;
          SDATASELInt_7                                           : in    std_logic;
          SDATASELInt_6                                           : in    std_logic;
          SDATASELInt_13                                          : in    std_logic;
          SDATASELInt_12                                          : in    std_logic;
          SDATASELInt_11                                          : in    std_logic;
          SDATASELInt_10                                          : in    std_logic;
          SDATASELInt_4                                           : in    std_logic;
          SDATASELInt_2                                           : in    std_logic;
          SDATASELInt_1                                           : in    std_logic;
          SDATASELInt_0                                           : in    std_logic;
          MSS_READY                                               : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                    : in    std_logic;
          N_236                                                   : in    std_logic;
          N_271                                                   : out   std_logic;
          N_235                                                   : in    std_logic;
          N_246                                                   : in    std_logic;
          N_276                                                   : in    std_logic;
          N_194_i_0                                               : in    std_logic;
          N_195_i_0                                               : in    std_logic;
          N_196_i_0                                               : in    std_logic;
          N_259                                                   : in    std_logic;
          N_258                                                   : in    std_logic;
          N_257                                                   : in    std_logic;
          N_256                                                   : in    std_logic;
          N_255                                                   : in    std_logic;
          N_244                                                   : in    std_logic;
          N_243                                                   : in    std_logic;
          N_242                                                   : in    std_logic;
          N_241                                                   : in    std_logic;
          N_247                                                   : in    std_logic;
          HWRITE_d                                                : out   std_logic;
          N_277                                                   : in    std_logic;
          ahbsram_req_d1                                          : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                     : out   std_logic;
          sram_done                                               : in    std_logic;
          hready_m_xhdl343_11                                     : in    std_logic;
          N_305                                                   : out   std_logic;
          hready_m_xhdl343_10                                     : in    std_logic;
          hready_m_xhdl344_7                                      : in    std_logic;
          N_335                                                   : out   std_logic;
          N_215                                                   : out   std_logic;
          N_216                                                   : out   std_logic;
          N_214                                                   : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                 : out   std_logic;
          N_157_i_i_o2_0                                          : in    std_logic;
          N_157_i_i_o2_0_out                                      : in    std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY              : in    std_logic;
          defSlaveSMNextState                                     : in    std_logic;
          hready_m_xhdl345                                        : in    std_logic;
          un8_hreadyin_i_0                                        : out   std_logic;
          N_225                                                   : in    std_logic;
          HTRANS_i_a2_0_0                                         : in    std_logic;
          N_120                                                   : in    std_logic;
          hsel2_i_4                                               : in    std_logic
        );

end CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf;

architecture DEF_ARCH of 
        CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \count[3]_net_1\, VCC_net_1, N_57_i_i_0, counte, 
        GND_net_1, \count[4]_net_1\, N_368_i_0, \count[1]_net_1\, 
        N_370_i_0, \count[2]_net_1\, N_928_i_0, \count[0]_net_1\, 
        N_400, \N_271\, \burst_count_reg[0]_net_1\, N_113_i_0, 
        \ahbcurr_state[1]_net_1\, \ahbcurr_state_ns[1]\, 
        \ahbcurr_state[0]_net_1\, \ahbcurr_state_ns[0]\, 
        ahbsram_req_d1_net_1, 
        \CoreAHBLite_0_AHBmslave3_HREADY_i_1\, m9_0_1, 
        \un8_hreadyin_i_1\, N_378, un1_sramahb_ack_i_i_0_o3_1, 
        N_381, m6_0_a4_0_0, N_408, N_391, N_403, 
        un8_hreadyin_i_0_net_1, \un8_hreadyin_i_0_0\ : std_logic;

begin 

    ahbcurr_state(1) <= \ahbcurr_state[1]_net_1\;
    ahbcurr_state(0) <= \ahbcurr_state[0]_net_1\;
    N_271 <= \N_271\;
    ahbsram_req_d1 <= ahbsram_req_d1_net_1;
    CoreAHBLite_0_AHBmslave3_HREADY_i_1 <= 
        \CoreAHBLite_0_AHBmslave3_HREADY_i_1\;
    un8_hreadyin_i_0 <= un8_hreadyin_i_0_net_1;

    \HWRITE_d\ : SLE
      port map(D => N_277, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => HWRITE_d);
    
    un1_hreadyin_i_a3_0 : CFG4
      generic map(INIT => x"2223")

      port map(A => arbRegSMCurrentState(15), B => 
        \CoreAHBLite_0_AHBmslave3_HREADY_i_1\, C => 
        N_157_i_i_o2_0, D => N_157_i_i_o2_0_out, Y => \N_271\);
    
    \count[1]\ : SLE
      port map(D => N_370_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => counte, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \count[1]_net_1\);
    
    \HADDR_d[1]\ : SLE
      port map(D => N_246, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(1));
    
    \HADDR_d[15]\ : SLE
      port map(D => N_241, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(15));
    
    \count[0]\ : SLE
      port map(D => N_400, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => counte, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \count[0]_net_1\);
    
    ahbsram_req_d1_RNI5FGD1 : CFG3
      generic map(INIT => x"08")

      port map(A => \ahbcurr_state[0]_net_1\, B => N_378, C => 
        ahbsram_req_d1_net_1, Y => N_408);
    
    un8_hreadyin_i_0_0 : CFG2
      generic map(INIT => x"D")

      port map(A => N_225, B => un8_hreadyin_i_0_net_1, Y => 
        \un8_hreadyin_i_0_0\);
    
    \HADDR_d[14]\ : SLE
      port map(D => N_242, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(14));
    
    count_n4_i_o3 : CFG3
      generic map(INIT => x"7F")

      port map(A => \count[2]_net_1\, B => \count[1]_net_1\, C
         => \count[0]_net_1\, Y => N_381);
    
    \HSIZE_d[1]\ : SLE
      port map(D => N_235, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_size(1));
    
    \count_RNO[2]\ : CFG3
      generic map(INIT => x"6A")

      port map(A => \count[2]_net_1\, B => \count[1]_net_1\, C
         => \count[0]_net_1\, Y => N_928_i_0);
    
    \ahbcurr_state_RNIOGBG3_0[0]\ : CFG4
      generic map(INIT => x"1311")

      port map(A => \ahbcurr_state[0]_net_1\, B => 
        \ahbcurr_state[1]_net_1\, C => N_378, D => N_391, Y => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \count_RNO[4]\ : CFG3
      generic map(INIT => x"D2")

      port map(A => \count[3]_net_1\, B => N_381, C => 
        \count[4]_net_1\, Y => N_368_i_0);
    
    \ahbcurr_state_ns_1_0_.m6_0_a4_0_0_0\ : CFG3
      generic map(INIT => x"10")

      port map(A => \ahbcurr_state[0]_net_1\, B => 
        \ahbcurr_state[1]_net_1\, C => N_277, Y => m6_0_a4_0_0);
    
    un8_hreadyin_i_1 : CFG4
      generic map(INIT => x"FAF8")

      port map(A => HTRANS_i_a2_0_0, B => N_120, C => 
        \un8_hreadyin_i_0_0\, D => N_157_i_i_o2_0_out, Y => 
        \un8_hreadyin_i_1\);
    
    \ahbcurr_state[0]\ : SLE
      port map(D => \ahbcurr_state_ns[0]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ahbcurr_state[0]_net_1\);
    
    un8_hreadyin_i_a3_7 : CFG3
      generic map(INIT => x"04")

      port map(A => xhdl1222_2, B => hready_m_xhdl343_11, C => 
        xhdl1222_0, Y => N_305);
    
    \ahbsram_req_d1\ : SLE
      port map(D => \CoreAHBLite_0_AHBmslave3_HREADY_i_1\, CLK
         => CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        ahbsram_req_d1_net_1);
    
    \HADDR_d[9]\ : SLE
      port map(D => N_256, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(9));
    
    \count_RNO[3]\ : CFG2
      generic map(INIT => x"9")

      port map(A => N_381, B => \count[3]_net_1\, Y => N_57_i_i_0);
    
    \ahbcurr_state_RNIOGBG3[0]\ : CFG4
      generic map(INIT => x"ECEE")

      port map(A => \ahbcurr_state[0]_net_1\, B => 
        \ahbcurr_state[1]_net_1\, C => N_378, D => N_391, Y => 
        \CoreAHBLite_0_AHBmslave3_HREADY_i_1\);
    
    \count_RNO[1]\ : CFG3
      generic map(INIT => x"48")

      port map(A => \count[0]_net_1\, B => N_391, C => 
        \count[1]_net_1\, Y => N_370_i_0);
    
    \HADDR_d[8]\ : SLE
      port map(D => N_257, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(8));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \count[2]\ : SLE
      port map(D => N_928_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => counte, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \count[2]_net_1\);
    
    \burst_count_reg_RNIJLC51[0]\ : CFG4
      generic map(INIT => x"FFBE")

      port map(A => \count[1]_net_1\, B => \count[0]_net_1\, C
         => \burst_count_reg[0]_net_1\, D => \count[2]_net_1\, Y
         => un1_sramahb_ack_i_i_0_o3_1);
    
    \ahbcurr_state[1]\ : SLE
      port map(D => \ahbcurr_state_ns[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ahbcurr_state[1]_net_1\);
    
    \count_RNIS3IO1[4]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \count[3]_net_1\, B => 
        un1_sramahb_ack_i_i_0_o3_1, C => \count[4]_net_1\, Y => 
        N_391);
    
    ahbsram_req_d1_RNIA0LG3 : CFG4
      generic map(INIT => x"F4FF")

      port map(A => ahbsram_req_d1_net_1, B => 
        \ahbcurr_state[1]_net_1\, C => N_408, D => N_391, Y => 
        counte);
    
    \ahbcurr_state_ns_1_0_.m9_0\ : CFG4
      generic map(INIT => x"8C88")

      port map(A => \ahbcurr_state[1]_net_1\, B => m9_0_1, C => 
        \un8_hreadyin_i_1\, D => \N_271\, Y => 
        \ahbcurr_state_ns[1]\);
    
    \ahbcurr_state_ns_1_0_.m6_0\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => \un8_hreadyin_i_1\, B => \N_271\, C => N_403, 
        D => m6_0_a4_0_0, Y => \ahbcurr_state_ns[0]\);
    
    \ahbcurr_state_ns_1_0_.m9_0_1\ : CFG4
      generic map(INIT => x"2301")

      port map(A => \ahbcurr_state[1]_net_1\, B => 
        \ahbcurr_state[0]_net_1\, C => N_277, D => N_378, Y => 
        m9_0_1);
    
    \HADDR_d[12]\ : SLE
      port map(D => N_244, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(12));
    
    \ahbcurr_state_ns_1_0_.m6_0_a4\ : CFG4
      generic map(INIT => x"2220")

      port map(A => \ahbcurr_state[0]_net_1\, B => 
        \ahbcurr_state[1]_net_1\, C => N_378, D => N_391, Y => 
        N_403);
    
    un8_hreadyin_i_a3_9 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl343_10, B => hready_m_xhdl344_7, 
        Y => N_335);
    
    \HADDR_d[13]\ : SLE
      port map(D => N_243, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(13));
    
    \HADDR_d[3]\ : SLE
      port map(D => N_194_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(3));
    
    count_n0_i_a4 : CFG2
      generic map(INIT => x"2")

      port map(A => N_391, B => \count[0]_net_1\, Y => N_400);
    
    \ahbcurr_state_ns_1_0_.m9_0_o3\ : CFG3
      generic map(INIT => x"37")

      port map(A => sramcurr_state(0), B => sram_done, C => 
        sramcurr_state(1), Y => N_378);
    
    un8_hreadyin_i_o2_1 : CFG4
      generic map(INIT => x"0116")

      port map(A => SDATASELInt_13, B => SDATASELInt_12, C => 
        SDATASELInt_11, D => SDATASELInt_10, Y => N_216);
    
    \HADDR_d[10]\ : SLE
      port map(D => N_255, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(10));
    
    un8_hreadyin_i_o2_0 : CFG4
      generic map(INIT => x"0116")

      port map(A => SDATASELInt_9, B => SDATASELInt_8, C => 
        SDATASELInt_7, D => SDATASELInt_6, Y => N_215);
    
    \count[3]\ : SLE
      port map(D => N_57_i_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => counte, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \count[3]_net_1\);
    
    \HSIZE_d[0]\ : SLE
      port map(D => N_236, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_size(0));
    
    \burst_count_reg[0]\ : SLE
      port map(D => VCC_net_1, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_113_i_0, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \burst_count_reg[0]_net_1\);
    
    \HADDR_d[7]\ : SLE
      port map(D => N_258, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(7));
    
    \HADDR_d[6]\ : SLE
      port map(D => N_259, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(6));
    
    \burst_count_reg_RNO[0]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \CoreAHBLite_0_AHBmslave3_HREADY_i_1\, B => 
        hsel2_i_4, C => \un8_hreadyin_i_1\, Y => N_113_i_0);
    
    \un8_hreadyin_i_0\ : CFG4
      generic map(INIT => x"DC50")

      port map(A => CertificationSystem_sb_0_AHBmslave5_HREADY, B
         => defSlaveSMNextState, C => hready_m_xhdl345, D => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        Y => un8_hreadyin_i_0_net_1);
    
    un8_hreadyin_i_o2 : CFG4
      generic map(INIT => x"0116")

      port map(A => SDATASELInt_4, B => SDATASELInt_2, C => 
        SDATASELInt_1, D => SDATASELInt_0, Y => N_214);
    
    \HADDR_d[2]\ : SLE
      port map(D => N_276, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(2));
    
    \HADDR_d[4]\ : SLE
      port map(D => N_195_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(4));
    
    \HADDR_d[5]\ : SLE
      port map(D => N_196_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(5));
    
    \HADDR_d[0]\ : SLE
      port map(D => N_247, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(0));
    
    \count[4]\ : SLE
      port map(D => N_368_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => counte, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \count[4]_net_1\);
    
    \HADDR_d[11]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave3_HADDR(11), CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => \N_271\, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => ahbsram_addr(11));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM is

    port( CoreAHBLite_0_AHBmslave3_HADDR                          : in    std_logic_vector(11 to 11);
          arbRegSMCurrentState                                    : in    std_logic_vector(15 to 15);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP : in    std_logic_vector(0 to 0);
          CoreAHBLite_0_AHBmslave3_HRDATA                         : out   std_logic_vector(31 downto 0);
          xhdl1222_2                                              : in    std_logic;
          xhdl1222_0                                              : in    std_logic;
          SDATASELInt_9                                           : in    std_logic;
          SDATASELInt_8                                           : in    std_logic;
          SDATASELInt_7                                           : in    std_logic;
          SDATASELInt_6                                           : in    std_logic;
          SDATASELInt_13                                          : in    std_logic;
          SDATASELInt_12                                          : in    std_logic;
          SDATASELInt_11                                          : in    std_logic;
          SDATASELInt_10                                          : in    std_logic;
          SDATASELInt_4                                           : in    std_logic;
          SDATASELInt_2                                           : in    std_logic;
          SDATASELInt_1                                           : in    std_logic;
          SDATASELInt_0                                           : in    std_logic;
          MSS_READY                                               : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                    : in    std_logic;
          N_236                                                   : in    std_logic;
          N_271                                                   : out   std_logic;
          N_235                                                   : in    std_logic;
          N_246                                                   : in    std_logic;
          N_276                                                   : in    std_logic;
          N_194_i_0                                               : in    std_logic;
          N_195_i_0                                               : in    std_logic;
          N_196_i_0                                               : in    std_logic;
          N_259                                                   : in    std_logic;
          N_258                                                   : in    std_logic;
          N_257                                                   : in    std_logic;
          N_256                                                   : in    std_logic;
          N_255                                                   : in    std_logic;
          N_244                                                   : in    std_logic;
          N_243                                                   : in    std_logic;
          N_242                                                   : in    std_logic;
          N_241                                                   : in    std_logic;
          N_247                                                   : in    std_logic;
          N_277                                                   : in    std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                     : out   std_logic;
          hready_m_xhdl343_11                                     : in    std_logic;
          N_305                                                   : out   std_logic;
          hready_m_xhdl343_10                                     : in    std_logic;
          hready_m_xhdl344_7                                      : in    std_logic;
          N_335                                                   : out   std_logic;
          N_215                                                   : out   std_logic;
          N_216                                                   : out   std_logic;
          N_214                                                   : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                 : out   std_logic;
          N_157_i_i_o2_0                                          : in    std_logic;
          N_157_i_i_o2_0_out                                      : in    std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY              : in    std_logic;
          defSlaveSMNextState                                     : in    std_logic;
          hready_m_xhdl345                                        : in    std_logic;
          un8_hreadyin_i_0                                        : out   std_logic;
          N_225                                                   : in    std_logic;
          HTRANS_i_a2_0_0                                         : in    std_logic;
          N_120                                                   : in    std_logic;
          hsel2_i_4                                               : in    std_logic;
          N_38_i_0                                                : in    std_logic;
          N_40_i_0                                                : in    std_logic;
          N_42_i_0                                                : in    std_logic;
          N_44_i_0                                                : in    std_logic;
          N_46_i_0                                                : in    std_logic;
          N_48_i_0                                                : in    std_logic;
          N_50_i_0                                                : in    std_logic;
          N_52_i_0                                                : in    std_logic;
          N_54_i_0                                                : in    std_logic;
          N_56_i_0                                                : in    std_logic;
          N_58_i_0                                                : in    std_logic;
          N_64_i_0                                                : in    std_logic;
          N_66_i_0                                                : in    std_logic;
          N_68_i_0                                                : in    std_logic;
          N_70_i_0                                                : in    std_logic;
          N_72_i_0                                                : in    std_logic;
          N_74_i_0                                                : in    std_logic;
          N_76_i_0                                                : in    std_logic;
          N_78_i_0                                                : in    std_logic;
          N_80_i_0                                                : in    std_logic;
          N_82_i_0                                                : in    std_logic;
          N_84_i_0                                                : in    std_logic;
          N_86_i_0                                                : in    std_logic;
          N_88_i_0                                                : in    std_logic;
          N_90_i_0                                                : in    std_logic;
          N_92_i_0                                                : in    std_logic;
          N_94_i_0                                                : in    std_logic;
          N_96_i_0                                                : in    std_logic;
          N_98_i_0                                                : in    std_logic;
          N_60_i_0                                                : in    std_logic;
          N_62_i_0                                                : in    std_logic;
          N_63_i_0                                                : in    std_logic
        );

end CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM;

architecture DEF_ARCH of 
        CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf
    port( CoreAHBLite_0_AHBmslave3_HRDATA      : out   std_logic_vector(31 downto 0);
          sramcurr_state                       : out   std_logic_vector(1 downto 0);
          ahbsram_size                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          ahbcurr_state                        : in    std_logic_vector(1 downto 0) := (others => 'U');
          ahbsram_addr                         : in    std_logic_vector(15 downto 0) := (others => 'U');
          MSS_READY                            : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0 : in    std_logic := 'U';
          sram_done                            : out   std_logic;
          HWRITE_d                             : in    std_logic := 'U';
          ahbsram_req_d1                       : in    std_logic := 'U';
          N_38_i_0                             : in    std_logic := 'U';
          N_40_i_0                             : in    std_logic := 'U';
          N_42_i_0                             : in    std_logic := 'U';
          N_44_i_0                             : in    std_logic := 'U';
          N_46_i_0                             : in    std_logic := 'U';
          N_48_i_0                             : in    std_logic := 'U';
          N_50_i_0                             : in    std_logic := 'U';
          N_52_i_0                             : in    std_logic := 'U';
          N_54_i_0                             : in    std_logic := 'U';
          N_56_i_0                             : in    std_logic := 'U';
          N_58_i_0                             : in    std_logic := 'U';
          N_64_i_0                             : in    std_logic := 'U';
          N_66_i_0                             : in    std_logic := 'U';
          N_68_i_0                             : in    std_logic := 'U';
          N_70_i_0                             : in    std_logic := 'U';
          N_72_i_0                             : in    std_logic := 'U';
          N_74_i_0                             : in    std_logic := 'U';
          N_76_i_0                             : in    std_logic := 'U';
          N_78_i_0                             : in    std_logic := 'U';
          N_80_i_0                             : in    std_logic := 'U';
          N_82_i_0                             : in    std_logic := 'U';
          N_84_i_0                             : in    std_logic := 'U';
          N_86_i_0                             : in    std_logic := 'U';
          N_88_i_0                             : in    std_logic := 'U';
          N_90_i_0                             : in    std_logic := 'U';
          N_92_i_0                             : in    std_logic := 'U';
          N_94_i_0                             : in    std_logic := 'U';
          N_96_i_0                             : in    std_logic := 'U';
          N_98_i_0                             : in    std_logic := 'U';
          N_60_i_0                             : in    std_logic := 'U';
          N_62_i_0                             : in    std_logic := 'U';
          N_63_i_0                             : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf
    port( ahbsram_size                                            : out   std_logic_vector(1 downto 0);
          CoreAHBLite_0_AHBmslave3_HADDR                          : in    std_logic_vector(11 to 11) := (others => 'U');
          ahbsram_addr                                            : out   std_logic_vector(15 downto 0);
          ahbcurr_state                                           : out   std_logic_vector(1 downto 0);
          sramcurr_state                                          : in    std_logic_vector(1 downto 0) := (others => 'U');
          arbRegSMCurrentState                                    : in    std_logic_vector(15 to 15) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP : in    std_logic_vector(0 to 0) := (others => 'U');
          xhdl1222_2                                              : in    std_logic := 'U';
          xhdl1222_0                                              : in    std_logic := 'U';
          SDATASELInt_9                                           : in    std_logic := 'U';
          SDATASELInt_8                                           : in    std_logic := 'U';
          SDATASELInt_7                                           : in    std_logic := 'U';
          SDATASELInt_6                                           : in    std_logic := 'U';
          SDATASELInt_13                                          : in    std_logic := 'U';
          SDATASELInt_12                                          : in    std_logic := 'U';
          SDATASELInt_11                                          : in    std_logic := 'U';
          SDATASELInt_10                                          : in    std_logic := 'U';
          SDATASELInt_4                                           : in    std_logic := 'U';
          SDATASELInt_2                                           : in    std_logic := 'U';
          SDATASELInt_1                                           : in    std_logic := 'U';
          SDATASELInt_0                                           : in    std_logic := 'U';
          MSS_READY                                               : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                    : in    std_logic := 'U';
          N_236                                                   : in    std_logic := 'U';
          N_271                                                   : out   std_logic;
          N_235                                                   : in    std_logic := 'U';
          N_246                                                   : in    std_logic := 'U';
          N_276                                                   : in    std_logic := 'U';
          N_194_i_0                                               : in    std_logic := 'U';
          N_195_i_0                                               : in    std_logic := 'U';
          N_196_i_0                                               : in    std_logic := 'U';
          N_259                                                   : in    std_logic := 'U';
          N_258                                                   : in    std_logic := 'U';
          N_257                                                   : in    std_logic := 'U';
          N_256                                                   : in    std_logic := 'U';
          N_255                                                   : in    std_logic := 'U';
          N_244                                                   : in    std_logic := 'U';
          N_243                                                   : in    std_logic := 'U';
          N_242                                                   : in    std_logic := 'U';
          N_241                                                   : in    std_logic := 'U';
          N_247                                                   : in    std_logic := 'U';
          HWRITE_d                                                : out   std_logic;
          N_277                                                   : in    std_logic := 'U';
          ahbsram_req_d1                                          : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                     : out   std_logic;
          sram_done                                               : in    std_logic := 'U';
          hready_m_xhdl343_11                                     : in    std_logic := 'U';
          N_305                                                   : out   std_logic;
          hready_m_xhdl343_10                                     : in    std_logic := 'U';
          hready_m_xhdl344_7                                      : in    std_logic := 'U';
          N_335                                                   : out   std_logic;
          N_215                                                   : out   std_logic;
          N_216                                                   : out   std_logic;
          N_214                                                   : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                 : out   std_logic;
          N_157_i_i_o2_0                                          : in    std_logic := 'U';
          N_157_i_i_o2_0_out                                      : in    std_logic := 'U';
          CertificationSystem_sb_0_AHBmslave5_HREADY              : in    std_logic := 'U';
          defSlaveSMNextState                                     : in    std_logic := 'U';
          hready_m_xhdl345                                        : in    std_logic := 'U';
          un8_hreadyin_i_0                                        : out   std_logic;
          N_225                                                   : in    std_logic := 'U';
          HTRANS_i_a2_0_0                                         : in    std_logic := 'U';
          N_120                                                   : in    std_logic := 'U';
          hsel2_i_4                                               : in    std_logic := 'U'
        );
  end component;

    signal \ahbsram_size[0]\, \ahbsram_size[1]\, 
        \ahbsram_addr[0]\, \ahbsram_addr[1]\, \ahbsram_addr[2]\, 
        \ahbsram_addr[3]\, \ahbsram_addr[4]\, \ahbsram_addr[5]\, 
        \ahbsram_addr[6]\, \ahbsram_addr[7]\, \ahbsram_addr[8]\, 
        \ahbsram_addr[9]\, \ahbsram_addr[10]\, \ahbsram_addr[11]\, 
        \ahbsram_addr[12]\, \ahbsram_addr[13]\, 
        \ahbsram_addr[14]\, \ahbsram_addr[15]\, 
        \ahbcurr_state[0]\, \ahbcurr_state[1]\, 
        \sramcurr_state[0]\, \sramcurr_state[1]\, HWRITE_d, 
        ahbsram_req_d1, sram_done, GND_net_1, VCC_net_1
         : std_logic;

    for all : CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf
	Use entity work.
        CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf(DEF_ARCH);
    for all : CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf
	Use entity work.
        CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    U_SramCtrlIf : 
        CertificationSystem_sb_COREAHBLSRAM_0_0_SramCtrlIf
      port map(CoreAHBLite_0_AHBmslave3_HRDATA(31) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(31), 
        CoreAHBLite_0_AHBmslave3_HRDATA(30) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(30), 
        CoreAHBLite_0_AHBmslave3_HRDATA(29) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(29), 
        CoreAHBLite_0_AHBmslave3_HRDATA(28) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(28), 
        CoreAHBLite_0_AHBmslave3_HRDATA(27) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(27), 
        CoreAHBLite_0_AHBmslave3_HRDATA(26) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(26), 
        CoreAHBLite_0_AHBmslave3_HRDATA(25) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(25), 
        CoreAHBLite_0_AHBmslave3_HRDATA(24) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(24), 
        CoreAHBLite_0_AHBmslave3_HRDATA(23) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(23), 
        CoreAHBLite_0_AHBmslave3_HRDATA(22) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(22), 
        CoreAHBLite_0_AHBmslave3_HRDATA(21) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(21), 
        CoreAHBLite_0_AHBmslave3_HRDATA(20) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(20), 
        CoreAHBLite_0_AHBmslave3_HRDATA(19) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(19), 
        CoreAHBLite_0_AHBmslave3_HRDATA(18) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(18), 
        CoreAHBLite_0_AHBmslave3_HRDATA(17) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(17), 
        CoreAHBLite_0_AHBmslave3_HRDATA(16) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(16), 
        CoreAHBLite_0_AHBmslave3_HRDATA(15) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(15), 
        CoreAHBLite_0_AHBmslave3_HRDATA(14) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(14), 
        CoreAHBLite_0_AHBmslave3_HRDATA(13) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(13), 
        CoreAHBLite_0_AHBmslave3_HRDATA(12) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(12), 
        CoreAHBLite_0_AHBmslave3_HRDATA(11) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(11), 
        CoreAHBLite_0_AHBmslave3_HRDATA(10) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(10), 
        CoreAHBLite_0_AHBmslave3_HRDATA(9) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(9), 
        CoreAHBLite_0_AHBmslave3_HRDATA(8) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(8), 
        CoreAHBLite_0_AHBmslave3_HRDATA(7) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(7), 
        CoreAHBLite_0_AHBmslave3_HRDATA(6) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(6), 
        CoreAHBLite_0_AHBmslave3_HRDATA(5) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(5), 
        CoreAHBLite_0_AHBmslave3_HRDATA(4) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(4), 
        CoreAHBLite_0_AHBmslave3_HRDATA(3) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(3), 
        CoreAHBLite_0_AHBmslave3_HRDATA(2) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(2), 
        CoreAHBLite_0_AHBmslave3_HRDATA(1) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(1), 
        CoreAHBLite_0_AHBmslave3_HRDATA(0) => 
        CoreAHBLite_0_AHBmslave3_HRDATA(0), sramcurr_state(1) => 
        \sramcurr_state[1]\, sramcurr_state(0) => 
        \sramcurr_state[0]\, ahbsram_size(1) => \ahbsram_size[1]\, 
        ahbsram_size(0) => \ahbsram_size[0]\, ahbcurr_state(1)
         => \ahbcurr_state[1]\, ahbcurr_state(0) => 
        \ahbcurr_state[0]\, ahbsram_addr(15) => 
        \ahbsram_addr[15]\, ahbsram_addr(14) => 
        \ahbsram_addr[14]\, ahbsram_addr(13) => 
        \ahbsram_addr[13]\, ahbsram_addr(12) => 
        \ahbsram_addr[12]\, ahbsram_addr(11) => 
        \ahbsram_addr[11]\, ahbsram_addr(10) => 
        \ahbsram_addr[10]\, ahbsram_addr(9) => \ahbsram_addr[9]\, 
        ahbsram_addr(8) => \ahbsram_addr[8]\, ahbsram_addr(7) => 
        \ahbsram_addr[7]\, ahbsram_addr(6) => \ahbsram_addr[6]\, 
        ahbsram_addr(5) => \ahbsram_addr[5]\, ahbsram_addr(4) => 
        \ahbsram_addr[4]\, ahbsram_addr(3) => \ahbsram_addr[3]\, 
        ahbsram_addr(2) => \ahbsram_addr[2]\, ahbsram_addr(1) => 
        \ahbsram_addr[1]\, ahbsram_addr(0) => \ahbsram_addr[0]\, 
        MSS_READY => MSS_READY, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, sram_done => 
        sram_done, HWRITE_d => HWRITE_d, ahbsram_req_d1 => 
        ahbsram_req_d1, N_38_i_0 => N_38_i_0, N_40_i_0 => 
        N_40_i_0, N_42_i_0 => N_42_i_0, N_44_i_0 => N_44_i_0, 
        N_46_i_0 => N_46_i_0, N_48_i_0 => N_48_i_0, N_50_i_0 => 
        N_50_i_0, N_52_i_0 => N_52_i_0, N_54_i_0 => N_54_i_0, 
        N_56_i_0 => N_56_i_0, N_58_i_0 => N_58_i_0, N_64_i_0 => 
        N_64_i_0, N_66_i_0 => N_66_i_0, N_68_i_0 => N_68_i_0, 
        N_70_i_0 => N_70_i_0, N_72_i_0 => N_72_i_0, N_74_i_0 => 
        N_74_i_0, N_76_i_0 => N_76_i_0, N_78_i_0 => N_78_i_0, 
        N_80_i_0 => N_80_i_0, N_82_i_0 => N_82_i_0, N_84_i_0 => 
        N_84_i_0, N_86_i_0 => N_86_i_0, N_88_i_0 => N_88_i_0, 
        N_90_i_0 => N_90_i_0, N_92_i_0 => N_92_i_0, N_94_i_0 => 
        N_94_i_0, N_96_i_0 => N_96_i_0, N_98_i_0 => N_98_i_0, 
        N_60_i_0 => N_60_i_0, N_62_i_0 => N_62_i_0, N_63_i_0 => 
        N_63_i_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    U_CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf : 
        CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf
      port map(ahbsram_size(1) => \ahbsram_size[1]\, 
        ahbsram_size(0) => \ahbsram_size[0]\, 
        CoreAHBLite_0_AHBmslave3_HADDR(11) => 
        CoreAHBLite_0_AHBmslave3_HADDR(11), ahbsram_addr(15) => 
        \ahbsram_addr[15]\, ahbsram_addr(14) => 
        \ahbsram_addr[14]\, ahbsram_addr(13) => 
        \ahbsram_addr[13]\, ahbsram_addr(12) => 
        \ahbsram_addr[12]\, ahbsram_addr(11) => 
        \ahbsram_addr[11]\, ahbsram_addr(10) => 
        \ahbsram_addr[10]\, ahbsram_addr(9) => \ahbsram_addr[9]\, 
        ahbsram_addr(8) => \ahbsram_addr[8]\, ahbsram_addr(7) => 
        \ahbsram_addr[7]\, ahbsram_addr(6) => \ahbsram_addr[6]\, 
        ahbsram_addr(5) => \ahbsram_addr[5]\, ahbsram_addr(4) => 
        \ahbsram_addr[4]\, ahbsram_addr(3) => \ahbsram_addr[3]\, 
        ahbsram_addr(2) => \ahbsram_addr[2]\, ahbsram_addr(1) => 
        \ahbsram_addr[1]\, ahbsram_addr(0) => \ahbsram_addr[0]\, 
        ahbcurr_state(1) => \ahbcurr_state[1]\, ahbcurr_state(0)
         => \ahbcurr_state[0]\, sramcurr_state(1) => 
        \sramcurr_state[1]\, sramcurr_state(0) => 
        \sramcurr_state[0]\, arbRegSMCurrentState(15) => 
        arbRegSMCurrentState(15), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0), 
        xhdl1222_2 => xhdl1222_2, xhdl1222_0 => xhdl1222_0, 
        SDATASELInt_9 => SDATASELInt_9, SDATASELInt_8 => 
        SDATASELInt_8, SDATASELInt_7 => SDATASELInt_7, 
        SDATASELInt_6 => SDATASELInt_6, SDATASELInt_13 => 
        SDATASELInt_13, SDATASELInt_12 => SDATASELInt_12, 
        SDATASELInt_11 => SDATASELInt_11, SDATASELInt_10 => 
        SDATASELInt_10, SDATASELInt_4 => SDATASELInt_4, 
        SDATASELInt_2 => SDATASELInt_2, SDATASELInt_1 => 
        SDATASELInt_1, SDATASELInt_0 => SDATASELInt_0, MSS_READY
         => MSS_READY, CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, N_236 => N_236, 
        N_271 => N_271, N_235 => N_235, N_246 => N_246, N_276 => 
        N_276, N_194_i_0 => N_194_i_0, N_195_i_0 => N_195_i_0, 
        N_196_i_0 => N_196_i_0, N_259 => N_259, N_258 => N_258, 
        N_257 => N_257, N_256 => N_256, N_255 => N_255, N_244 => 
        N_244, N_243 => N_243, N_242 => N_242, N_241 => N_241, 
        N_247 => N_247, HWRITE_d => HWRITE_d, N_277 => N_277, 
        ahbsram_req_d1 => ahbsram_req_d1, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, sram_done => 
        sram_done, hready_m_xhdl343_11 => hready_m_xhdl343_11, 
        N_305 => N_305, hready_m_xhdl343_10 => 
        hready_m_xhdl343_10, hready_m_xhdl344_7 => 
        hready_m_xhdl344_7, N_335 => N_335, N_215 => N_215, N_216
         => N_216, N_214 => N_214, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, N_157_i_i_o2_0
         => N_157_i_i_o2_0, N_157_i_i_o2_0_out => 
        N_157_i_i_o2_0_out, 
        CertificationSystem_sb_0_AHBmslave5_HREADY => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, 
        defSlaveSMNextState => defSlaveSMNextState, 
        hready_m_xhdl345 => hready_m_xhdl345, un8_hreadyin_i_0
         => un8_hreadyin_i_0, N_225 => N_225, HTRANS_i_a2_0_0 => 
        HTRANS_i_a2_0_0, N_120 => N_120, hsel2_i_4 => hsel2_i_4);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem_sb is

    port( result_addr_net_0                          : in    std_logic_vector(3 downto 0);
          line_7                                     : in    std_logic_vector(2 downto 1);
          xhdl1222_2                                 : out   std_logic;
          line_13                                    : in    std_logic;
          line_10                                    : in    std_logic;
          line_21                                    : in    std_logic;
          line_24                                    : in    std_logic;
          line_18                                    : in    std_logic;
          line_23                                    : in    std_logic;
          line_16                                    : in    std_logic;
          line_28                                    : in    std_logic;
          line_9                                     : in    std_logic;
          line_3_d0                                  : in    std_logic;
          line_5_d0                                  : in    std_logic;
          line_15                                    : in    std_logic;
          line_26                                    : in    std_logic;
          line_14                                    : in    std_logic;
          line_20                                    : in    std_logic;
          line_2_d0                                  : in    std_logic;
          line_25                                    : in    std_logic;
          line_29                                    : in    std_logic;
          line_19                                    : in    std_logic;
          line_27                                    : in    std_logic;
          line_30                                    : in    std_logic;
          line_17                                    : in    std_logic;
          line_8                                     : in    std_logic;
          line_0_d0                                  : in    std_logic;
          line_6_d0                                  : in    std_logic;
          line_1_d0                                  : in    std_logic;
          line_0_10                                  : in    std_logic;
          line_0_21                                  : in    std_logic;
          line_0_24                                  : in    std_logic;
          line_0_18                                  : in    std_logic;
          line_0_23                                  : in    std_logic;
          line_0_16                                  : in    std_logic;
          line_0_28                                  : in    std_logic;
          line_0_9                                   : in    std_logic;
          line_0_3                                   : in    std_logic;
          line_0_5                                   : in    std_logic;
          line_0_15                                  : in    std_logic;
          line_0_26                                  : in    std_logic;
          line_0_14                                  : in    std_logic;
          line_0_20                                  : in    std_logic;
          line_0_2                                   : in    std_logic;
          line_0_25                                  : in    std_logic;
          line_0_29                                  : in    std_logic;
          line_0_19                                  : in    std_logic;
          line_0_27                                  : in    std_logic;
          line_0_30                                  : in    std_logic;
          line_0_17                                  : in    std_logic;
          line_0_8                                   : in    std_logic;
          line_0_0                                   : in    std_logic;
          line_0_1                                   : in    std_logic;
          line_0_6                                   : in    std_logic;
          line_0_13                                  : in    std_logic;
          line_1_10                                  : in    std_logic;
          line_1_21                                  : in    std_logic;
          line_1_24                                  : in    std_logic;
          line_1_18                                  : in    std_logic;
          line_1_23                                  : in    std_logic;
          line_1_16                                  : in    std_logic;
          line_1_28                                  : in    std_logic;
          line_1_9                                   : in    std_logic;
          line_1_3                                   : in    std_logic;
          line_1_5                                   : in    std_logic;
          line_1_15                                  : in    std_logic;
          line_1_26                                  : in    std_logic;
          line_1_14                                  : in    std_logic;
          line_1_20                                  : in    std_logic;
          line_1_2                                   : in    std_logic;
          line_1_25                                  : in    std_logic;
          line_1_29                                  : in    std_logic;
          line_1_19                                  : in    std_logic;
          line_1_27                                  : in    std_logic;
          line_1_30                                  : in    std_logic;
          line_1_17                                  : in    std_logic;
          line_1_8                                   : in    std_logic;
          line_1_0                                   : in    std_logic;
          line_1_1                                   : in    std_logic;
          line_1_6                                   : in    std_logic;
          line_1_13                                  : in    std_logic;
          line_2_19                                  : in    std_logic;
          line_2_27                                  : in    std_logic;
          line_2_30                                  : in    std_logic;
          line_2_17                                  : in    std_logic;
          line_2_8                                   : in    std_logic;
          line_2_10                                  : in    std_logic;
          line_2_15                                  : in    std_logic;
          line_2_26                                  : in    std_logic;
          line_2_20                                  : in    std_logic;
          line_2_0                                   : in    std_logic;
          line_2_1                                   : in    std_logic;
          line_2_29                                  : in    std_logic;
          line_2_25                                  : in    std_logic;
          line_2_2                                   : in    std_logic;
          line_2_6                                   : in    std_logic;
          line_2_13                                  : in    std_logic;
          line_2_14                                  : in    std_logic;
          line_2_5                                   : in    std_logic;
          line_2_3                                   : in    std_logic;
          line_2_9                                   : in    std_logic;
          line_2_28                                  : in    std_logic;
          line_2_16                                  : in    std_logic;
          line_2_23                                  : in    std_logic;
          line_2_18                                  : in    std_logic;
          line_2_24                                  : in    std_logic;
          line_2_21                                  : in    std_logic;
          line_3_19                                  : in    std_logic;
          line_3_17                                  : in    std_logic;
          line_3_8                                   : in    std_logic;
          line_3_0                                   : in    std_logic;
          line_3_1                                   : in    std_logic;
          line_3_29                                  : in    std_logic;
          line_3_25                                  : in    std_logic;
          line_3_2                                   : in    std_logic;
          line_3_20                                  : in    std_logic;
          line_3_6                                   : in    std_logic;
          line_3_13                                  : in    std_logic;
          line_3_14                                  : in    std_logic;
          line_3_26                                  : in    std_logic;
          line_3_15                                  : in    std_logic;
          line_3_5                                   : in    std_logic;
          line_3_3                                   : in    std_logic;
          line_3_9                                   : in    std_logic;
          line_3_28                                  : in    std_logic;
          line_3_16                                  : in    std_logic;
          line_3_23                                  : in    std_logic;
          line_3_18                                  : in    std_logic;
          line_3_24                                  : in    std_logic;
          line_3_21                                  : in    std_logic;
          line_3_10                                  : in    std_logic;
          SHA256_Module_0_data_out_5                 : in    std_logic;
          SHA256_Module_0_data_out_13                : in    std_logic;
          SHA256_Module_0_data_out_12                : in    std_logic;
          SHA256_Module_0_data_out_8                 : in    std_logic;
          SHA256_Module_0_data_out_23                : in    std_logic;
          SHA256_Module_0_data_out_0                 : in    std_logic;
          line_4_19                                  : in    std_logic;
          line_4_17                                  : in    std_logic;
          line_4_8                                   : in    std_logic;
          line_4_0                                   : in    std_logic;
          line_4_1                                   : in    std_logic;
          line_4_29                                  : in    std_logic;
          line_4_25                                  : in    std_logic;
          line_4_2                                   : in    std_logic;
          line_4_20                                  : in    std_logic;
          line_4_14                                  : in    std_logic;
          line_4_26                                  : in    std_logic;
          line_4_15                                  : in    std_logic;
          line_4_5                                   : in    std_logic;
          line_4_3                                   : in    std_logic;
          line_4_9                                   : in    std_logic;
          line_4_28                                  : in    std_logic;
          line_4_16                                  : in    std_logic;
          line_4_23                                  : in    std_logic;
          line_4_18                                  : in    std_logic;
          line_4_24                                  : in    std_logic;
          line_4_21                                  : in    std_logic;
          line_4_10                                  : in    std_logic;
          line_4_6                                   : in    std_logic;
          line_4_13                                  : in    std_logic;
          line_5_19                                  : in    std_logic;
          line_5_17                                  : in    std_logic;
          line_5_8                                   : in    std_logic;
          line_5_0                                   : in    std_logic;
          line_5_1                                   : in    std_logic;
          line_5_29                                  : in    std_logic;
          line_5_25                                  : in    std_logic;
          line_5_2                                   : in    std_logic;
          line_5_20                                  : in    std_logic;
          line_5_6                                   : in    std_logic;
          line_5_13                                  : in    std_logic;
          line_5_14                                  : in    std_logic;
          line_5_26                                  : in    std_logic;
          line_5_15                                  : in    std_logic;
          line_5_5                                   : in    std_logic;
          line_5_3                                   : in    std_logic;
          line_5_9                                   : in    std_logic;
          line_5_28                                  : in    std_logic;
          line_5_16                                  : in    std_logic;
          line_5_23                                  : in    std_logic;
          line_5_18                                  : in    std_logic;
          line_5_24                                  : in    std_logic;
          line_5_21                                  : in    std_logic;
          line_5_10                                  : in    std_logic;
          line_6_19                                  : in    std_logic;
          line_6_17                                  : in    std_logic;
          line_6_8                                   : in    std_logic;
          line_6_0                                   : in    std_logic;
          line_6_1                                   : in    std_logic;
          line_6_29                                  : in    std_logic;
          line_6_25                                  : in    std_logic;
          line_6_2                                   : in    std_logic;
          line_6_20                                  : in    std_logic;
          line_6_6                                   : in    std_logic;
          line_6_13                                  : in    std_logic;
          line_6_14                                  : in    std_logic;
          line_6_26                                  : in    std_logic;
          line_6_15                                  : in    std_logic;
          line_6_5                                   : in    std_logic;
          line_6_3                                   : in    std_logic;
          line_6_9                                   : in    std_logic;
          line_6_28                                  : in    std_logic;
          line_6_16                                  : in    std_logic;
          line_6_23                                  : in    std_logic;
          line_6_18                                  : in    std_logic;
          line_6_24                                  : in    std_logic;
          line_6_21                                  : in    std_logic;
          line_6_10                                  : in    std_logic;
          CertificationSystem_sb_0_POWER_ON_RESET_N  : out   std_logic;
          DEVRST_N                                   : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0       : out   std_logic;
          SPI_0_SS0                                  : inout std_logic := 'Z';
          SPI_0_DO                                   : out   std_logic;
          SPI_0_DI                                   : in    std_logic;
          SPI_0_CLK                                  : inout std_logic := 'Z';
          MMUART_1_TXD                               : out   std_logic;
          MMUART_1_RXD                               : in    std_logic;
          CertificationSystem_sb_0_GPIO_1_M2F        : out   std_logic;
          GPIO_0_M2F_c                               : out   std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F        : out   std_logic;
          SHA256_Module_0_waiting_data               : in    std_logic;
          SHA256_Module_0_data_available_lastbank_8  : in    std_logic;
          SHA256_Module_0_di_req_o                   : in    std_logic;
          SHA256_Module_0_do_valid_o                 : in    std_logic;
          SHA256_Module_0_data_available             : in    std_logic;
          SHA256_Module_0_error_o                    : in    std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY : in    std_logic;
          N_225                                      : out   std_logic;
          N_276                                      : out   std_logic;
          N_259                                      : out   std_logic;
          N_277                                      : out   std_logic;
          ren_pos                                    : in    std_logic;
          N_206                                      : out   std_logic;
          N_508                                      : in    std_logic;
          N_507                                      : in    std_logic;
          un8_hreadyin_i_0                           : out   std_logic;
          N_226                                      : out   std_logic;
          N_65_i_0                                   : out   std_logic;
          N_67_i_0                                   : out   std_logic;
          N_110_i_0                                  : out   std_logic;
          N_112_i_0                                  : out   std_logic;
          N_114_i_0                                  : out   std_logic;
          N_116_i_0                                  : out   std_logic;
          N_69_i_0                                   : out   std_logic;
          N_71_i_0                                   : out   std_logic;
          N_73_i_0                                   : out   std_logic;
          N_75_i_0                                   : out   std_logic;
          N_77_i_0                                   : out   std_logic;
          N_83_i_0                                   : out   std_logic;
          N_85_i_0                                   : out   std_logic;
          N_133_i_0                                  : out   std_logic;
          N_87_i_0                                   : out   std_logic;
          N_89_i_0                                   : out   std_logic;
          N_140_i_0                                  : out   std_logic;
          N_91_i_0                                   : out   std_logic;
          N_93_i_0                                   : out   std_logic;
          N_95_i_0                                   : out   std_logic;
          N_97_i_0                                   : out   std_logic;
          N_99_i_0                                   : out   std_logic;
          N_152_i_0                                  : out   std_logic;
          N_101_i_0                                  : out   std_logic;
          N_156_i_0                                  : out   std_logic;
          N_158_i_0                                  : out   std_logic;
          N_103_i_0                                  : out   std_logic;
          N_105_i_0                                  : out   std_logic;
          N_107_i_0                                  : out   std_logic;
          N_168_i_0                                  : out   std_logic;
          N_109_i_0                                  : out   std_logic;
          N_111_i_0                                  : out   std_logic;
          N_218_i_0                                  : out   std_logic;
          N_217_i_0                                  : out   std_logic;
          N_203_i_0                                  : out   std_logic
        );

end CertificationSystem_sb;

architecture DEF_ARCH of CertificationSystem_sb is 

  component CertificationSystem_sb_FABOSC_0_OSC
    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );
  end component;

  component CoreResetP
    port( MSS_READY                                             : out   std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0                  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic := 'U';
          CertificationSystem_sb_0_POWER_ON_RESET_N             : in    std_logic := 'U'
        );
  end component;

  component CoreAHBLite
    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE     : in    std_logic_vector(1 downto 0) := (others => 'U');
          arbRegSMCurrentState                                        : out   std_logic_vector(15 to 15);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS    : in    std_logic_vector(1 to 1) := (others => 'U');
          result_addr_net_0                                           : in    std_logic_vector(3 downto 0) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP     : out   std_logic_vector(0 to 0);
          CoreAHBLite_0_AHBmslave3_HRDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          line_7                                                      : in    std_logic_vector(2 downto 1) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA    : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HADDR                              : out   std_logic_vector(11 to 11);
          xhdl1222_0                                                  : out   std_logic;
          xhdl1222_2                                                  : out   std_logic;
          SDATASELInt_0                                               : out   std_logic;
          SDATASELInt_1                                               : out   std_logic;
          SDATASELInt_2                                               : out   std_logic;
          SDATASELInt_4                                               : out   std_logic;
          SDATASELInt_6                                               : out   std_logic;
          SDATASELInt_7                                               : out   std_logic;
          SDATASELInt_8                                               : out   std_logic;
          SDATASELInt_9                                               : out   std_logic;
          SDATASELInt_10                                              : out   std_logic;
          SDATASELInt_11                                              : out   std_logic;
          SDATASELInt_12                                              : out   std_logic;
          SDATASELInt_13                                              : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31  : in    std_logic := 'U';
          line_13                                                     : in    std_logic := 'U';
          line_10                                                     : in    std_logic := 'U';
          line_21                                                     : in    std_logic := 'U';
          line_24                                                     : in    std_logic := 'U';
          line_18                                                     : in    std_logic := 'U';
          line_23                                                     : in    std_logic := 'U';
          line_16                                                     : in    std_logic := 'U';
          line_28                                                     : in    std_logic := 'U';
          line_9                                                      : in    std_logic := 'U';
          line_3_d0                                                   : in    std_logic := 'U';
          line_5_d0                                                   : in    std_logic := 'U';
          line_15                                                     : in    std_logic := 'U';
          line_26                                                     : in    std_logic := 'U';
          line_14                                                     : in    std_logic := 'U';
          line_20                                                     : in    std_logic := 'U';
          line_2_d0                                                   : in    std_logic := 'U';
          line_25                                                     : in    std_logic := 'U';
          line_29                                                     : in    std_logic := 'U';
          line_19                                                     : in    std_logic := 'U';
          line_27                                                     : in    std_logic := 'U';
          line_30                                                     : in    std_logic := 'U';
          line_17                                                     : in    std_logic := 'U';
          line_8                                                      : in    std_logic := 'U';
          line_0_d0                                                   : in    std_logic := 'U';
          line_6_d0                                                   : in    std_logic := 'U';
          line_1_d0                                                   : in    std_logic := 'U';
          line_0_10                                                   : in    std_logic := 'U';
          line_0_21                                                   : in    std_logic := 'U';
          line_0_24                                                   : in    std_logic := 'U';
          line_0_18                                                   : in    std_logic := 'U';
          line_0_23                                                   : in    std_logic := 'U';
          line_0_16                                                   : in    std_logic := 'U';
          line_0_28                                                   : in    std_logic := 'U';
          line_0_9                                                    : in    std_logic := 'U';
          line_0_3                                                    : in    std_logic := 'U';
          line_0_5                                                    : in    std_logic := 'U';
          line_0_15                                                   : in    std_logic := 'U';
          line_0_26                                                   : in    std_logic := 'U';
          line_0_14                                                   : in    std_logic := 'U';
          line_0_20                                                   : in    std_logic := 'U';
          line_0_2                                                    : in    std_logic := 'U';
          line_0_25                                                   : in    std_logic := 'U';
          line_0_29                                                   : in    std_logic := 'U';
          line_0_19                                                   : in    std_logic := 'U';
          line_0_27                                                   : in    std_logic := 'U';
          line_0_30                                                   : in    std_logic := 'U';
          line_0_17                                                   : in    std_logic := 'U';
          line_0_8                                                    : in    std_logic := 'U';
          line_0_0                                                    : in    std_logic := 'U';
          line_0_1                                                    : in    std_logic := 'U';
          line_0_6                                                    : in    std_logic := 'U';
          line_0_13                                                   : in    std_logic := 'U';
          line_1_10                                                   : in    std_logic := 'U';
          line_1_21                                                   : in    std_logic := 'U';
          line_1_24                                                   : in    std_logic := 'U';
          line_1_18                                                   : in    std_logic := 'U';
          line_1_23                                                   : in    std_logic := 'U';
          line_1_16                                                   : in    std_logic := 'U';
          line_1_28                                                   : in    std_logic := 'U';
          line_1_9                                                    : in    std_logic := 'U';
          line_1_3                                                    : in    std_logic := 'U';
          line_1_5                                                    : in    std_logic := 'U';
          line_1_15                                                   : in    std_logic := 'U';
          line_1_26                                                   : in    std_logic := 'U';
          line_1_14                                                   : in    std_logic := 'U';
          line_1_20                                                   : in    std_logic := 'U';
          line_1_2                                                    : in    std_logic := 'U';
          line_1_25                                                   : in    std_logic := 'U';
          line_1_29                                                   : in    std_logic := 'U';
          line_1_19                                                   : in    std_logic := 'U';
          line_1_27                                                   : in    std_logic := 'U';
          line_1_30                                                   : in    std_logic := 'U';
          line_1_17                                                   : in    std_logic := 'U';
          line_1_8                                                    : in    std_logic := 'U';
          line_1_0                                                    : in    std_logic := 'U';
          line_1_1                                                    : in    std_logic := 'U';
          line_1_6                                                    : in    std_logic := 'U';
          line_1_13                                                   : in    std_logic := 'U';
          line_2_19                                                   : in    std_logic := 'U';
          line_2_27                                                   : in    std_logic := 'U';
          line_2_30                                                   : in    std_logic := 'U';
          line_2_17                                                   : in    std_logic := 'U';
          line_2_8                                                    : in    std_logic := 'U';
          line_2_10                                                   : in    std_logic := 'U';
          line_2_15                                                   : in    std_logic := 'U';
          line_2_26                                                   : in    std_logic := 'U';
          line_2_20                                                   : in    std_logic := 'U';
          line_2_0                                                    : in    std_logic := 'U';
          line_2_1                                                    : in    std_logic := 'U';
          line_2_29                                                   : in    std_logic := 'U';
          line_2_25                                                   : in    std_logic := 'U';
          line_2_2                                                    : in    std_logic := 'U';
          line_2_6                                                    : in    std_logic := 'U';
          line_2_13                                                   : in    std_logic := 'U';
          line_2_14                                                   : in    std_logic := 'U';
          line_2_5                                                    : in    std_logic := 'U';
          line_2_3                                                    : in    std_logic := 'U';
          line_2_9                                                    : in    std_logic := 'U';
          line_2_28                                                   : in    std_logic := 'U';
          line_2_16                                                   : in    std_logic := 'U';
          line_2_23                                                   : in    std_logic := 'U';
          line_2_18                                                   : in    std_logic := 'U';
          line_2_24                                                   : in    std_logic := 'U';
          line_2_21                                                   : in    std_logic := 'U';
          line_3_19                                                   : in    std_logic := 'U';
          line_3_17                                                   : in    std_logic := 'U';
          line_3_8                                                    : in    std_logic := 'U';
          line_3_0                                                    : in    std_logic := 'U';
          line_3_1                                                    : in    std_logic := 'U';
          line_3_29                                                   : in    std_logic := 'U';
          line_3_25                                                   : in    std_logic := 'U';
          line_3_2                                                    : in    std_logic := 'U';
          line_3_20                                                   : in    std_logic := 'U';
          line_3_6                                                    : in    std_logic := 'U';
          line_3_13                                                   : in    std_logic := 'U';
          line_3_14                                                   : in    std_logic := 'U';
          line_3_26                                                   : in    std_logic := 'U';
          line_3_15                                                   : in    std_logic := 'U';
          line_3_5                                                    : in    std_logic := 'U';
          line_3_3                                                    : in    std_logic := 'U';
          line_3_9                                                    : in    std_logic := 'U';
          line_3_28                                                   : in    std_logic := 'U';
          line_3_16                                                   : in    std_logic := 'U';
          line_3_23                                                   : in    std_logic := 'U';
          line_3_18                                                   : in    std_logic := 'U';
          line_3_24                                                   : in    std_logic := 'U';
          line_3_21                                                   : in    std_logic := 'U';
          line_3_10                                                   : in    std_logic := 'U';
          SHA256_Module_0_data_out_5                                  : in    std_logic := 'U';
          SHA256_Module_0_data_out_13                                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_12                                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_8                                  : in    std_logic := 'U';
          SHA256_Module_0_data_out_23                                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_0                                  : in    std_logic := 'U';
          line_4_19                                                   : in    std_logic := 'U';
          line_4_17                                                   : in    std_logic := 'U';
          line_4_8                                                    : in    std_logic := 'U';
          line_4_0                                                    : in    std_logic := 'U';
          line_4_1                                                    : in    std_logic := 'U';
          line_4_29                                                   : in    std_logic := 'U';
          line_4_25                                                   : in    std_logic := 'U';
          line_4_2                                                    : in    std_logic := 'U';
          line_4_20                                                   : in    std_logic := 'U';
          line_4_14                                                   : in    std_logic := 'U';
          line_4_26                                                   : in    std_logic := 'U';
          line_4_15                                                   : in    std_logic := 'U';
          line_4_5                                                    : in    std_logic := 'U';
          line_4_3                                                    : in    std_logic := 'U';
          line_4_9                                                    : in    std_logic := 'U';
          line_4_28                                                   : in    std_logic := 'U';
          line_4_16                                                   : in    std_logic := 'U';
          line_4_23                                                   : in    std_logic := 'U';
          line_4_18                                                   : in    std_logic := 'U';
          line_4_24                                                   : in    std_logic := 'U';
          line_4_21                                                   : in    std_logic := 'U';
          line_4_10                                                   : in    std_logic := 'U';
          line_4_6                                                    : in    std_logic := 'U';
          line_4_13                                                   : in    std_logic := 'U';
          line_5_19                                                   : in    std_logic := 'U';
          line_5_17                                                   : in    std_logic := 'U';
          line_5_8                                                    : in    std_logic := 'U';
          line_5_0                                                    : in    std_logic := 'U';
          line_5_1                                                    : in    std_logic := 'U';
          line_5_29                                                   : in    std_logic := 'U';
          line_5_25                                                   : in    std_logic := 'U';
          line_5_2                                                    : in    std_logic := 'U';
          line_5_20                                                   : in    std_logic := 'U';
          line_5_6                                                    : in    std_logic := 'U';
          line_5_13                                                   : in    std_logic := 'U';
          line_5_14                                                   : in    std_logic := 'U';
          line_5_26                                                   : in    std_logic := 'U';
          line_5_15                                                   : in    std_logic := 'U';
          line_5_5                                                    : in    std_logic := 'U';
          line_5_3                                                    : in    std_logic := 'U';
          line_5_9                                                    : in    std_logic := 'U';
          line_5_28                                                   : in    std_logic := 'U';
          line_5_16                                                   : in    std_logic := 'U';
          line_5_23                                                   : in    std_logic := 'U';
          line_5_18                                                   : in    std_logic := 'U';
          line_5_24                                                   : in    std_logic := 'U';
          line_5_21                                                   : in    std_logic := 'U';
          line_5_10                                                   : in    std_logic := 'U';
          line_6_19                                                   : in    std_logic := 'U';
          line_6_17                                                   : in    std_logic := 'U';
          line_6_8                                                    : in    std_logic := 'U';
          line_6_0                                                    : in    std_logic := 'U';
          line_6_1                                                    : in    std_logic := 'U';
          line_6_29                                                   : in    std_logic := 'U';
          line_6_25                                                   : in    std_logic := 'U';
          line_6_2                                                    : in    std_logic := 'U';
          line_6_20                                                   : in    std_logic := 'U';
          line_6_6                                                    : in    std_logic := 'U';
          line_6_13                                                   : in    std_logic := 'U';
          line_6_14                                                   : in    std_logic := 'U';
          line_6_26                                                   : in    std_logic := 'U';
          line_6_15                                                   : in    std_logic := 'U';
          line_6_5                                                    : in    std_logic := 'U';
          line_6_3                                                    : in    std_logic := 'U';
          line_6_9                                                    : in    std_logic := 'U';
          line_6_28                                                   : in    std_logic := 'U';
          line_6_16                                                   : in    std_logic := 'U';
          line_6_23                                                   : in    std_logic := 'U';
          line_6_18                                                   : in    std_logic := 'U';
          line_6_24                                                   : in    std_logic := 'U';
          line_6_21                                                   : in    std_logic := 'U';
          line_6_10                                                   : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16 : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11 : out   std_logic;
          MSS_READY                                                   : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                        : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE    : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                         : in    std_logic := 'U';
          CertificationSystem_sb_0_AHBmslave5_HREADY                  : in    std_logic := 'U';
          hready_m_xhdl344_7                                          : out   std_logic;
          N_225                                                       : out   std_logic;
          N_276                                                       : out   std_logic;
          N_259                                                       : out   std_logic;
          N_243                                                       : out   std_logic;
          N_236                                                       : out   std_logic;
          N_235                                                       : out   std_logic;
          N_277                                                       : out   std_logic;
          N_255                                                       : out   std_logic;
          N_241                                                       : out   std_logic;
          N_242                                                       : out   std_logic;
          N_244                                                       : out   std_logic;
          N_246                                                       : out   std_logic;
          N_247                                                       : out   std_logic;
          N_256                                                       : out   std_logic;
          N_257                                                       : out   std_logic;
          N_258                                                       : out   std_logic;
          ren_pos                                                     : in    std_logic := 'U';
          hready_m_xhdl343_10                                         : out   std_logic;
          hready_m_xhdl343_11                                         : out   std_logic;
          N_120                                                       : out   std_logic;
          N_216                                                       : in    std_logic := 'U';
          N_215                                                       : in    std_logic := 'U';
          hready_m_xhdl345                                            : out   std_logic;
          N_335                                                       : in    std_logic := 'U';
          N_214                                                       : in    std_logic := 'U';
          N_305                                                       : in    std_logic := 'U';
          N_206                                                       : out   std_logic;
          N_508                                                       : in    std_logic := 'U';
          N_478_i_0                                                   : out   std_logic;
          N_507                                                       : in    std_logic := 'U';
          N_477_i_0                                                   : out   std_logic;
          N_479_i_0                                                   : out   std_logic;
          N_480_i_0                                                   : out   std_logic;
          N_481_i_0                                                   : out   std_logic;
          un8_hreadyin_i_0                                            : in    std_logic := 'U';
          N_9_i_0                                                     : out   std_logic;
          N_226                                                       : out   std_logic;
          defSlaveSMNextState                                         : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                     : in    std_logic := 'U';
          N_63_i_0                                                    : out   std_logic;
          N_62_i_0                                                    : out   std_logic;
          N_60_i_0                                                    : out   std_logic;
          N_98_i_0                                                    : out   std_logic;
          N_96_i_0                                                    : out   std_logic;
          N_94_i_0                                                    : out   std_logic;
          N_92_i_0                                                    : out   std_logic;
          N_90_i_0                                                    : out   std_logic;
          N_88_i_0                                                    : out   std_logic;
          N_86_i_0                                                    : out   std_logic;
          N_84_i_0                                                    : out   std_logic;
          N_82_i_0                                                    : out   std_logic;
          N_80_i_0                                                    : out   std_logic;
          N_78_i_0                                                    : out   std_logic;
          N_76_i_0                                                    : out   std_logic;
          N_74_i_0                                                    : out   std_logic;
          N_72_i_0                                                    : out   std_logic;
          N_70_i_0                                                    : out   std_logic;
          N_68_i_0                                                    : out   std_logic;
          N_66_i_0                                                    : out   std_logic;
          N_64_i_0                                                    : out   std_logic;
          N_58_i_0                                                    : out   std_logic;
          N_56_i_0                                                    : out   std_logic;
          N_54_i_0                                                    : out   std_logic;
          N_52_i_0                                                    : out   std_logic;
          N_50_i_0                                                    : out   std_logic;
          N_48_i_0                                                    : out   std_logic;
          N_46_i_0                                                    : out   std_logic;
          N_44_i_0                                                    : out   std_logic;
          N_42_i_0                                                    : out   std_logic;
          N_40_i_0                                                    : out   std_logic;
          N_38_i_0                                                    : out   std_logic;
          HTRANS_i_a2_0_0                                             : out   std_logic;
          N_271                                                       : in    std_logic := 'U';
          N_157_i_i_o2_0                                              : out   std_logic;
          N_157_i_i_o2_0_out                                          : out   std_logic;
          hsel2_i_4                                                   : out   std_logic;
          N_196_i_0                                                   : out   std_logic;
          N_195_i_0                                                   : out   std_logic;
          N_194_i_0                                                   : out   std_logic;
          N_65_i_0                                                    : out   std_logic;
          N_67_i_0                                                    : out   std_logic;
          N_110_i_0                                                   : out   std_logic;
          N_112_i_0                                                   : out   std_logic;
          N_114_i_0                                                   : out   std_logic;
          N_116_i_0                                                   : out   std_logic;
          N_69_i_0                                                    : out   std_logic;
          N_71_i_0                                                    : out   std_logic;
          N_73_i_0                                                    : out   std_logic;
          N_75_i_0                                                    : out   std_logic;
          N_77_i_0                                                    : out   std_logic;
          N_83_i_0                                                    : out   std_logic;
          N_85_i_0                                                    : out   std_logic;
          N_133_i_0                                                   : out   std_logic;
          N_87_i_0                                                    : out   std_logic;
          N_89_i_0                                                    : out   std_logic;
          N_140_i_0                                                   : out   std_logic;
          N_91_i_0                                                    : out   std_logic;
          N_93_i_0                                                    : out   std_logic;
          N_95_i_0                                                    : out   std_logic;
          N_97_i_0                                                    : out   std_logic;
          N_99_i_0                                                    : out   std_logic;
          N_152_i_0                                                   : out   std_logic;
          N_101_i_0                                                   : out   std_logic;
          N_156_i_0                                                   : out   std_logic;
          N_158_i_0                                                   : out   std_logic;
          N_103_i_0                                                   : out   std_logic;
          N_105_i_0                                                   : out   std_logic;
          N_107_i_0                                                   : out   std_logic;
          N_168_i_0                                                   : out   std_logic;
          N_109_i_0                                                   : out   std_logic;
          N_111_i_0                                                   : out   std_logic;
          N_218_i_0                                                   : out   std_logic;
          N_217_i_0                                                   : out   std_logic;
          N_203_i_0                                                   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CertificationSystem_sb_MSS
    port( CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE     : out   std_logic_vector(1 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS    : out   std_logic_vector(1 to 1);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA    : out   std_logic_vector(31 downto 0);
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP     : in    std_logic_vector(0 to 0) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9   : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31  : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8  : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29 : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30 : in    std_logic := 'U';
          SPI_0_SS0                                                   : inout   std_logic;
          SPI_0_DO                                                    : out   std_logic;
          SPI_0_DI                                                    : in    std_logic := 'U';
          SPI_0_CLK                                                   : inout   std_logic;
          MMUART_1_TXD                                                : out   std_logic;
          MMUART_1_RXD                                                : in    std_logic := 'U';
          CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N       : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE    : out   std_logic;
          CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F            : out   std_logic;
          CertificationSystem_sb_0_GPIO_1_M2F                         : out   std_logic;
          GPIO_0_M2F_c                                                : out   std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F                         : out   std_logic;
          N_481_i_0                                                   : in    std_logic := 'U';
          N_480_i_0                                                   : in    std_logic := 'U';
          N_479_i_0                                                   : in    std_logic := 'U';
          N_478_i_0                                                   : in    std_logic := 'U';
          N_477_i_0                                                   : in    std_logic := 'U';
          N_9_i_0                                                     : in    std_logic := 'U';
          FAB_CCC_LOCK                                                : in    std_logic := 'U';
          SHA256_Module_0_waiting_data                                : in    std_logic := 'U';
          SHA256_Module_0_data_available_lastbank_8                   : in    std_logic := 'U';
          SHA256_Module_0_di_req_o                                    : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o                                  : in    std_logic := 'U';
          SHA256_Module_0_data_available                              : in    std_logic := 'U';
          SHA256_Module_0_error_o                                     : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                        : in    std_logic := 'U'
        );
  end component;

  component CertificationSystem_sb_CCC_0_FCCC
    port( CertificationSystem_sb_0_FAB_CCC_GL0               : out   std_logic;
          FAB_CCC_LOCK                                       : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

  component CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM
    port( CoreAHBLite_0_AHBmslave3_HADDR                          : in    std_logic_vector(11 to 11) := (others => 'U');
          arbRegSMCurrentState                                    : in    std_logic_vector(15 to 15) := (others => 'U');
          CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP : in    std_logic_vector(0 to 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave3_HRDATA                         : out   std_logic_vector(31 downto 0);
          xhdl1222_2                                              : in    std_logic := 'U';
          xhdl1222_0                                              : in    std_logic := 'U';
          SDATASELInt_9                                           : in    std_logic := 'U';
          SDATASELInt_8                                           : in    std_logic := 'U';
          SDATASELInt_7                                           : in    std_logic := 'U';
          SDATASELInt_6                                           : in    std_logic := 'U';
          SDATASELInt_13                                          : in    std_logic := 'U';
          SDATASELInt_12                                          : in    std_logic := 'U';
          SDATASELInt_11                                          : in    std_logic := 'U';
          SDATASELInt_10                                          : in    std_logic := 'U';
          SDATASELInt_4                                           : in    std_logic := 'U';
          SDATASELInt_2                                           : in    std_logic := 'U';
          SDATASELInt_1                                           : in    std_logic := 'U';
          SDATASELInt_0                                           : in    std_logic := 'U';
          MSS_READY                                               : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0                    : in    std_logic := 'U';
          N_236                                                   : in    std_logic := 'U';
          N_271                                                   : out   std_logic;
          N_235                                                   : in    std_logic := 'U';
          N_246                                                   : in    std_logic := 'U';
          N_276                                                   : in    std_logic := 'U';
          N_194_i_0                                               : in    std_logic := 'U';
          N_195_i_0                                               : in    std_logic := 'U';
          N_196_i_0                                               : in    std_logic := 'U';
          N_259                                                   : in    std_logic := 'U';
          N_258                                                   : in    std_logic := 'U';
          N_257                                                   : in    std_logic := 'U';
          N_256                                                   : in    std_logic := 'U';
          N_255                                                   : in    std_logic := 'U';
          N_244                                                   : in    std_logic := 'U';
          N_243                                                   : in    std_logic := 'U';
          N_242                                                   : in    std_logic := 'U';
          N_241                                                   : in    std_logic := 'U';
          N_247                                                   : in    std_logic := 'U';
          N_277                                                   : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave3_HREADY_i_1                     : out   std_logic;
          hready_m_xhdl343_11                                     : in    std_logic := 'U';
          N_305                                                   : out   std_logic;
          hready_m_xhdl343_10                                     : in    std_logic := 'U';
          hready_m_xhdl344_7                                      : in    std_logic := 'U';
          N_335                                                   : out   std_logic;
          N_215                                                   : out   std_logic;
          N_216                                                   : out   std_logic;
          N_214                                                   : out   std_logic;
          CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0                 : out   std_logic;
          N_157_i_i_o2_0                                          : in    std_logic := 'U';
          N_157_i_i_o2_0_out                                      : in    std_logic := 'U';
          CertificationSystem_sb_0_AHBmslave5_HREADY              : in    std_logic := 'U';
          defSlaveSMNextState                                     : in    std_logic := 'U';
          hready_m_xhdl345                                        : in    std_logic := 'U';
          un8_hreadyin_i_0                                        : out   std_logic;
          N_225                                                   : in    std_logic := 'U';
          HTRANS_i_a2_0_0                                         : in    std_logic := 'U';
          N_120                                                   : in    std_logic := 'U';
          hsel2_i_4                                               : in    std_logic := 'U';
          N_38_i_0                                                : in    std_logic := 'U';
          N_40_i_0                                                : in    std_logic := 'U';
          N_42_i_0                                                : in    std_logic := 'U';
          N_44_i_0                                                : in    std_logic := 'U';
          N_46_i_0                                                : in    std_logic := 'U';
          N_48_i_0                                                : in    std_logic := 'U';
          N_50_i_0                                                : in    std_logic := 'U';
          N_52_i_0                                                : in    std_logic := 'U';
          N_54_i_0                                                : in    std_logic := 'U';
          N_56_i_0                                                : in    std_logic := 'U';
          N_58_i_0                                                : in    std_logic := 'U';
          N_64_i_0                                                : in    std_logic := 'U';
          N_66_i_0                                                : in    std_logic := 'U';
          N_68_i_0                                                : in    std_logic := 'U';
          N_70_i_0                                                : in    std_logic := 'U';
          N_72_i_0                                                : in    std_logic := 'U';
          N_74_i_0                                                : in    std_logic := 'U';
          N_76_i_0                                                : in    std_logic := 'U';
          N_78_i_0                                                : in    std_logic := 'U';
          N_80_i_0                                                : in    std_logic := 'U';
          N_82_i_0                                                : in    std_logic := 'U';
          N_84_i_0                                                : in    std_logic := 'U';
          N_86_i_0                                                : in    std_logic := 'U';
          N_88_i_0                                                : in    std_logic := 'U';
          N_90_i_0                                                : in    std_logic := 'U';
          N_92_i_0                                                : in    std_logic := 'U';
          N_94_i_0                                                : in    std_logic := 'U';
          N_96_i_0                                                : in    std_logic := 'U';
          N_98_i_0                                                : in    std_logic := 'U';
          N_60_i_0                                                : in    std_logic := 'U';
          N_62_i_0                                                : in    std_logic := 'U';
          N_63_i_0                                                : in    std_logic := 'U'
        );
  end component;

    signal \CertificationSystem_sb_0_POWER_ON_RESET_N\, 
        \SYSRESET_POR\, \CertificationSystem_sb_0_FAB_CCC_GL0\, 
        FAB_CCC_LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[0]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[1]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[6]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[7]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[8]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[9]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[10]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[11]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[12]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[13]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[14]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[15]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[28]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[29]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[30]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[31]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[0]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[1]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[0]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[1]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[2]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[3]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[4]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[5]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[6]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[7]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[8]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[10]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[11]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[12]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[13]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[14]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[15]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[16]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[17]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[19]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[21]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[22]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[23]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[24]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[25]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[26]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[27]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[29]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[30]\, 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        N_481_i_0, N_480_i_0, N_479_i_0, N_478_i_0, N_477_i_0, 
        N_9_i_0, \xhdl1222[3]\, \xhdl1222_2\, \SDATASELInt[0]\, 
        \SDATASELInt[1]\, \SDATASELInt[2]\, \SDATASELInt[4]\, 
        \SDATASELInt[6]\, \SDATASELInt[7]\, \SDATASELInt[8]\, 
        \SDATASELInt[9]\, \SDATASELInt[10]\, \SDATASELInt[11]\, 
        \SDATASELInt[12]\, \SDATASELInt[13]\, 
        \arbRegSMCurrentState[15]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[0]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[1]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[2]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[3]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[4]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[5]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[6]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[7]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[8]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[9]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[10]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[11]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[12]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[13]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[14]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[15]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[16]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[17]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[18]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[19]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[20]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[21]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[22]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[23]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[24]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[25]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[26]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[27]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[28]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[29]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[30]\, 
        \CoreAHBLite_0_AHBmslave3_HRDATA[31]\, 
        \CoreAHBLite_0_AHBmslave3_HADDR[11]\, MSS_READY, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, hready_m_xhdl344_7, 
        \N_225\, \N_276\, \N_259\, N_243, N_236, N_235, \N_277\, 
        N_255, N_241, N_242, N_244, N_246, N_247, N_256, N_257, 
        N_258, hready_m_xhdl343_10, hready_m_xhdl343_11, N_120, 
        N_216, N_215, hready_m_xhdl345, N_335, N_214, N_305, 
        \un8_hreadyin_i_0\, defSlaveSMNextState, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, N_63_i_0, 
        N_62_i_0, N_60_i_0, N_98_i_0, N_96_i_0, N_94_i_0, 
        N_92_i_0, N_90_i_0, N_88_i_0, N_86_i_0, N_84_i_0, 
        N_82_i_0, N_80_i_0, N_78_i_0, N_76_i_0, N_74_i_0, 
        N_72_i_0, N_70_i_0, N_68_i_0, N_66_i_0, N_64_i_0, 
        N_58_i_0, N_56_i_0, N_54_i_0, N_52_i_0, N_50_i_0, 
        N_48_i_0, N_46_i_0, N_44_i_0, N_42_i_0, N_40_i_0, 
        N_38_i_0, HTRANS_i_a2_0_0, N_271, N_157_i_i_o2_0, 
        N_157_i_i_o2_0_out, hsel2_i_4, N_196_i_0, N_195_i_0, 
        N_194_i_0, GND_net_1, VCC_net_1 : std_logic;

    for all : CertificationSystem_sb_FABOSC_0_OSC
	Use entity work.CertificationSystem_sb_FABOSC_0_OSC(DEF_ARCH);
    for all : CoreResetP
	Use entity work.CoreResetP(DEF_ARCH);
    for all : CoreAHBLite
	Use entity work.CoreAHBLite(DEF_ARCH);
    for all : CertificationSystem_sb_MSS
	Use entity work.CertificationSystem_sb_MSS(DEF_ARCH);
    for all : CertificationSystem_sb_CCC_0_FCCC
	Use entity work.CertificationSystem_sb_CCC_0_FCCC(DEF_ARCH);
    for all : CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM
	Use entity work.
        CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM(DEF_ARCH);
begin 

    xhdl1222_2 <= \xhdl1222_2\;
    CertificationSystem_sb_0_POWER_ON_RESET_N <= 
        \CertificationSystem_sb_0_POWER_ON_RESET_N\;
    CertificationSystem_sb_0_FAB_CCC_GL0 <= 
        \CertificationSystem_sb_0_FAB_CCC_GL0\;
    N_225 <= \N_225\;
    N_276 <= \N_276\;
    N_259 <= \N_259\;
    N_277 <= \N_277\;
    un8_hreadyin_i_0 <= \un8_hreadyin_i_0\;

    FABOSC_0 : CertificationSystem_sb_FABOSC_0_OSC
      port map(FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
         => FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    CORERESETP_0 : CoreResetP
      port map(MSS_READY => MSS_READY, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        \CertificationSystem_sb_0_FAB_CCC_GL0\, 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        CertificationSystem_sb_0_POWER_ON_RESET_N => 
        \CertificationSystem_sb_0_POWER_ON_RESET_N\);
    
    CoreAHBLite_0 : CoreAHBLite
      port map(
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[0]\, 
        arbRegSMCurrentState(15) => \arbRegSMCurrentState[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        result_addr_net_0(3) => result_addr_net_0(3), 
        result_addr_net_0(2) => result_addr_net_0(2), 
        result_addr_net_0(1) => result_addr_net_0(1), 
        result_addr_net_0(0) => result_addr_net_0(0), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(31) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[31]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(30) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[30]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(29) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[29]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(28) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[28]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(27) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[27]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(26) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[26]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(25) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[25]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(24) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[24]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(23) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[23]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(22) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[22]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(21) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[21]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(20) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[20]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(19) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[19]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(18) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[18]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(17) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[17]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(16) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[16]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(15) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[15]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(14) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[14]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(13) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[13]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(12) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[12]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(11) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[11]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(10) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[10]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(9) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[9]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(8) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[8]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(7) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[7]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(6) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[6]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(5) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[5]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(4) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[4]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(3) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[3]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(2) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[2]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(1) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[1]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(0) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[0]\, line_7(2) => 
        line_7(2), line_7(1) => line_7(1), 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        CoreAHBLite_0_AHBmslave3_HADDR(11) => 
        \CoreAHBLite_0_AHBmslave3_HADDR[11]\, xhdl1222_0 => 
        \xhdl1222[3]\, xhdl1222_2 => \xhdl1222_2\, SDATASELInt_0
         => \SDATASELInt[0]\, SDATASELInt_1 => \SDATASELInt[1]\, 
        SDATASELInt_2 => \SDATASELInt[2]\, SDATASELInt_4 => 
        \SDATASELInt[4]\, SDATASELInt_6 => \SDATASELInt[6]\, 
        SDATASELInt_7 => \SDATASELInt[7]\, SDATASELInt_8 => 
        \SDATASELInt[8]\, SDATASELInt_9 => \SDATASELInt[9]\, 
        SDATASELInt_10 => \SDATASELInt[10]\, SDATASELInt_11 => 
        \SDATASELInt[11]\, SDATASELInt_12 => \SDATASELInt[12]\, 
        SDATASELInt_13 => \SDATASELInt[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[11]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[12]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[14]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[29]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[30]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[6]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[7]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[8]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[9]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[10]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[28]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[31]\, 
        line_13 => line_13, line_10 => line_10, line_21 => 
        line_21, line_24 => line_24, line_18 => line_18, line_23
         => line_23, line_16 => line_16, line_28 => line_28, 
        line_9 => line_9, line_3_d0 => line_3_d0, line_5_d0 => 
        line_5_d0, line_15 => line_15, line_26 => line_26, 
        line_14 => line_14, line_20 => line_20, line_2_d0 => 
        line_2_d0, line_25 => line_25, line_29 => line_29, 
        line_19 => line_19, line_27 => line_27, line_30 => 
        line_30, line_17 => line_17, line_8 => line_8, line_0_d0
         => line_0_d0, line_6_d0 => line_6_d0, line_1_d0 => 
        line_1_d0, line_0_10 => line_0_10, line_0_21 => line_0_21, 
        line_0_24 => line_0_24, line_0_18 => line_0_18, line_0_23
         => line_0_23, line_0_16 => line_0_16, line_0_28 => 
        line_0_28, line_0_9 => line_0_9, line_0_3 => line_0_3, 
        line_0_5 => line_0_5, line_0_15 => line_0_15, line_0_26
         => line_0_26, line_0_14 => line_0_14, line_0_20 => 
        line_0_20, line_0_2 => line_0_2, line_0_25 => line_0_25, 
        line_0_29 => line_0_29, line_0_19 => line_0_19, line_0_27
         => line_0_27, line_0_30 => line_0_30, line_0_17 => 
        line_0_17, line_0_8 => line_0_8, line_0_0 => line_0_0, 
        line_0_1 => line_0_1, line_0_6 => line_0_6, line_0_13 => 
        line_0_13, line_1_10 => line_1_10, line_1_21 => line_1_21, 
        line_1_24 => line_1_24, line_1_18 => line_1_18, line_1_23
         => line_1_23, line_1_16 => line_1_16, line_1_28 => 
        line_1_28, line_1_9 => line_1_9, line_1_3 => line_1_3, 
        line_1_5 => line_1_5, line_1_15 => line_1_15, line_1_26
         => line_1_26, line_1_14 => line_1_14, line_1_20 => 
        line_1_20, line_1_2 => line_1_2, line_1_25 => line_1_25, 
        line_1_29 => line_1_29, line_1_19 => line_1_19, line_1_27
         => line_1_27, line_1_30 => line_1_30, line_1_17 => 
        line_1_17, line_1_8 => line_1_8, line_1_0 => line_1_0, 
        line_1_1 => line_1_1, line_1_6 => line_1_6, line_1_13 => 
        line_1_13, line_2_19 => line_2_19, line_2_27 => line_2_27, 
        line_2_30 => line_2_30, line_2_17 => line_2_17, line_2_8
         => line_2_8, line_2_10 => line_2_10, line_2_15 => 
        line_2_15, line_2_26 => line_2_26, line_2_20 => line_2_20, 
        line_2_0 => line_2_0, line_2_1 => line_2_1, line_2_29 => 
        line_2_29, line_2_25 => line_2_25, line_2_2 => line_2_2, 
        line_2_6 => line_2_6, line_2_13 => line_2_13, line_2_14
         => line_2_14, line_2_5 => line_2_5, line_2_3 => line_2_3, 
        line_2_9 => line_2_9, line_2_28 => line_2_28, line_2_16
         => line_2_16, line_2_23 => line_2_23, line_2_18 => 
        line_2_18, line_2_24 => line_2_24, line_2_21 => line_2_21, 
        line_3_19 => line_3_19, line_3_17 => line_3_17, line_3_8
         => line_3_8, line_3_0 => line_3_0, line_3_1 => line_3_1, 
        line_3_29 => line_3_29, line_3_25 => line_3_25, line_3_2
         => line_3_2, line_3_20 => line_3_20, line_3_6 => 
        line_3_6, line_3_13 => line_3_13, line_3_14 => line_3_14, 
        line_3_26 => line_3_26, line_3_15 => line_3_15, line_3_5
         => line_3_5, line_3_3 => line_3_3, line_3_9 => line_3_9, 
        line_3_28 => line_3_28, line_3_16 => line_3_16, line_3_23
         => line_3_23, line_3_18 => line_3_18, line_3_24 => 
        line_3_24, line_3_21 => line_3_21, line_3_10 => line_3_10, 
        SHA256_Module_0_data_out_5 => SHA256_Module_0_data_out_5, 
        SHA256_Module_0_data_out_13 => 
        SHA256_Module_0_data_out_13, SHA256_Module_0_data_out_12
         => SHA256_Module_0_data_out_12, 
        SHA256_Module_0_data_out_8 => SHA256_Module_0_data_out_8, 
        SHA256_Module_0_data_out_23 => 
        SHA256_Module_0_data_out_23, SHA256_Module_0_data_out_0
         => SHA256_Module_0_data_out_0, line_4_19 => line_4_19, 
        line_4_17 => line_4_17, line_4_8 => line_4_8, line_4_0
         => line_4_0, line_4_1 => line_4_1, line_4_29 => 
        line_4_29, line_4_25 => line_4_25, line_4_2 => line_4_2, 
        line_4_20 => line_4_20, line_4_14 => line_4_14, line_4_26
         => line_4_26, line_4_15 => line_4_15, line_4_5 => 
        line_4_5, line_4_3 => line_4_3, line_4_9 => line_4_9, 
        line_4_28 => line_4_28, line_4_16 => line_4_16, line_4_23
         => line_4_23, line_4_18 => line_4_18, line_4_24 => 
        line_4_24, line_4_21 => line_4_21, line_4_10 => line_4_10, 
        line_4_6 => line_4_6, line_4_13 => line_4_13, line_5_19
         => line_5_19, line_5_17 => line_5_17, line_5_8 => 
        line_5_8, line_5_0 => line_5_0, line_5_1 => line_5_1, 
        line_5_29 => line_5_29, line_5_25 => line_5_25, line_5_2
         => line_5_2, line_5_20 => line_5_20, line_5_6 => 
        line_5_6, line_5_13 => line_5_13, line_5_14 => line_5_14, 
        line_5_26 => line_5_26, line_5_15 => line_5_15, line_5_5
         => line_5_5, line_5_3 => line_5_3, line_5_9 => line_5_9, 
        line_5_28 => line_5_28, line_5_16 => line_5_16, line_5_23
         => line_5_23, line_5_18 => line_5_18, line_5_24 => 
        line_5_24, line_5_21 => line_5_21, line_5_10 => line_5_10, 
        line_6_19 => line_6_19, line_6_17 => line_6_17, line_6_8
         => line_6_8, line_6_0 => line_6_0, line_6_1 => line_6_1, 
        line_6_29 => line_6_29, line_6_25 => line_6_25, line_6_2
         => line_6_2, line_6_20 => line_6_20, line_6_6 => 
        line_6_6, line_6_13 => line_6_13, line_6_14 => line_6_14, 
        line_6_26 => line_6_26, line_6_15 => line_6_15, line_6_5
         => line_6_5, line_6_3 => line_6_3, line_6_9 => line_6_9, 
        line_6_28 => line_6_28, line_6_16 => line_6_16, line_6_23
         => line_6_23, line_6_18 => line_6_18, line_6_24 => 
        line_6_24, line_6_21 => line_6_21, line_6_10 => line_6_10, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[5]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[12]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[8]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[23]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[10]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[6]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[25]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[17]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[19]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[21]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[24]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[26]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[29]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[30]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[4]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[7]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[22]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[27]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[14]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[16]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[11]\, 
        MSS_READY => MSS_READY, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        \CertificationSystem_sb_0_FAB_CCC_GL0\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, 
        CertificationSystem_sb_0_AHBmslave5_HREADY => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, 
        hready_m_xhdl344_7 => hready_m_xhdl344_7, N_225 => 
        \N_225\, N_276 => \N_276\, N_259 => \N_259\, N_243 => 
        N_243, N_236 => N_236, N_235 => N_235, N_277 => \N_277\, 
        N_255 => N_255, N_241 => N_241, N_242 => N_242, N_244 => 
        N_244, N_246 => N_246, N_247 => N_247, N_256 => N_256, 
        N_257 => N_257, N_258 => N_258, ren_pos => ren_pos, 
        hready_m_xhdl343_10 => hready_m_xhdl343_10, 
        hready_m_xhdl343_11 => hready_m_xhdl343_11, N_120 => 
        N_120, N_216 => N_216, N_215 => N_215, hready_m_xhdl345
         => hready_m_xhdl345, N_335 => N_335, N_214 => N_214, 
        N_305 => N_305, N_206 => N_206, N_508 => N_508, N_478_i_0
         => N_478_i_0, N_507 => N_507, N_477_i_0 => N_477_i_0, 
        N_479_i_0 => N_479_i_0, N_480_i_0 => N_480_i_0, N_481_i_0
         => N_481_i_0, un8_hreadyin_i_0 => \un8_hreadyin_i_0\, 
        N_9_i_0 => N_9_i_0, N_226 => N_226, defSlaveSMNextState
         => defSlaveSMNextState, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, N_63_i_0 => 
        N_63_i_0, N_62_i_0 => N_62_i_0, N_60_i_0 => N_60_i_0, 
        N_98_i_0 => N_98_i_0, N_96_i_0 => N_96_i_0, N_94_i_0 => 
        N_94_i_0, N_92_i_0 => N_92_i_0, N_90_i_0 => N_90_i_0, 
        N_88_i_0 => N_88_i_0, N_86_i_0 => N_86_i_0, N_84_i_0 => 
        N_84_i_0, N_82_i_0 => N_82_i_0, N_80_i_0 => N_80_i_0, 
        N_78_i_0 => N_78_i_0, N_76_i_0 => N_76_i_0, N_74_i_0 => 
        N_74_i_0, N_72_i_0 => N_72_i_0, N_70_i_0 => N_70_i_0, 
        N_68_i_0 => N_68_i_0, N_66_i_0 => N_66_i_0, N_64_i_0 => 
        N_64_i_0, N_58_i_0 => N_58_i_0, N_56_i_0 => N_56_i_0, 
        N_54_i_0 => N_54_i_0, N_52_i_0 => N_52_i_0, N_50_i_0 => 
        N_50_i_0, N_48_i_0 => N_48_i_0, N_46_i_0 => N_46_i_0, 
        N_44_i_0 => N_44_i_0, N_42_i_0 => N_42_i_0, N_40_i_0 => 
        N_40_i_0, N_38_i_0 => N_38_i_0, HTRANS_i_a2_0_0 => 
        HTRANS_i_a2_0_0, N_271 => N_271, N_157_i_i_o2_0 => 
        N_157_i_i_o2_0, N_157_i_i_o2_0_out => N_157_i_i_o2_0_out, 
        hsel2_i_4 => hsel2_i_4, N_196_i_0 => N_196_i_0, N_195_i_0
         => N_195_i_0, N_194_i_0 => N_194_i_0, N_65_i_0 => 
        N_65_i_0, N_67_i_0 => N_67_i_0, N_110_i_0 => N_110_i_0, 
        N_112_i_0 => N_112_i_0, N_114_i_0 => N_114_i_0, N_116_i_0
         => N_116_i_0, N_69_i_0 => N_69_i_0, N_71_i_0 => N_71_i_0, 
        N_73_i_0 => N_73_i_0, N_75_i_0 => N_75_i_0, N_77_i_0 => 
        N_77_i_0, N_83_i_0 => N_83_i_0, N_85_i_0 => N_85_i_0, 
        N_133_i_0 => N_133_i_0, N_87_i_0 => N_87_i_0, N_89_i_0
         => N_89_i_0, N_140_i_0 => N_140_i_0, N_91_i_0 => 
        N_91_i_0, N_93_i_0 => N_93_i_0, N_95_i_0 => N_95_i_0, 
        N_97_i_0 => N_97_i_0, N_99_i_0 => N_99_i_0, N_152_i_0 => 
        N_152_i_0, N_101_i_0 => N_101_i_0, N_156_i_0 => N_156_i_0, 
        N_158_i_0 => N_158_i_0, N_103_i_0 => N_103_i_0, N_105_i_0
         => N_105_i_0, N_107_i_0 => N_107_i_0, N_168_i_0 => 
        N_168_i_0, N_109_i_0 => N_109_i_0, N_111_i_0 => N_111_i_0, 
        N_218_i_0 => N_218_i_0, N_217_i_0 => N_217_i_0, N_203_i_0
         => N_203_i_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    CertificationSystem_sb_MSS_0 : CertificationSystem_sb_MSS
      port map(
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HSIZE[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HTRANS[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(31)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[31]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(30)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[30]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(29)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[29]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(28)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[28]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(27)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[27]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(26)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[26]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(25)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[25]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(24)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[24]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(23)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[23]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(22)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[22]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(21)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[21]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(20)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[20]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(19)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[19]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(18)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[18]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(17)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[17]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(16)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[16]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(15)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(14)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[14]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(13)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(12)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[12]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(11)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[11]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(10)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[10]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(9)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[9]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(8)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[8]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(7)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[7]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(6)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[6]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(5)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[5]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(4)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[4]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(3)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(2)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(1)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWDATA[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_0
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_1
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_2
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_3
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_4
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[4]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_5
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[5]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_6
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[6]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_7
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[7]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_8
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[8]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_9
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[9]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_10
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[10]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_11
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[11]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_12
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[12]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_13
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_14
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[14]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_15
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_28
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[28]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_29
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[29]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_30
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[30]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR_31
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HADDR[31]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_0
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[0]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_1
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[1]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_2
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[2]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_3
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[3]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_4
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[4]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_5
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[5]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_6
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[6]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_7
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[7]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_8
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[8]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_10
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[10]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_11
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[11]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_12
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[12]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_13
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[13]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_14
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[14]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_15
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_16
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[16]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_17
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[17]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_19
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[19]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_21
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[21]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_22
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[22]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_23
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[23]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_24
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[24]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_25
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[25]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_26
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[26]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_27
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[27]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_29
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[29]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA_30
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRDATA[30]\, 
        SPI_0_SS0 => SPI_0_SS0, SPI_0_DO => SPI_0_DO, SPI_0_DI
         => SPI_0_DI, SPI_0_CLK => SPI_0_CLK, MMUART_1_TXD => 
        MMUART_1_TXD, MMUART_1_RXD => MMUART_1_RXD, 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        CertificationSystem_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE
         => 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HWRITE, 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        CertificationSystem_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        CertificationSystem_sb_0_GPIO_1_M2F => 
        CertificationSystem_sb_0_GPIO_1_M2F, GPIO_0_M2F_c => 
        GPIO_0_M2F_c, CertificationSystem_sb_0_GPIO_9_M2F => 
        CertificationSystem_sb_0_GPIO_9_M2F, N_481_i_0 => 
        N_481_i_0, N_480_i_0 => N_480_i_0, N_479_i_0 => N_479_i_0, 
        N_478_i_0 => N_478_i_0, N_477_i_0 => N_477_i_0, N_9_i_0
         => N_9_i_0, FAB_CCC_LOCK => FAB_CCC_LOCK, 
        SHA256_Module_0_waiting_data => 
        SHA256_Module_0_waiting_data, 
        SHA256_Module_0_data_available_lastbank_8 => 
        SHA256_Module_0_data_available_lastbank_8, 
        SHA256_Module_0_di_req_o => SHA256_Module_0_di_req_o, 
        SHA256_Module_0_do_valid_o => SHA256_Module_0_do_valid_o, 
        SHA256_Module_0_data_available => 
        SHA256_Module_0_data_available, SHA256_Module_0_error_o
         => SHA256_Module_0_error_o, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        \CertificationSystem_sb_0_FAB_CCC_GL0\);
    
    CCC_0 : CertificationSystem_sb_CCC_0_FCCC
      port map(CertificationSystem_sb_0_FAB_CCC_GL0 => 
        \CertificationSystem_sb_0_FAB_CCC_GL0\, FAB_CCC_LOCK => 
        FAB_CCC_LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    SYSRESET_POR_RNIC1R5 : CLKINT
      port map(A => \SYSRESET_POR\, Y => 
        \CertificationSystem_sb_0_POWER_ON_RESET_N\);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => \SYSRESET_POR\, DEVRST_N => 
        DEVRST_N);
    
    COREAHBLSRAM_0_0 : 
        CertificationSystem_sb_COREAHBLSRAM_0_0_COREAHBLSRAM
      port map(CoreAHBLite_0_AHBmslave3_HADDR(11) => 
        \CoreAHBLite_0_AHBmslave3_HADDR[11]\, 
        arbRegSMCurrentState(15) => \arbRegSMCurrentState[15]\, 
        CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP(0)
         => 
        \CertificationSystem_sb_MSS_TMP_0_FIC_0_AHB_MASTER_HRESP[0]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(31) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[31]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(30) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[30]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(29) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[29]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(28) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[28]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(27) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[27]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(26) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[26]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(25) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[25]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(24) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[24]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(23) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[23]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(22) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[22]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(21) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[21]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(20) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[20]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(19) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[19]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(18) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[18]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(17) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[17]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(16) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[16]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(15) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[15]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(14) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[14]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(13) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[13]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(12) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[12]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(11) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[11]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(10) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[10]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(9) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[9]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(8) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[8]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(7) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[7]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(6) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[6]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(5) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[5]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(4) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[4]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(3) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[3]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(2) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[2]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(1) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[1]\, 
        CoreAHBLite_0_AHBmslave3_HRDATA(0) => 
        \CoreAHBLite_0_AHBmslave3_HRDATA[0]\, xhdl1222_2 => 
        \xhdl1222_2\, xhdl1222_0 => \xhdl1222[3]\, SDATASELInt_9
         => \SDATASELInt[9]\, SDATASELInt_8 => \SDATASELInt[8]\, 
        SDATASELInt_7 => \SDATASELInt[7]\, SDATASELInt_6 => 
        \SDATASELInt[6]\, SDATASELInt_13 => \SDATASELInt[13]\, 
        SDATASELInt_12 => \SDATASELInt[12]\, SDATASELInt_11 => 
        \SDATASELInt[11]\, SDATASELInt_10 => \SDATASELInt[10]\, 
        SDATASELInt_4 => \SDATASELInt[4]\, SDATASELInt_2 => 
        \SDATASELInt[2]\, SDATASELInt_1 => \SDATASELInt[1]\, 
        SDATASELInt_0 => \SDATASELInt[0]\, MSS_READY => MSS_READY, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        \CertificationSystem_sb_0_FAB_CCC_GL0\, N_236 => N_236, 
        N_271 => N_271, N_235 => N_235, N_246 => N_246, N_276 => 
        \N_276\, N_194_i_0 => N_194_i_0, N_195_i_0 => N_195_i_0, 
        N_196_i_0 => N_196_i_0, N_259 => \N_259\, N_258 => N_258, 
        N_257 => N_257, N_256 => N_256, N_255 => N_255, N_244 => 
        N_244, N_243 => N_243, N_242 => N_242, N_241 => N_241, 
        N_247 => N_247, N_277 => \N_277\, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1, hready_m_xhdl343_11
         => hready_m_xhdl343_11, N_305 => N_305, 
        hready_m_xhdl343_10 => hready_m_xhdl343_10, 
        hready_m_xhdl344_7 => hready_m_xhdl344_7, N_335 => N_335, 
        N_215 => N_215, N_216 => N_216, N_214 => N_214, 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0 => 
        CoreAHBLite_0_AHBmslave3_HREADY_i_1_i_0, N_157_i_i_o2_0
         => N_157_i_i_o2_0, N_157_i_i_o2_0_out => 
        N_157_i_i_o2_0_out, 
        CertificationSystem_sb_0_AHBmslave5_HREADY => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, 
        defSlaveSMNextState => defSlaveSMNextState, 
        hready_m_xhdl345 => hready_m_xhdl345, un8_hreadyin_i_0
         => \un8_hreadyin_i_0\, N_225 => \N_225\, HTRANS_i_a2_0_0
         => HTRANS_i_a2_0_0, N_120 => N_120, hsel2_i_4 => 
        hsel2_i_4, N_38_i_0 => N_38_i_0, N_40_i_0 => N_40_i_0, 
        N_42_i_0 => N_42_i_0, N_44_i_0 => N_44_i_0, N_46_i_0 => 
        N_46_i_0, N_48_i_0 => N_48_i_0, N_50_i_0 => N_50_i_0, 
        N_52_i_0 => N_52_i_0, N_54_i_0 => N_54_i_0, N_56_i_0 => 
        N_56_i_0, N_58_i_0 => N_58_i_0, N_64_i_0 => N_64_i_0, 
        N_66_i_0 => N_66_i_0, N_68_i_0 => N_68_i_0, N_70_i_0 => 
        N_70_i_0, N_72_i_0 => N_72_i_0, N_74_i_0 => N_74_i_0, 
        N_76_i_0 => N_76_i_0, N_78_i_0 => N_78_i_0, N_80_i_0 => 
        N_80_i_0, N_82_i_0 => N_82_i_0, N_84_i_0 => N_84_i_0, 
        N_86_i_0 => N_86_i_0, N_88_i_0 => N_88_i_0, N_90_i_0 => 
        N_90_i_0, N_92_i_0 => N_92_i_0, N_94_i_0 => N_94_i_0, 
        N_96_i_0 => N_96_i_0, N_98_i_0 => N_98_i_0, N_60_i_0 => 
        N_60_i_0, N_62_i_0 => N_62_i_0, N_63_i_0 => N_63_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity AHB_slave_dummy is

    port( waddr_in_net_0                             : out   std_logic_vector(4 downto 0);
          result_addr_net_0                          : out   std_logic_vector(3 downto 0);
          xhdl1222                                   : in    std_logic_vector(5 to 5);
          CertificationSystem_sb_0_POWER_ON_RESET_N  : in    std_logic;
          CertificationSystem_sb_0_FAB_CCC_GL0       : in    std_logic;
          N_276                                      : in    std_logic;
          N_203_i_0                                  : in    std_logic;
          N_217_i_0                                  : in    std_logic;
          N_218_i_0                                  : in    std_logic;
          N_259                                      : in    std_logic;
          CertificationSystem_sb_0_AHBmslave5_HREADY : out   std_logic;
          AHB_slave_dummy_0_write_en                 : out   std_logic;
          AHB_slave_dummy_0_read_en                  : out   std_logic;
          N_277                                      : in    std_logic;
          N_225                                      : in    std_logic;
          N_206                                      : in    std_logic;
          un8_hreadyin_i_0                           : in    std_logic;
          N_226                                      : in    std_logic
        );

end AHB_slave_dummy;

architecture DEF_ARCH of AHB_slave_dummy is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, N_222_i_0, GND_net_1, N_221_i_0, 
        \CertificationSystem_sb_0_AHBmslave5_HREADY\, 
        \ready_ldmx\, N_311_i_0, \AHB_slave_dummy_0_write_en\, 
        \write_en_ldmx\, \AHB_slave_dummy_0_read_en\, 
        \read_en_ldmx\, \hwrite_r\, N_279_i_0, \FSM[0]_net_1\, 
        \FSM[1]_net_1\, \FSM_ns[1]\, 
        \un1_lsram_raddr_1_sqmuxa_i_o3_2_1\, N_314, 
        \lsram_raddr_1_sqmuxa_i_o2_0\ : std_logic;

begin 

    CertificationSystem_sb_0_AHBmslave5_HREADY <= 
        \CertificationSystem_sb_0_AHBmslave5_HREADY\;
    AHB_slave_dummy_0_write_en <= \AHB_slave_dummy_0_write_en\;
    AHB_slave_dummy_0_read_en <= \AHB_slave_dummy_0_read_en\;

    ready_ldmx : CFG4
      generic map(INIT => x"FA22")

      port map(A => \FSM[0]_net_1\, B => \hwrite_r\, C => N_277, 
        D => \CertificationSystem_sb_0_AHBmslave5_HREADY\, Y => 
        \ready_ldmx\);
    
    \lsram_raddr[2]\ : SLE
      port map(D => N_217_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_221_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => result_addr_net_0(2));
    
    hwrite_r : SLE
      port map(D => N_277, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_279_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \hwrite_r\);
    
    \FSM[1]\ : SLE
      port map(D => \FSM_ns[1]\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FSM[1]_net_1\);
    
    \lsram_waddr[0]\ : SLE
      port map(D => N_276, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_222_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => waddr_in_net_0(0));
    
    write_en_ldmx : CFG4
      generic map(INIT => x"54F4")

      port map(A => \FSM[0]_net_1\, B => N_277, C => 
        \AHB_slave_dummy_0_write_en\, D => \hwrite_r\, Y => 
        \write_en_ldmx\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \lsram_raddr[1]\ : SLE
      port map(D => N_203_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_221_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => result_addr_net_0(1));
    
    lsram_raddr_1_sqmuxa_i_o2_0_RNI1UDV_0 : CFG3
      generic map(INIT => x"01")

      port map(A => N_226, B => N_277, C => 
        \lsram_raddr_1_sqmuxa_i_o2_0\, Y => N_221_i_0);
    
    \lsram_waddr[1]\ : SLE
      port map(D => N_203_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_222_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => waddr_in_net_0(1));
    
    lsram_raddr_1_sqmuxa_i_o2_0_RNIMURK : CFG2
      generic map(INIT => x"1")

      port map(A => N_226, B => \lsram_raddr_1_sqmuxa_i_o2_0\, Y
         => N_279_i_0);
    
    \lsram_raddr[0]\ : SLE
      port map(D => N_276, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_221_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => result_addr_net_0(0));
    
    lsram_raddr_1_sqmuxa_i_o2_0_RNI1UDV : CFG3
      generic map(INIT => x"04")

      port map(A => N_226, B => N_277, C => 
        \lsram_raddr_1_sqmuxa_i_o2_0\, Y => N_222_i_0);
    
    \lsram_waddr[3]\ : SLE
      port map(D => N_218_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_222_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => waddr_in_net_0(3));
    
    \FSM_ns_0_a2_0_a2[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \FSM[0]_net_1\, B => \hwrite_r\, Y => 
        \FSM_ns[1]\);
    
    un1_lsram_raddr_1_sqmuxa_i_o3_2_1_RNIBAEP : CFG4
      generic map(INIT => x"F0F1")

      port map(A => \un1_lsram_raddr_1_sqmuxa_i_o3_2_1\, B => 
        N_226, C => \FSM[0]_net_1\, D => N_314, Y => N_311_i_0);
    
    \FSM[0]\ : SLE
      port map(D => N_279_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FSM[0]_net_1\);
    
    un1_lsram_raddr_1_sqmuxa_i_a3 : CFG3
      generic map(INIT => x"0E")

      port map(A => N_206, B => un8_hreadyin_i_0, C => 
        xhdl1222(5), Y => N_314);
    
    un1_lsram_raddr_1_sqmuxa_i_o3_2_1 : CFG3
      generic map(INIT => x"BF")

      port map(A => \FSM[1]_net_1\, B => 
        \CertificationSystem_sb_0_AHBmslave5_HREADY\, C => N_225, 
        Y => \un1_lsram_raddr_1_sqmuxa_i_o3_2_1\);
    
    lsram_raddr_1_sqmuxa_i_o2_0 : CFG3
      generic map(INIT => x"FE")

      port map(A => \un1_lsram_raddr_1_sqmuxa_i_o3_2_1\, B => 
        \FSM[0]_net_1\, C => N_314, Y => 
        \lsram_raddr_1_sqmuxa_i_o2_0\);
    
    write_en : SLE
      port map(D => \write_en_ldmx\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_311_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AHB_slave_dummy_0_write_en\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    read_en : SLE
      port map(D => \read_en_ldmx\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_311_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AHB_slave_dummy_0_read_en\);
    
    ready : SLE
      port map(D => \ready_ldmx\, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_311_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        \CertificationSystem_sb_0_AHBmslave5_HREADY\);
    
    \lsram_raddr[3]\ : SLE
      port map(D => N_218_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_221_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => result_addr_net_0(3));
    
    \lsram_waddr[4]\ : SLE
      port map(D => N_259, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_222_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => waddr_in_net_0(4));
    
    \lsram_waddr[2]\ : SLE
      port map(D => N_217_i_0, CLK => 
        CertificationSystem_sb_0_FAB_CCC_GL0, EN => N_222_i_0, 
        ALn => CertificationSystem_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => waddr_in_net_0(2));
    
    read_en_ldmx : CFG4
      generic map(INIT => x"F151")

      port map(A => \FSM[0]_net_1\, B => N_277, C => 
        \AHB_slave_dummy_0_read_en\, D => \hwrite_r\, Y => 
        \read_en_ldmx\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CertificationSystem is

    port( DEVRST_N     : in    std_logic;
          MMUART_1_RXD : in    std_logic;
          SPI_0_DI     : in    std_logic;
          GPIO_0_M2F   : out   std_logic;
          MMUART_1_TXD : out   std_logic;
          SPI_0_DO     : out   std_logic;
          SPI_0_CLK    : inout std_logic := 'Z';
          SPI_0_SS0    : inout std_logic := 'Z'
        );

end CertificationSystem;

architecture DEF_ARCH of CertificationSystem is 

  component SHA256_Module
    port( result_addr_net_0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          line_7                                    : out   std_logic_vector(2 downto 1);
          waddr_in_net_0                            : in    std_logic_vector(4 downto 0) := (others => 'U');
          SHA256_Module_0_data_out_5                : out   std_logic;
          SHA256_Module_0_data_out_13               : out   std_logic;
          SHA256_Module_0_data_out_12               : out   std_logic;
          SHA256_Module_0_data_out_23               : out   std_logic;
          SHA256_Module_0_data_out_8                : out   std_logic;
          SHA256_Module_0_data_out_0                : out   std_logic;
          line_0_d0                                 : out   std_logic;
          line_1_d0                                 : out   std_logic;
          line_2_d0                                 : out   std_logic;
          line_3_d0                                 : out   std_logic;
          line_5_d0                                 : out   std_logic;
          line_6_d0                                 : out   std_logic;
          line_8                                    : out   std_logic;
          line_9                                    : out   std_logic;
          line_10                                   : out   std_logic;
          line_13                                   : out   std_logic;
          line_14                                   : out   std_logic;
          line_15                                   : out   std_logic;
          line_16                                   : out   std_logic;
          line_17                                   : out   std_logic;
          line_18                                   : out   std_logic;
          line_19                                   : out   std_logic;
          line_20                                   : out   std_logic;
          line_21                                   : out   std_logic;
          line_23                                   : out   std_logic;
          line_24                                   : out   std_logic;
          line_25                                   : out   std_logic;
          line_26                                   : out   std_logic;
          line_28                                   : out   std_logic;
          line_29                                   : out   std_logic;
          line_27                                   : out   std_logic;
          line_30                                   : out   std_logic;
          line_3_0                                  : out   std_logic;
          line_3_1                                  : out   std_logic;
          line_3_2                                  : out   std_logic;
          line_3_3                                  : out   std_logic;
          line_3_5                                  : out   std_logic;
          line_3_6                                  : out   std_logic;
          line_3_8                                  : out   std_logic;
          line_3_9                                  : out   std_logic;
          line_3_10                                 : out   std_logic;
          line_3_13                                 : out   std_logic;
          line_3_14                                 : out   std_logic;
          line_3_15                                 : out   std_logic;
          line_3_16                                 : out   std_logic;
          line_3_17                                 : out   std_logic;
          line_3_18                                 : out   std_logic;
          line_3_19                                 : out   std_logic;
          line_3_20                                 : out   std_logic;
          line_3_21                                 : out   std_logic;
          line_3_23                                 : out   std_logic;
          line_3_24                                 : out   std_logic;
          line_3_25                                 : out   std_logic;
          line_3_26                                 : out   std_logic;
          line_3_28                                 : out   std_logic;
          line_3_29                                 : out   std_logic;
          line_0_0                                  : out   std_logic;
          line_0_1                                  : out   std_logic;
          line_0_2                                  : out   std_logic;
          line_0_3                                  : out   std_logic;
          line_0_5                                  : out   std_logic;
          line_0_6                                  : out   std_logic;
          line_0_8                                  : out   std_logic;
          line_0_9                                  : out   std_logic;
          line_0_10                                 : out   std_logic;
          line_0_13                                 : out   std_logic;
          line_0_14                                 : out   std_logic;
          line_0_15                                 : out   std_logic;
          line_0_16                                 : out   std_logic;
          line_0_17                                 : out   std_logic;
          line_0_18                                 : out   std_logic;
          line_0_19                                 : out   std_logic;
          line_0_20                                 : out   std_logic;
          line_0_21                                 : out   std_logic;
          line_0_23                                 : out   std_logic;
          line_0_24                                 : out   std_logic;
          line_0_25                                 : out   std_logic;
          line_0_26                                 : out   std_logic;
          line_0_28                                 : out   std_logic;
          line_0_29                                 : out   std_logic;
          line_0_27                                 : out   std_logic;
          line_0_30                                 : out   std_logic;
          line_4_0                                  : out   std_logic;
          line_4_1                                  : out   std_logic;
          line_4_2                                  : out   std_logic;
          line_4_3                                  : out   std_logic;
          line_4_5                                  : out   std_logic;
          line_4_6                                  : out   std_logic;
          line_4_8                                  : out   std_logic;
          line_4_9                                  : out   std_logic;
          line_4_10                                 : out   std_logic;
          line_4_13                                 : out   std_logic;
          line_4_14                                 : out   std_logic;
          line_4_15                                 : out   std_logic;
          line_4_16                                 : out   std_logic;
          line_4_17                                 : out   std_logic;
          line_4_18                                 : out   std_logic;
          line_4_19                                 : out   std_logic;
          line_4_20                                 : out   std_logic;
          line_4_21                                 : out   std_logic;
          line_4_23                                 : out   std_logic;
          line_4_24                                 : out   std_logic;
          line_4_25                                 : out   std_logic;
          line_4_26                                 : out   std_logic;
          line_4_28                                 : out   std_logic;
          line_4_29                                 : out   std_logic;
          line_1_0                                  : out   std_logic;
          line_1_1                                  : out   std_logic;
          line_1_2                                  : out   std_logic;
          line_1_3                                  : out   std_logic;
          line_1_5                                  : out   std_logic;
          line_1_6                                  : out   std_logic;
          line_1_8                                  : out   std_logic;
          line_1_9                                  : out   std_logic;
          line_1_10                                 : out   std_logic;
          line_1_13                                 : out   std_logic;
          line_1_14                                 : out   std_logic;
          line_1_15                                 : out   std_logic;
          line_1_16                                 : out   std_logic;
          line_1_17                                 : out   std_logic;
          line_1_18                                 : out   std_logic;
          line_1_19                                 : out   std_logic;
          line_1_20                                 : out   std_logic;
          line_1_21                                 : out   std_logic;
          line_1_23                                 : out   std_logic;
          line_1_24                                 : out   std_logic;
          line_1_25                                 : out   std_logic;
          line_1_26                                 : out   std_logic;
          line_1_28                                 : out   std_logic;
          line_1_29                                 : out   std_logic;
          line_1_27                                 : out   std_logic;
          line_1_30                                 : out   std_logic;
          line_5_0                                  : out   std_logic;
          line_5_1                                  : out   std_logic;
          line_5_2                                  : out   std_logic;
          line_5_3                                  : out   std_logic;
          line_5_5                                  : out   std_logic;
          line_5_6                                  : out   std_logic;
          line_5_8                                  : out   std_logic;
          line_5_9                                  : out   std_logic;
          line_5_10                                 : out   std_logic;
          line_5_13                                 : out   std_logic;
          line_5_14                                 : out   std_logic;
          line_5_15                                 : out   std_logic;
          line_5_16                                 : out   std_logic;
          line_5_17                                 : out   std_logic;
          line_5_18                                 : out   std_logic;
          line_5_19                                 : out   std_logic;
          line_5_20                                 : out   std_logic;
          line_5_21                                 : out   std_logic;
          line_5_23                                 : out   std_logic;
          line_5_24                                 : out   std_logic;
          line_5_25                                 : out   std_logic;
          line_5_26                                 : out   std_logic;
          line_5_28                                 : out   std_logic;
          line_5_29                                 : out   std_logic;
          line_6_0                                  : out   std_logic;
          line_6_1                                  : out   std_logic;
          line_6_2                                  : out   std_logic;
          line_6_3                                  : out   std_logic;
          line_6_5                                  : out   std_logic;
          line_6_6                                  : out   std_logic;
          line_6_8                                  : out   std_logic;
          line_6_9                                  : out   std_logic;
          line_6_10                                 : out   std_logic;
          line_6_13                                 : out   std_logic;
          line_6_14                                 : out   std_logic;
          line_6_15                                 : out   std_logic;
          line_6_16                                 : out   std_logic;
          line_6_17                                 : out   std_logic;
          line_6_18                                 : out   std_logic;
          line_6_19                                 : out   std_logic;
          line_6_20                                 : out   std_logic;
          line_6_21                                 : out   std_logic;
          line_6_23                                 : out   std_logic;
          line_6_24                                 : out   std_logic;
          line_6_25                                 : out   std_logic;
          line_6_26                                 : out   std_logic;
          line_6_28                                 : out   std_logic;
          line_6_29                                 : out   std_logic;
          line_2_0                                  : out   std_logic;
          line_2_1                                  : out   std_logic;
          line_2_2                                  : out   std_logic;
          line_2_3                                  : out   std_logic;
          line_2_5                                  : out   std_logic;
          line_2_6                                  : out   std_logic;
          line_2_8                                  : out   std_logic;
          line_2_9                                  : out   std_logic;
          line_2_10                                 : out   std_logic;
          line_2_13                                 : out   std_logic;
          line_2_14                                 : out   std_logic;
          line_2_15                                 : out   std_logic;
          line_2_16                                 : out   std_logic;
          line_2_17                                 : out   std_logic;
          line_2_18                                 : out   std_logic;
          line_2_19                                 : out   std_logic;
          line_2_20                                 : out   std_logic;
          line_2_21                                 : out   std_logic;
          line_2_23                                 : out   std_logic;
          line_2_24                                 : out   std_logic;
          line_2_25                                 : out   std_logic;
          line_2_26                                 : out   std_logic;
          line_2_28                                 : out   std_logic;
          line_2_29                                 : out   std_logic;
          line_2_27                                 : out   std_logic;
          line_2_30                                 : out   std_logic;
          SHA256_Module_0_do_valid_o                : out   std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F       : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0      : in    std_logic := 'U';
          N_507                                     : out   std_logic;
          N_508                                     : out   std_logic;
          ren_pos                                   : out   std_logic;
          AHB_slave_dummy_0_read_en                 : in    std_logic := 'U';
          SHA256_Module_0_error_o                   : out   std_logic;
          SHA256_Module_0_di_req_o                  : out   std_logic;
          SHA256_Module_0_waiting_data              : out   std_logic;
          SHA256_Module_0_data_available_lastbank_8 : out   std_logic;
          SHA256_Module_0_data_available            : out   std_logic;
          N_111_i_0                                 : in    std_logic := 'U';
          N_109_i_0                                 : in    std_logic := 'U';
          N_168_i_0                                 : in    std_logic := 'U';
          N_107_i_0                                 : in    std_logic := 'U';
          N_99_i_0                                  : in    std_logic := 'U';
          N_97_i_0                                  : in    std_logic := 'U';
          N_67_i_0                                  : in    std_logic := 'U';
          N_65_i_0                                  : in    std_logic := 'U';
          N_105_i_0                                 : in    std_logic := 'U';
          N_103_i_0                                 : in    std_logic := 'U';
          N_158_i_0                                 : in    std_logic := 'U';
          N_156_i_0                                 : in    std_logic := 'U';
          N_101_i_0                                 : in    std_logic := 'U';
          N_152_i_0                                 : in    std_logic := 'U';
          N_95_i_0                                  : in    std_logic := 'U';
          N_93_i_0                                  : in    std_logic := 'U';
          N_91_i_0                                  : in    std_logic := 'U';
          N_140_i_0                                 : in    std_logic := 'U';
          N_89_i_0                                  : in    std_logic := 'U';
          N_87_i_0                                  : in    std_logic := 'U';
          N_133_i_0                                 : in    std_logic := 'U';
          N_85_i_0                                  : in    std_logic := 'U';
          N_83_i_0                                  : in    std_logic := 'U';
          N_77_i_0                                  : in    std_logic := 'U';
          N_75_i_0                                  : in    std_logic := 'U';
          N_73_i_0                                  : in    std_logic := 'U';
          N_71_i_0                                  : in    std_logic := 'U';
          N_69_i_0                                  : in    std_logic := 'U';
          N_116_i_0                                 : in    std_logic := 'U';
          N_114_i_0                                 : in    std_logic := 'U';
          N_112_i_0                                 : in    std_logic := 'U';
          N_110_i_0                                 : in    std_logic := 'U';
          CertificationSystem_sb_0_GPIO_1_M2F       : in    std_logic := 'U';
          AHB_slave_dummy_0_write_en                : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CertificationSystem_sb
    port( result_addr_net_0                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          line_7                                     : in    std_logic_vector(2 downto 1) := (others => 'U');
          xhdl1222_2                                 : out   std_logic;
          line_13                                    : in    std_logic := 'U';
          line_10                                    : in    std_logic := 'U';
          line_21                                    : in    std_logic := 'U';
          line_24                                    : in    std_logic := 'U';
          line_18                                    : in    std_logic := 'U';
          line_23                                    : in    std_logic := 'U';
          line_16                                    : in    std_logic := 'U';
          line_28                                    : in    std_logic := 'U';
          line_9                                     : in    std_logic := 'U';
          line_3_d0                                  : in    std_logic := 'U';
          line_5_d0                                  : in    std_logic := 'U';
          line_15                                    : in    std_logic := 'U';
          line_26                                    : in    std_logic := 'U';
          line_14                                    : in    std_logic := 'U';
          line_20                                    : in    std_logic := 'U';
          line_2_d0                                  : in    std_logic := 'U';
          line_25                                    : in    std_logic := 'U';
          line_29                                    : in    std_logic := 'U';
          line_19                                    : in    std_logic := 'U';
          line_27                                    : in    std_logic := 'U';
          line_30                                    : in    std_logic := 'U';
          line_17                                    : in    std_logic := 'U';
          line_8                                     : in    std_logic := 'U';
          line_0_d0                                  : in    std_logic := 'U';
          line_6_d0                                  : in    std_logic := 'U';
          line_1_d0                                  : in    std_logic := 'U';
          line_0_10                                  : in    std_logic := 'U';
          line_0_21                                  : in    std_logic := 'U';
          line_0_24                                  : in    std_logic := 'U';
          line_0_18                                  : in    std_logic := 'U';
          line_0_23                                  : in    std_logic := 'U';
          line_0_16                                  : in    std_logic := 'U';
          line_0_28                                  : in    std_logic := 'U';
          line_0_9                                   : in    std_logic := 'U';
          line_0_3                                   : in    std_logic := 'U';
          line_0_5                                   : in    std_logic := 'U';
          line_0_15                                  : in    std_logic := 'U';
          line_0_26                                  : in    std_logic := 'U';
          line_0_14                                  : in    std_logic := 'U';
          line_0_20                                  : in    std_logic := 'U';
          line_0_2                                   : in    std_logic := 'U';
          line_0_25                                  : in    std_logic := 'U';
          line_0_29                                  : in    std_logic := 'U';
          line_0_19                                  : in    std_logic := 'U';
          line_0_27                                  : in    std_logic := 'U';
          line_0_30                                  : in    std_logic := 'U';
          line_0_17                                  : in    std_logic := 'U';
          line_0_8                                   : in    std_logic := 'U';
          line_0_0                                   : in    std_logic := 'U';
          line_0_1                                   : in    std_logic := 'U';
          line_0_6                                   : in    std_logic := 'U';
          line_0_13                                  : in    std_logic := 'U';
          line_1_10                                  : in    std_logic := 'U';
          line_1_21                                  : in    std_logic := 'U';
          line_1_24                                  : in    std_logic := 'U';
          line_1_18                                  : in    std_logic := 'U';
          line_1_23                                  : in    std_logic := 'U';
          line_1_16                                  : in    std_logic := 'U';
          line_1_28                                  : in    std_logic := 'U';
          line_1_9                                   : in    std_logic := 'U';
          line_1_3                                   : in    std_logic := 'U';
          line_1_5                                   : in    std_logic := 'U';
          line_1_15                                  : in    std_logic := 'U';
          line_1_26                                  : in    std_logic := 'U';
          line_1_14                                  : in    std_logic := 'U';
          line_1_20                                  : in    std_logic := 'U';
          line_1_2                                   : in    std_logic := 'U';
          line_1_25                                  : in    std_logic := 'U';
          line_1_29                                  : in    std_logic := 'U';
          line_1_19                                  : in    std_logic := 'U';
          line_1_27                                  : in    std_logic := 'U';
          line_1_30                                  : in    std_logic := 'U';
          line_1_17                                  : in    std_logic := 'U';
          line_1_8                                   : in    std_logic := 'U';
          line_1_0                                   : in    std_logic := 'U';
          line_1_1                                   : in    std_logic := 'U';
          line_1_6                                   : in    std_logic := 'U';
          line_1_13                                  : in    std_logic := 'U';
          line_2_19                                  : in    std_logic := 'U';
          line_2_27                                  : in    std_logic := 'U';
          line_2_30                                  : in    std_logic := 'U';
          line_2_17                                  : in    std_logic := 'U';
          line_2_8                                   : in    std_logic := 'U';
          line_2_10                                  : in    std_logic := 'U';
          line_2_15                                  : in    std_logic := 'U';
          line_2_26                                  : in    std_logic := 'U';
          line_2_20                                  : in    std_logic := 'U';
          line_2_0                                   : in    std_logic := 'U';
          line_2_1                                   : in    std_logic := 'U';
          line_2_29                                  : in    std_logic := 'U';
          line_2_25                                  : in    std_logic := 'U';
          line_2_2                                   : in    std_logic := 'U';
          line_2_6                                   : in    std_logic := 'U';
          line_2_13                                  : in    std_logic := 'U';
          line_2_14                                  : in    std_logic := 'U';
          line_2_5                                   : in    std_logic := 'U';
          line_2_3                                   : in    std_logic := 'U';
          line_2_9                                   : in    std_logic := 'U';
          line_2_28                                  : in    std_logic := 'U';
          line_2_16                                  : in    std_logic := 'U';
          line_2_23                                  : in    std_logic := 'U';
          line_2_18                                  : in    std_logic := 'U';
          line_2_24                                  : in    std_logic := 'U';
          line_2_21                                  : in    std_logic := 'U';
          line_3_19                                  : in    std_logic := 'U';
          line_3_17                                  : in    std_logic := 'U';
          line_3_8                                   : in    std_logic := 'U';
          line_3_0                                   : in    std_logic := 'U';
          line_3_1                                   : in    std_logic := 'U';
          line_3_29                                  : in    std_logic := 'U';
          line_3_25                                  : in    std_logic := 'U';
          line_3_2                                   : in    std_logic := 'U';
          line_3_20                                  : in    std_logic := 'U';
          line_3_6                                   : in    std_logic := 'U';
          line_3_13                                  : in    std_logic := 'U';
          line_3_14                                  : in    std_logic := 'U';
          line_3_26                                  : in    std_logic := 'U';
          line_3_15                                  : in    std_logic := 'U';
          line_3_5                                   : in    std_logic := 'U';
          line_3_3                                   : in    std_logic := 'U';
          line_3_9                                   : in    std_logic := 'U';
          line_3_28                                  : in    std_logic := 'U';
          line_3_16                                  : in    std_logic := 'U';
          line_3_23                                  : in    std_logic := 'U';
          line_3_18                                  : in    std_logic := 'U';
          line_3_24                                  : in    std_logic := 'U';
          line_3_21                                  : in    std_logic := 'U';
          line_3_10                                  : in    std_logic := 'U';
          SHA256_Module_0_data_out_5                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_13                : in    std_logic := 'U';
          SHA256_Module_0_data_out_12                : in    std_logic := 'U';
          SHA256_Module_0_data_out_8                 : in    std_logic := 'U';
          SHA256_Module_0_data_out_23                : in    std_logic := 'U';
          SHA256_Module_0_data_out_0                 : in    std_logic := 'U';
          line_4_19                                  : in    std_logic := 'U';
          line_4_17                                  : in    std_logic := 'U';
          line_4_8                                   : in    std_logic := 'U';
          line_4_0                                   : in    std_logic := 'U';
          line_4_1                                   : in    std_logic := 'U';
          line_4_29                                  : in    std_logic := 'U';
          line_4_25                                  : in    std_logic := 'U';
          line_4_2                                   : in    std_logic := 'U';
          line_4_20                                  : in    std_logic := 'U';
          line_4_14                                  : in    std_logic := 'U';
          line_4_26                                  : in    std_logic := 'U';
          line_4_15                                  : in    std_logic := 'U';
          line_4_5                                   : in    std_logic := 'U';
          line_4_3                                   : in    std_logic := 'U';
          line_4_9                                   : in    std_logic := 'U';
          line_4_28                                  : in    std_logic := 'U';
          line_4_16                                  : in    std_logic := 'U';
          line_4_23                                  : in    std_logic := 'U';
          line_4_18                                  : in    std_logic := 'U';
          line_4_24                                  : in    std_logic := 'U';
          line_4_21                                  : in    std_logic := 'U';
          line_4_10                                  : in    std_logic := 'U';
          line_4_6                                   : in    std_logic := 'U';
          line_4_13                                  : in    std_logic := 'U';
          line_5_19                                  : in    std_logic := 'U';
          line_5_17                                  : in    std_logic := 'U';
          line_5_8                                   : in    std_logic := 'U';
          line_5_0                                   : in    std_logic := 'U';
          line_5_1                                   : in    std_logic := 'U';
          line_5_29                                  : in    std_logic := 'U';
          line_5_25                                  : in    std_logic := 'U';
          line_5_2                                   : in    std_logic := 'U';
          line_5_20                                  : in    std_logic := 'U';
          line_5_6                                   : in    std_logic := 'U';
          line_5_13                                  : in    std_logic := 'U';
          line_5_14                                  : in    std_logic := 'U';
          line_5_26                                  : in    std_logic := 'U';
          line_5_15                                  : in    std_logic := 'U';
          line_5_5                                   : in    std_logic := 'U';
          line_5_3                                   : in    std_logic := 'U';
          line_5_9                                   : in    std_logic := 'U';
          line_5_28                                  : in    std_logic := 'U';
          line_5_16                                  : in    std_logic := 'U';
          line_5_23                                  : in    std_logic := 'U';
          line_5_18                                  : in    std_logic := 'U';
          line_5_24                                  : in    std_logic := 'U';
          line_5_21                                  : in    std_logic := 'U';
          line_5_10                                  : in    std_logic := 'U';
          line_6_19                                  : in    std_logic := 'U';
          line_6_17                                  : in    std_logic := 'U';
          line_6_8                                   : in    std_logic := 'U';
          line_6_0                                   : in    std_logic := 'U';
          line_6_1                                   : in    std_logic := 'U';
          line_6_29                                  : in    std_logic := 'U';
          line_6_25                                  : in    std_logic := 'U';
          line_6_2                                   : in    std_logic := 'U';
          line_6_20                                  : in    std_logic := 'U';
          line_6_6                                   : in    std_logic := 'U';
          line_6_13                                  : in    std_logic := 'U';
          line_6_14                                  : in    std_logic := 'U';
          line_6_26                                  : in    std_logic := 'U';
          line_6_15                                  : in    std_logic := 'U';
          line_6_5                                   : in    std_logic := 'U';
          line_6_3                                   : in    std_logic := 'U';
          line_6_9                                   : in    std_logic := 'U';
          line_6_28                                  : in    std_logic := 'U';
          line_6_16                                  : in    std_logic := 'U';
          line_6_23                                  : in    std_logic := 'U';
          line_6_18                                  : in    std_logic := 'U';
          line_6_24                                  : in    std_logic := 'U';
          line_6_21                                  : in    std_logic := 'U';
          line_6_10                                  : in    std_logic := 'U';
          CertificationSystem_sb_0_POWER_ON_RESET_N  : out   std_logic;
          DEVRST_N                                   : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0       : out   std_logic;
          SPI_0_SS0                                  : inout   std_logic;
          SPI_0_DO                                   : out   std_logic;
          SPI_0_DI                                   : in    std_logic := 'U';
          SPI_0_CLK                                  : inout   std_logic;
          MMUART_1_TXD                               : out   std_logic;
          MMUART_1_RXD                               : in    std_logic := 'U';
          CertificationSystem_sb_0_GPIO_1_M2F        : out   std_logic;
          GPIO_0_M2F_c                               : out   std_logic;
          CertificationSystem_sb_0_GPIO_9_M2F        : out   std_logic;
          SHA256_Module_0_waiting_data               : in    std_logic := 'U';
          SHA256_Module_0_data_available_lastbank_8  : in    std_logic := 'U';
          SHA256_Module_0_di_req_o                   : in    std_logic := 'U';
          SHA256_Module_0_do_valid_o                 : in    std_logic := 'U';
          SHA256_Module_0_data_available             : in    std_logic := 'U';
          SHA256_Module_0_error_o                    : in    std_logic := 'U';
          CertificationSystem_sb_0_AHBmslave5_HREADY : in    std_logic := 'U';
          N_225                                      : out   std_logic;
          N_276                                      : out   std_logic;
          N_259                                      : out   std_logic;
          N_277                                      : out   std_logic;
          ren_pos                                    : in    std_logic := 'U';
          N_206                                      : out   std_logic;
          N_508                                      : in    std_logic := 'U';
          N_507                                      : in    std_logic := 'U';
          un8_hreadyin_i_0                           : out   std_logic;
          N_226                                      : out   std_logic;
          N_65_i_0                                   : out   std_logic;
          N_67_i_0                                   : out   std_logic;
          N_110_i_0                                  : out   std_logic;
          N_112_i_0                                  : out   std_logic;
          N_114_i_0                                  : out   std_logic;
          N_116_i_0                                  : out   std_logic;
          N_69_i_0                                   : out   std_logic;
          N_71_i_0                                   : out   std_logic;
          N_73_i_0                                   : out   std_logic;
          N_75_i_0                                   : out   std_logic;
          N_77_i_0                                   : out   std_logic;
          N_83_i_0                                   : out   std_logic;
          N_85_i_0                                   : out   std_logic;
          N_133_i_0                                  : out   std_logic;
          N_87_i_0                                   : out   std_logic;
          N_89_i_0                                   : out   std_logic;
          N_140_i_0                                  : out   std_logic;
          N_91_i_0                                   : out   std_logic;
          N_93_i_0                                   : out   std_logic;
          N_95_i_0                                   : out   std_logic;
          N_97_i_0                                   : out   std_logic;
          N_99_i_0                                   : out   std_logic;
          N_152_i_0                                  : out   std_logic;
          N_101_i_0                                  : out   std_logic;
          N_156_i_0                                  : out   std_logic;
          N_158_i_0                                  : out   std_logic;
          N_103_i_0                                  : out   std_logic;
          N_105_i_0                                  : out   std_logic;
          N_107_i_0                                  : out   std_logic;
          N_168_i_0                                  : out   std_logic;
          N_109_i_0                                  : out   std_logic;
          N_111_i_0                                  : out   std_logic;
          N_218_i_0                                  : out   std_logic;
          N_217_i_0                                  : out   std_logic;
          N_203_i_0                                  : out   std_logic
        );
  end component;

  component AHB_slave_dummy
    port( waddr_in_net_0                             : out   std_logic_vector(4 downto 0);
          result_addr_net_0                          : out   std_logic_vector(3 downto 0);
          xhdl1222                                   : in    std_logic_vector(5 to 5) := (others => 'U');
          CertificationSystem_sb_0_POWER_ON_RESET_N  : in    std_logic := 'U';
          CertificationSystem_sb_0_FAB_CCC_GL0       : in    std_logic := 'U';
          N_276                                      : in    std_logic := 'U';
          N_203_i_0                                  : in    std_logic := 'U';
          N_217_i_0                                  : in    std_logic := 'U';
          N_218_i_0                                  : in    std_logic := 'U';
          N_259                                      : in    std_logic := 'U';
          CertificationSystem_sb_0_AHBmslave5_HREADY : out   std_logic;
          AHB_slave_dummy_0_write_en                 : out   std_logic;
          AHB_slave_dummy_0_read_en                  : out   std_logic;
          N_277                                      : in    std_logic := 'U';
          N_225                                      : in    std_logic := 'U';
          N_206                                      : in    std_logic := 'U';
          un8_hreadyin_i_0                           : in    std_logic := 'U';
          N_226                                      : in    std_logic := 'U'
        );
  end component;

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

    signal CertificationSystem_sb_0_FAB_CCC_GL0, 
        CertificationSystem_sb_0_POWER_ON_RESET_N, 
        CertificationSystem_sb_0_AHBmslave5_HREADY, 
        \waddr_in_net_0[0]\, \waddr_in_net_0[1]\, 
        \waddr_in_net_0[2]\, \waddr_in_net_0[3]\, 
        \waddr_in_net_0[4]\, \result_addr_net_0[0]\, 
        \result_addr_net_0[1]\, \result_addr_net_0[2]\, 
        \result_addr_net_0[3]\, AHB_slave_dummy_0_write_en, 
        AHB_slave_dummy_0_read_en, VCC_net_1, 
        SHA256_Module_0_waiting_data, 
        SHA256_Module_0_data_available_lastbank_8, 
        SHA256_Module_0_di_req_o, GND_net_1, 
        SHA256_Module_0_do_valid_o, 
        SHA256_Module_0_data_available, SHA256_Module_0_error_o, 
        CertificationSystem_sb_0_GPIO_1_M2F, 
        CertificationSystem_sb_0_GPIO_9_M2F, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[1]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[2]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[1]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[2]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[3]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[4]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[6]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[9]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[14]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[15]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[16]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[17]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[18]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[19]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[21]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[22]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[24]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[25]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[26]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[27]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[29]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[30]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[1]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[2]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[3]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[4]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[6]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[9]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[14]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[15]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[16]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[17]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[18]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[19]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[21]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[22]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[24]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[25]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[26]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[27]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[29]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[30]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[1]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[2]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[3]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[4]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[6]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[9]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[14]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[15]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[16]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[17]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[18]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[19]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[21]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[22]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[24]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[25]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[26]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[27]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[29]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[30]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[1]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[2]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[3]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[4]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[6]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[9]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[14]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[15]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[16]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[17]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[18]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[19]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[21]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[22]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[24]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[25]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[26]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[27]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[29]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[30]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[1]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[2]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[3]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[4]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[6]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[9]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[14]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[15]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[16]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[17]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[18]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[19]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[21]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[22]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[24]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[25]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[26]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[27]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[29]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[30]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[1]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[2]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[3]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[4]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[6]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[9]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[14]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[15]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[16]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[17]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[18]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[19]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[21]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[22]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[24]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[25]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[26]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[27]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[29]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[30]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[1]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[2]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[3]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[4]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[6]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[9]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[14]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[15]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[16]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[17]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[18]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[19]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[21]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[22]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[24]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[25]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[26]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[27]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[28]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[29]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[30]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[31]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.ren_pos\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[1]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[2]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[3]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[4]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[6]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[7]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[9]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[10]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[11]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[14]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[15]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[16]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[17]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[18]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[19]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[20]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[21]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[22]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[24]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[25]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[26]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[27]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[29]\, 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[30]\, 
        \CertificationSystem_sb_0.CoreAHBLite_0.matrix4x16.xhdl1222[5]\, 
        N_226, GPIO_0_M2F_c, N_276, N_259, N_277, 
        \SHA256_Module_0_data_out[8]\, N_206, N_225, 
        \SHA256_Module_0_data_out[23]\, 
        \SHA256_Module_0_data_out[0]\, 
        \SHA256_Module_0_data_out[12]\, N_508, 
        \SHA256_Module_0_data_out[13]\, 
        \SHA256_Module_0_data_out[5]\, N_507, 
        \CertificationSystem_sb_0.COREAHBLSRAM_0_0.U_CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf.un8_hreadyin_i_0\, 
        N_65_i_0, N_67_i_0, N_110_i_0, N_112_i_0, N_114_i_0, 
        N_116_i_0, N_69_i_0, N_71_i_0, N_73_i_0, N_75_i_0, 
        N_77_i_0, N_83_i_0, N_85_i_0, N_133_i_0, N_87_i_0, 
        N_89_i_0, N_140_i_0, N_91_i_0, N_93_i_0, N_95_i_0, 
        N_97_i_0, N_99_i_0, N_152_i_0, N_101_i_0, N_156_i_0, 
        N_158_i_0, N_103_i_0, N_105_i_0, N_107_i_0, N_168_i_0, 
        N_109_i_0, N_111_i_0, N_218_i_0, N_217_i_0, N_203_i_0
         : std_logic;

    for all : SHA256_Module
	Use entity work.SHA256_Module(DEF_ARCH);
    for all : CertificationSystem_sb
	Use entity work.CertificationSystem_sb(DEF_ARCH);
    for all : AHB_slave_dummy
	Use entity work.AHB_slave_dummy(DEF_ARCH);
begin 


    SHA256_Module_0 : SHA256_Module
      port map(result_addr_net_0(3) => \result_addr_net_0[3]\, 
        result_addr_net_0(2) => \result_addr_net_0[2]\, 
        result_addr_net_0(1) => \result_addr_net_0[1]\, 
        result_addr_net_0(0) => \result_addr_net_0[0]\, line_7(2)
         => \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[2]\, 
        line_7(1) => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[1]\, 
        waddr_in_net_0(4) => \waddr_in_net_0[4]\, 
        waddr_in_net_0(3) => \waddr_in_net_0[3]\, 
        waddr_in_net_0(2) => \waddr_in_net_0[2]\, 
        waddr_in_net_0(1) => \waddr_in_net_0[1]\, 
        waddr_in_net_0(0) => \waddr_in_net_0[0]\, 
        SHA256_Module_0_data_out_5 => 
        \SHA256_Module_0_data_out[5]\, 
        SHA256_Module_0_data_out_13 => 
        \SHA256_Module_0_data_out[13]\, 
        SHA256_Module_0_data_out_12 => 
        \SHA256_Module_0_data_out[12]\, 
        SHA256_Module_0_data_out_23 => 
        \SHA256_Module_0_data_out[23]\, 
        SHA256_Module_0_data_out_8 => 
        \SHA256_Module_0_data_out[8]\, SHA256_Module_0_data_out_0
         => \SHA256_Module_0_data_out[0]\, line_0_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[1]\, 
        line_1_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[2]\, 
        line_2_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[3]\, 
        line_3_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[4]\, 
        line_5_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[6]\, 
        line_6_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[7]\, line_8
         => \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[9]\, 
        line_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[10]\, 
        line_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[11]\, 
        line_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[14]\, 
        line_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[15]\, 
        line_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[16]\, 
        line_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[17]\, 
        line_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[18]\, 
        line_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[19]\, 
        line_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[20]\, 
        line_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[21]\, 
        line_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[22]\, 
        line_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[24]\, 
        line_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[25]\, 
        line_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[26]\, 
        line_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[27]\, 
        line_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[29]\, 
        line_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[30]\, 
        line_27 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[28]\, 
        line_30 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[31]\, 
        line_3_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[1]\, 
        line_3_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[2]\, 
        line_3_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[3]\, 
        line_3_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[4]\, 
        line_3_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[6]\, 
        line_3_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[7]\, 
        line_3_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[9]\, 
        line_3_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[10]\, 
        line_3_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[11]\, 
        line_3_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[14]\, 
        line_3_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[15]\, 
        line_3_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[16]\, 
        line_3_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[17]\, 
        line_3_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[18]\, 
        line_3_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[19]\, 
        line_3_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[20]\, 
        line_3_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[21]\, 
        line_3_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[22]\, 
        line_3_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[24]\, 
        line_3_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[25]\, 
        line_3_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[26]\, 
        line_3_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[27]\, 
        line_3_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[29]\, 
        line_3_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[30]\, 
        line_0_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[1]\, 
        line_0_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[2]\, 
        line_0_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[3]\, 
        line_0_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[4]\, 
        line_0_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[6]\, 
        line_0_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[7]\, 
        line_0_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[9]\, 
        line_0_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[10]\, 
        line_0_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[11]\, 
        line_0_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[14]\, 
        line_0_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[15]\, 
        line_0_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[16]\, 
        line_0_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[17]\, 
        line_0_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[18]\, 
        line_0_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[19]\, 
        line_0_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[20]\, 
        line_0_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[21]\, 
        line_0_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[22]\, 
        line_0_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[24]\, 
        line_0_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[25]\, 
        line_0_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[26]\, 
        line_0_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[27]\, 
        line_0_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[29]\, 
        line_0_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[30]\, 
        line_0_27 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[28]\, 
        line_0_30 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[31]\, 
        line_4_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[1]\, 
        line_4_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[2]\, 
        line_4_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[3]\, 
        line_4_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[4]\, 
        line_4_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[6]\, 
        line_4_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[7]\, 
        line_4_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[9]\, 
        line_4_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[10]\, 
        line_4_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[11]\, 
        line_4_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[14]\, 
        line_4_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[15]\, 
        line_4_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[16]\, 
        line_4_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[17]\, 
        line_4_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[18]\, 
        line_4_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[19]\, 
        line_4_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[20]\, 
        line_4_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[21]\, 
        line_4_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[22]\, 
        line_4_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[24]\, 
        line_4_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[25]\, 
        line_4_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[26]\, 
        line_4_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[27]\, 
        line_4_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[29]\, 
        line_4_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[30]\, 
        line_1_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[1]\, 
        line_1_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[2]\, 
        line_1_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[3]\, 
        line_1_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[4]\, 
        line_1_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[6]\, 
        line_1_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[7]\, 
        line_1_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[9]\, 
        line_1_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[10]\, 
        line_1_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[11]\, 
        line_1_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[14]\, 
        line_1_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[15]\, 
        line_1_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[16]\, 
        line_1_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[17]\, 
        line_1_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[18]\, 
        line_1_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[19]\, 
        line_1_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[20]\, 
        line_1_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[21]\, 
        line_1_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[22]\, 
        line_1_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[24]\, 
        line_1_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[25]\, 
        line_1_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[26]\, 
        line_1_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[27]\, 
        line_1_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[29]\, 
        line_1_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[30]\, 
        line_1_27 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[28]\, 
        line_1_30 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[31]\, 
        line_5_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[1]\, 
        line_5_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[2]\, 
        line_5_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[3]\, 
        line_5_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[4]\, 
        line_5_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[6]\, 
        line_5_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[7]\, 
        line_5_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[9]\, 
        line_5_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[10]\, 
        line_5_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[11]\, 
        line_5_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[14]\, 
        line_5_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[15]\, 
        line_5_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[16]\, 
        line_5_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[17]\, 
        line_5_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[18]\, 
        line_5_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[19]\, 
        line_5_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[20]\, 
        line_5_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[21]\, 
        line_5_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[22]\, 
        line_5_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[24]\, 
        line_5_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[25]\, 
        line_5_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[26]\, 
        line_5_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[27]\, 
        line_5_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[29]\, 
        line_5_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[30]\, 
        line_6_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[1]\, 
        line_6_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[2]\, 
        line_6_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[3]\, 
        line_6_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[4]\, 
        line_6_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[6]\, 
        line_6_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[7]\, 
        line_6_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[9]\, 
        line_6_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[10]\, 
        line_6_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[11]\, 
        line_6_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[14]\, 
        line_6_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[15]\, 
        line_6_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[16]\, 
        line_6_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[17]\, 
        line_6_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[18]\, 
        line_6_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[19]\, 
        line_6_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[20]\, 
        line_6_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[21]\, 
        line_6_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[22]\, 
        line_6_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[24]\, 
        line_6_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[25]\, 
        line_6_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[26]\, 
        line_6_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[27]\, 
        line_6_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[29]\, 
        line_6_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[30]\, 
        line_2_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[1]\, 
        line_2_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[2]\, 
        line_2_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[3]\, 
        line_2_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[4]\, 
        line_2_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[6]\, 
        line_2_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[7]\, 
        line_2_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[9]\, 
        line_2_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[10]\, 
        line_2_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[11]\, 
        line_2_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[14]\, 
        line_2_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[15]\, 
        line_2_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[16]\, 
        line_2_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[17]\, 
        line_2_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[18]\, 
        line_2_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[19]\, 
        line_2_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[20]\, 
        line_2_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[21]\, 
        line_2_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[22]\, 
        line_2_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[24]\, 
        line_2_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[25]\, 
        line_2_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[26]\, 
        line_2_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[27]\, 
        line_2_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[29]\, 
        line_2_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[30]\, 
        line_2_27 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[28]\, 
        line_2_30 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[31]\, 
        SHA256_Module_0_do_valid_o => SHA256_Module_0_do_valid_o, 
        CertificationSystem_sb_0_GPIO_9_M2F => 
        CertificationSystem_sb_0_GPIO_9_M2F, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, N_507 => N_507, 
        N_508 => N_508, ren_pos => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.ren_pos\, 
        AHB_slave_dummy_0_read_en => AHB_slave_dummy_0_read_en, 
        SHA256_Module_0_error_o => SHA256_Module_0_error_o, 
        SHA256_Module_0_di_req_o => SHA256_Module_0_di_req_o, 
        SHA256_Module_0_waiting_data => 
        SHA256_Module_0_waiting_data, 
        SHA256_Module_0_data_available_lastbank_8 => 
        SHA256_Module_0_data_available_lastbank_8, 
        SHA256_Module_0_data_available => 
        SHA256_Module_0_data_available, N_111_i_0 => N_111_i_0, 
        N_109_i_0 => N_109_i_0, N_168_i_0 => N_168_i_0, N_107_i_0
         => N_107_i_0, N_99_i_0 => N_99_i_0, N_97_i_0 => N_97_i_0, 
        N_67_i_0 => N_67_i_0, N_65_i_0 => N_65_i_0, N_105_i_0 => 
        N_105_i_0, N_103_i_0 => N_103_i_0, N_158_i_0 => N_158_i_0, 
        N_156_i_0 => N_156_i_0, N_101_i_0 => N_101_i_0, N_152_i_0
         => N_152_i_0, N_95_i_0 => N_95_i_0, N_93_i_0 => N_93_i_0, 
        N_91_i_0 => N_91_i_0, N_140_i_0 => N_140_i_0, N_89_i_0
         => N_89_i_0, N_87_i_0 => N_87_i_0, N_133_i_0 => 
        N_133_i_0, N_85_i_0 => N_85_i_0, N_83_i_0 => N_83_i_0, 
        N_77_i_0 => N_77_i_0, N_75_i_0 => N_75_i_0, N_73_i_0 => 
        N_73_i_0, N_71_i_0 => N_71_i_0, N_69_i_0 => N_69_i_0, 
        N_116_i_0 => N_116_i_0, N_114_i_0 => N_114_i_0, N_112_i_0
         => N_112_i_0, N_110_i_0 => N_110_i_0, 
        CertificationSystem_sb_0_GPIO_1_M2F => 
        CertificationSystem_sb_0_GPIO_1_M2F, 
        AHB_slave_dummy_0_write_en => AHB_slave_dummy_0_write_en);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    CertificationSystem_sb_0 : CertificationSystem_sb
      port map(result_addr_net_0(3) => \result_addr_net_0[3]\, 
        result_addr_net_0(2) => \result_addr_net_0[2]\, 
        result_addr_net_0(1) => \result_addr_net_0[1]\, 
        result_addr_net_0(0) => \result_addr_net_0[0]\, line_7(2)
         => \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[2]\, 
        line_7(1) => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[1]\, 
        xhdl1222_2 => 
        \CertificationSystem_sb_0.CoreAHBLite_0.matrix4x16.xhdl1222[5]\, 
        line_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[14]\, 
        line_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[11]\, 
        line_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[22]\, 
        line_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[25]\, 
        line_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[19]\, 
        line_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[24]\, 
        line_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[17]\, 
        line_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[29]\, line_9
         => \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[10]\, 
        line_3_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[4]\, 
        line_5_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[6]\, line_15
         => \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[16]\, 
        line_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[27]\, 
        line_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[15]\, 
        line_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[21]\, 
        line_2_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[3]\, line_25
         => \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[26]\, 
        line_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[30]\, 
        line_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[20]\, 
        line_27 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[28]\, 
        line_30 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[31]\, 
        line_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[18]\, line_8
         => \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[9]\, 
        line_0_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[1]\, 
        line_6_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[7]\, 
        line_1_d0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[2]\, 
        line_0_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[11]\, 
        line_0_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[22]\, 
        line_0_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[25]\, 
        line_0_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[19]\, 
        line_0_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[24]\, 
        line_0_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[17]\, 
        line_0_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[29]\, 
        line_0_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[10]\, 
        line_0_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[4]\, 
        line_0_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[6]\, 
        line_0_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[16]\, 
        line_0_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[27]\, 
        line_0_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[15]\, 
        line_0_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[21]\, 
        line_0_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[3]\, 
        line_0_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[26]\, 
        line_0_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[30]\, 
        line_0_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[20]\, 
        line_0_27 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[28]\, 
        line_0_30 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[31]\, 
        line_0_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[18]\, 
        line_0_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[9]\, 
        line_0_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[1]\, 
        line_0_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[2]\, 
        line_0_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[7]\, 
        line_0_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[14]\, 
        line_1_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[11]\, 
        line_1_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[22]\, 
        line_1_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[25]\, 
        line_1_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[19]\, 
        line_1_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[24]\, 
        line_1_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[17]\, 
        line_1_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[29]\, 
        line_1_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[10]\, 
        line_1_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[4]\, 
        line_1_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[6]\, 
        line_1_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[16]\, 
        line_1_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[27]\, 
        line_1_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[15]\, 
        line_1_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[21]\, 
        line_1_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[3]\, 
        line_1_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[26]\, 
        line_1_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[30]\, 
        line_1_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[20]\, 
        line_1_27 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[28]\, 
        line_1_30 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[31]\, 
        line_1_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[18]\, 
        line_1_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[9]\, 
        line_1_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[1]\, 
        line_1_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[2]\, 
        line_1_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[7]\, 
        line_1_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[14]\, 
        line_2_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[20]\, 
        line_2_27 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[28]\, 
        line_2_30 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[31]\, 
        line_2_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[18]\, 
        line_2_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[9]\, 
        line_2_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[11]\, 
        line_2_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[16]\, 
        line_2_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[27]\, 
        line_2_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[21]\, 
        line_2_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[1]\, 
        line_2_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[2]\, 
        line_2_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[30]\, 
        line_2_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[26]\, 
        line_2_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[3]\, 
        line_2_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[7]\, 
        line_2_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[14]\, 
        line_2_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[15]\, 
        line_2_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[6]\, 
        line_2_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[4]\, 
        line_2_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[10]\, 
        line_2_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[29]\, 
        line_2_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[17]\, 
        line_2_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[24]\, 
        line_2_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[19]\, 
        line_2_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[25]\, 
        line_2_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[22]\, 
        line_3_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[20]\, 
        line_3_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[18]\, 
        line_3_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[9]\, 
        line_3_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[1]\, 
        line_3_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[2]\, 
        line_3_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[30]\, 
        line_3_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[26]\, 
        line_3_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[3]\, 
        line_3_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[21]\, 
        line_3_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[7]\, 
        line_3_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[14]\, 
        line_3_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[15]\, 
        line_3_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[27]\, 
        line_3_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[16]\, 
        line_3_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[6]\, 
        line_3_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[4]\, 
        line_3_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[10]\, 
        line_3_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[29]\, 
        line_3_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[17]\, 
        line_3_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[24]\, 
        line_3_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[19]\, 
        line_3_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[25]\, 
        line_3_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[22]\, 
        line_3_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[11]\, 
        SHA256_Module_0_data_out_5 => 
        \SHA256_Module_0_data_out[5]\, 
        SHA256_Module_0_data_out_13 => 
        \SHA256_Module_0_data_out[13]\, 
        SHA256_Module_0_data_out_12 => 
        \SHA256_Module_0_data_out[12]\, 
        SHA256_Module_0_data_out_8 => 
        \SHA256_Module_0_data_out[8]\, 
        SHA256_Module_0_data_out_23 => 
        \SHA256_Module_0_data_out[23]\, 
        SHA256_Module_0_data_out_0 => 
        \SHA256_Module_0_data_out[0]\, line_4_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[20]\, 
        line_4_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_2.line[18]\, 
        line_4_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_3.line[9]\, 
        line_4_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[1]\, 
        line_4_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.line[2]\, 
        line_4_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[30]\, 
        line_4_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[26]\, 
        line_4_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[3]\, 
        line_4_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[21]\, 
        line_4_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[15]\, 
        line_4_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[27]\, 
        line_4_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[16]\, 
        line_4_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[6]\, 
        line_4_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[4]\, 
        line_4_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[10]\, 
        line_4_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[29]\, 
        line_4_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[17]\, 
        line_4_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[24]\, 
        line_4_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[19]\, 
        line_4_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[25]\, 
        line_4_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_7.line[22]\, 
        line_4_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[11]\, 
        line_4_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[7]\, 
        line_4_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[14]\, 
        line_5_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[20]\, 
        line_5_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[18]\, 
        line_5_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_1.line[9]\, 
        line_5_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[1]\, 
        line_5_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[2]\, 
        line_5_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[30]\, 
        line_5_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[26]\, 
        line_5_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[3]\, 
        line_5_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[21]\, 
        line_5_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[7]\, 
        line_5_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[14]\, 
        line_5_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[15]\, 
        line_5_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[27]\, 
        line_5_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[16]\, 
        line_5_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[6]\, 
        line_5_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[4]\, 
        line_5_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[10]\, 
        line_5_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[29]\, 
        line_5_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[17]\, 
        line_5_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[24]\, 
        line_5_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[19]\, 
        line_5_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[25]\, 
        line_5_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[22]\, 
        line_5_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_6.line[11]\, 
        line_6_19 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[20]\, 
        line_6_17 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[18]\, 
        line_6_8 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_5.line[9]\, 
        line_6_0 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[1]\, 
        line_6_1 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[2]\, 
        line_6_29 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[30]\, 
        line_6_25 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[26]\, 
        line_6_2 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[3]\, 
        line_6_20 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[21]\, 
        line_6_6 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[7]\, 
        line_6_13 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_0.line[14]\, 
        line_6_14 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[15]\, 
        line_6_26 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[27]\, 
        line_6_15 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[16]\, 
        line_6_5 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[6]\, 
        line_6_3 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[4]\, 
        line_6_9 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[10]\, 
        line_6_28 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[29]\, 
        line_6_16 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[17]\, 
        line_6_23 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[24]\, 
        line_6_18 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[19]\, 
        line_6_24 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[25]\, 
        line_6_21 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[22]\, 
        line_6_10 => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_4.line[11]\, 
        CertificationSystem_sb_0_POWER_ON_RESET_N => 
        CertificationSystem_sb_0_POWER_ON_RESET_N, DEVRST_N => 
        DEVRST_N, CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, SPI_0_SS0 => 
        SPI_0_SS0, SPI_0_DO => SPI_0_DO, SPI_0_DI => SPI_0_DI, 
        SPI_0_CLK => SPI_0_CLK, MMUART_1_TXD => MMUART_1_TXD, 
        MMUART_1_RXD => MMUART_1_RXD, 
        CertificationSystem_sb_0_GPIO_1_M2F => 
        CertificationSystem_sb_0_GPIO_1_M2F, GPIO_0_M2F_c => 
        GPIO_0_M2F_c, CertificationSystem_sb_0_GPIO_9_M2F => 
        CertificationSystem_sb_0_GPIO_9_M2F, 
        SHA256_Module_0_waiting_data => 
        SHA256_Module_0_waiting_data, 
        SHA256_Module_0_data_available_lastbank_8 => 
        SHA256_Module_0_data_available_lastbank_8, 
        SHA256_Module_0_di_req_o => SHA256_Module_0_di_req_o, 
        SHA256_Module_0_do_valid_o => SHA256_Module_0_do_valid_o, 
        SHA256_Module_0_data_available => 
        SHA256_Module_0_data_available, SHA256_Module_0_error_o
         => SHA256_Module_0_error_o, 
        CertificationSystem_sb_0_AHBmslave5_HREADY => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, N_225 => 
        N_225, N_276 => N_276, N_259 => N_259, N_277 => N_277, 
        ren_pos => 
        \SHA256_Module_0.reg9_1x32_0.reg_1x32_8.ren_pos\, N_206
         => N_206, N_508 => N_508, N_507 => N_507, 
        un8_hreadyin_i_0 => 
        \CertificationSystem_sb_0.COREAHBLSRAM_0_0.U_CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf.un8_hreadyin_i_0\, 
        N_226 => N_226, N_65_i_0 => N_65_i_0, N_67_i_0 => 
        N_67_i_0, N_110_i_0 => N_110_i_0, N_112_i_0 => N_112_i_0, 
        N_114_i_0 => N_114_i_0, N_116_i_0 => N_116_i_0, N_69_i_0
         => N_69_i_0, N_71_i_0 => N_71_i_0, N_73_i_0 => N_73_i_0, 
        N_75_i_0 => N_75_i_0, N_77_i_0 => N_77_i_0, N_83_i_0 => 
        N_83_i_0, N_85_i_0 => N_85_i_0, N_133_i_0 => N_133_i_0, 
        N_87_i_0 => N_87_i_0, N_89_i_0 => N_89_i_0, N_140_i_0 => 
        N_140_i_0, N_91_i_0 => N_91_i_0, N_93_i_0 => N_93_i_0, 
        N_95_i_0 => N_95_i_0, N_97_i_0 => N_97_i_0, N_99_i_0 => 
        N_99_i_0, N_152_i_0 => N_152_i_0, N_101_i_0 => N_101_i_0, 
        N_156_i_0 => N_156_i_0, N_158_i_0 => N_158_i_0, N_103_i_0
         => N_103_i_0, N_105_i_0 => N_105_i_0, N_107_i_0 => 
        N_107_i_0, N_168_i_0 => N_168_i_0, N_109_i_0 => N_109_i_0, 
        N_111_i_0 => N_111_i_0, N_218_i_0 => N_218_i_0, N_217_i_0
         => N_217_i_0, N_203_i_0 => N_203_i_0);
    
    AHB_slave_dummy_0 : AHB_slave_dummy
      port map(waddr_in_net_0(4) => \waddr_in_net_0[4]\, 
        waddr_in_net_0(3) => \waddr_in_net_0[3]\, 
        waddr_in_net_0(2) => \waddr_in_net_0[2]\, 
        waddr_in_net_0(1) => \waddr_in_net_0[1]\, 
        waddr_in_net_0(0) => \waddr_in_net_0[0]\, 
        result_addr_net_0(3) => \result_addr_net_0[3]\, 
        result_addr_net_0(2) => \result_addr_net_0[2]\, 
        result_addr_net_0(1) => \result_addr_net_0[1]\, 
        result_addr_net_0(0) => \result_addr_net_0[0]\, 
        xhdl1222(5) => 
        \CertificationSystem_sb_0.CoreAHBLite_0.matrix4x16.xhdl1222[5]\, 
        CertificationSystem_sb_0_POWER_ON_RESET_N => 
        CertificationSystem_sb_0_POWER_ON_RESET_N, 
        CertificationSystem_sb_0_FAB_CCC_GL0 => 
        CertificationSystem_sb_0_FAB_CCC_GL0, N_276 => N_276, 
        N_203_i_0 => N_203_i_0, N_217_i_0 => N_217_i_0, N_218_i_0
         => N_218_i_0, N_259 => N_259, 
        CertificationSystem_sb_0_AHBmslave5_HREADY => 
        CertificationSystem_sb_0_AHBmslave5_HREADY, 
        AHB_slave_dummy_0_write_en => AHB_slave_dummy_0_write_en, 
        AHB_slave_dummy_0_read_en => AHB_slave_dummy_0_read_en, 
        N_277 => N_277, N_225 => N_225, N_206 => N_206, 
        un8_hreadyin_i_0 => 
        \CertificationSystem_sb_0.COREAHBLSRAM_0_0.U_CertificationSystem_sb_COREAHBLSRAM_0_0_AHBLSramIf.un8_hreadyin_i_0\, 
        N_226 => N_226);
    
    GPIO_0_M2F_obuf : OUTBUF
      port map(D => GPIO_0_M2F_c, PAD => GPIO_0_M2F);
    

end DEF_ARCH; 
